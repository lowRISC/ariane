/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module etherboot (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 5970;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h87fe7052_00000000,
        64'h87fe7090_00000000,
        64'h00000000_ffffffff,
        64'h00000006_00000000,
        64'h87feb3b0_cc33aa55,
        64'h00000000_2f7c5c2d,
        64'h00000000_87feb1f8,
        64'h00000000_ffffffff,
        64'h00006772_615f6473,
        64'h0000646d_635f6473,
        64'h00000000_0c000000,
        64'h00000000_ffffffff,
        64'h00000000_00000000,
        64'h00000000_30000000,
        64'h00000000_004b4d47,
        64'h00004b4d_47545045,
        64'h00000003_0f060301,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'haaaaaaaa_aaaaaaaa,
        64'h55555555_55555555,
        64'h5851f42d_4c957f2d,
        64'h10000000_20000000,
        64'h10325476_98badcfe,
        64'hefcdab89_67452301,
        64'h00000002_464c457f,
        64'hcccccccc_cccccccd,
        64'h00000a0d_70617274,
        64'h00000000_000a7473,
        64'h65742065_68636143,
        64'h00000000_00000a74,
        64'h6f6f6220_50544654,
        64'h00000000_00000a74,
        64'h73657420_4d415244,
        64'h00000000_00000a74,
        64'h6f6f6220_49505351,
        64'h00000000_00000000,
        64'h0a746f6f_62204453,
        64'h00000000_0000000a,
        64'h5825203d_20646565,
        64'h73206d6f_646e6152,
        64'h000a5825_2c582520,
        64'h3d20676e_69747465,
        64'h73206863_74697753,
        64'h0000000a_5825203d,
        64'h205d6425_5b707773,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h0a646c25_2e646c25,
        64'h203d2049_5043202c,
        64'h73656c63_79632064,
        64'h6c25202c_736e6f69,
        64'h74637572_74736e69,
        64'h20646c25_202c424b,
        64'h6425203d_20746573,
        64'h5f676e69_6b726f77,
        64'h00000000_00000000,
        64'h0a2e2979_6c6e6f28,
        64'h2032206e_6f697372,
        64'h65762065_736e6563,
        64'h694c2063_696c6275,
        64'h50206c61_72656e65,
        64'h4720554e_47206568,
        64'h74207265_646e7520,
        64'h6465736e_6563694c,
        64'h00000000_0000000a,
        64'h2e6e6f62_617a6143,
        64'h2073656c_72616843,
        64'h20323130_322d3130,
        64'h30322029_43282074,
        64'h68676972_79706f43,
        64'h00000000_0000000a,
        64'h29746962_2d642528,
        64'h20302e33_2e34206e,
        64'h6f697372_65762072,
        64'h65747365_746d656d,
        64'h00000a74_73657420,
        64'h4d415244_206c6174,
        64'h656d2065_7261420a,
        64'h00000a2e_656e6f44,
        64'h00000000_000a6b6f,
        64'h0000203a_73252020,
        64'h00000073_73657264,
        64'h6441206b_63757453,
        64'h00000000_00000a3a,
        64'h00000000_0075252f,
        64'h00752520_706f6f4c,
        64'h00000000_000a7025,
        64'h7830206f_74207025,
        64'h78302073_69206567,
        64'h6e617220_74736574,
        64'h00000000_00082008,
        64'h00000000_00000008,
        64'h08080808_08080808,
        64'h08082020_20202020,
        64'h20202020_20080808,
        64'h08080808_08080808,
        64'h00000000_0000000a,
        64'h2e2e2e74_73657420,
        64'h7478656e_206f7420,
        64'h676e6970_70696b53,
        64'h00000000_000a2e78,
        64'h25783020_74657366,
        64'h666f2074_6120656e,
        64'h696c2073_73657264,
        64'h64612064_61622065,
        64'h6c626973_736f7020,
        64'h3a455255_4c494146,
        64'h00000000_00007525,
        64'h20676e69_74736574,
        64'h00000000_00007525,
        64'h20676e69_74746573,
        64'h00000000_00080808,
        64'h08080808_08080808,
        64'h00000000_00202020,
        64'h20202020_20202020,
        64'h00000000_0000000a,
        64'h7025203d_20327020,
        64'h2c702520_3d203170,
        64'h00000a2e_78257830,
        64'h20746573_66666f20,
        64'h74612078_25783020,
        64'h3d212078_25783020,
        64'h3a455255_4c494146,
        64'h00000000_000a7325,
        64'h206e6f69_74636e75,
        64'h66202c64_2520656e,
        64'h696c202c_73252065,
        64'h6c696620_2c64656c,
        64'h69616620_7325206e,
        64'h6f697472_65737361,
        64'h00000a72_6564616f,
        64'h6c20746f_6f622065,
        64'h67617473_20747372,
        64'h69662064_65736162,
        64'h20746f6f_622d750a,
        64'h00000000_216b7369,
        64'h6420746e_756f6d75,
        64'h206f7420_6c696166,
        64'h00000000_0021656c,
        64'h69662065_736f6c63,
        64'h206f7420_6c696166,
        64'h0000000a_21746f6f,
        64'h62206e65_706f206f,
        64'h74206465_6c696146,
        64'h00000000_00000000,
        64'h6e69622e_746f6f62,
        64'h00000000_00000a79,
        64'h726f6d65_6d206f74,
        64'h6e69206e_69622e74,
        64'h6f6f6220_64616f4c,
        64'h00000000_0000000a,
        64'h21726576_69726420,
        64'h44532074_6e756f6d,
        64'h206f7420_6c696146,
        64'h00000000_0000000a,
        64'h2e2e2e70_25207373,
        64'h65726464_61207461,
        64'h206d6172_676f7270,
        64'h20646564_616f6c20,
        64'h65687420_746f6f42,
        64'h00000000_5c2d2f7c,
        64'h000a7825_203d206c,
        64'h61757463_61202c58,
        64'h25203d20_64657269,
        64'h75716572_206e656c,
        64'h00000000_00000000,
        64'h0a2e6e6f_69746172,
        64'h65706f20_50544654,
        64'h206c6167_656c6c49,
        64'h00000000_000a2e64,
        64'h656c6c61_63207172,
        64'h775f656c_646e6168,
        64'h00000000_00000a2e,
        64'h646e6520_656c6966,
        64'h20657669_65636552,
        64'h00000000_00000000,
        64'h0a64253d_657a6973,
        64'h6b636f6c_62202c22,
        64'h73252220_3a717277,
        64'h00000000_0000002f,
        64'h00000000_000a646c,
        64'h25202e67_6e6f6c20,
        64'h6f6f7420_68746170,
        64'h20747365_75716552,
        64'h00000064_6c252065,
        64'h646f6320_68746977,
        64'h2064656c_69616620,
        64'h64616572_20666c65,
        64'h000a7972_6f6d656d,
        64'h20524444_206f7420,
        64'h666c6520_64616f6c,
        64'h00000000_00000000,
        64'h0a732520_3d202964,
        64'h252c7025_2835646d,
        64'h00000000_0000000a,
        64'h6425203d_20687467,
        64'h6e656c20_656c6946,
        64'h00000000_00636d6d,
        64'h00000029_73252820,
        64'h00006425_203a7325,
        64'h00000000_00004453,
        64'h00000000_434d4d65,
        64'h00000000_00000000,
        64'h0a646e75_6f662074,
        64'h6f6e2064_25206563,
        64'h69766544_20434d4d,
        64'h0000297a_484d3030,
        64'h32282030_30325348,
        64'h00000000_00297a48,
        64'h4d383032_28203430,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282030,
        64'h35524444_20534855,
        64'h00000000_0000297a,
        64'h484d3030_31282030,
        64'h35524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282035,
        64'h32524453_20534855,
        64'h00000000_00000029,
        64'h7a484d35_32282032,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d32_35282032,
        64'h35524444_20434d4d,
        64'h0000297a_484d3235,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000029_7a484d30,
        64'h35282064_65657053,
        64'h20686769_48204453,
        64'h0000297a_484d3632,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000000_00000079,
        64'h63616765_4c204453,
        64'h00000000_00007963,
        64'h6167656c_20434d4d,
        64'h00000064_252e6425,
        64'h00000000_63256325,
        64'h63256325_63256325,
        64'h00000078_34302578,
        64'h34302520_726e5320,
        64'h78363025_206e614d,
        64'h00000000_00000a21,
        64'h646e756f_66206473,
        64'h635f7478_65206f4e,
        64'h00000000_00000000,
        64'h0a65646f_6d206120,
        64'h7463656c_6573206f,
        64'h7420656c_62616e75,
        64'h00000000_00000000,
        64'h0a217463_656c6573,
        64'h20656761_746c6f76,
        64'h206f7420_646e6f70,
        64'h73657220_746f6e20,
        64'h64696420_64726143,
        64'h0000000a_746e6573,
        64'h65727020_64726163,
        64'h206f6e20_3a434d4d,
        64'h00000000_0000000a,
        64'h64656e6f_69746974,
        64'h72617020_79646165,
        64'h726c6120_64726143,
        64'h00000000_000a7367,
        64'h6e697474_65732079,
        64'h74696c69_6261696c,
        64'h65722065_74697277,
        64'h206e6f69_74697472,
        64'h61702064_656c6c6f,
        64'h72746e6f_63207473,
        64'h6f682074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000a29_7525203e,
        64'h20752528_206d756d,
        64'h6978616d_20736465,
        64'h65637865_20657a69,
        64'h73206465_636e6168,
        64'h6e65206c_61746f54,
        64'h00000000_0000000a,
        64'h65747562_69727474,
        64'h61206465_636e6168,
        64'h6e652074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0a64656e,
        64'h67696c61_20657a69,
        64'h73207075_6f726720,
        64'h50572043_4820746f,
        64'h6e206e6f_69746974,
        64'h72617020_69255047,
        64'h0000000a_64656e67,
        64'h696c6120_657a6973,
        64'h2070756f_72672050,
        64'h57204348_20746f6e,
        64'h20616572_61206465,
        64'h636e6168_6e652061,
        64'h74616420_72657355,
        64'h00000a65_7a697320,
        64'h70756f72_67205057,
        64'h20434820_656e6966,
        64'h65642074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_000a676e,
        64'h696e6f69_74697472,
        64'h61702074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0000000a,
        64'h61657261_20617461,
        64'h64207265_73752064,
        64'h65636e61_686e6520,
        64'h726f6620_64657269,
        64'h75716572_20342e34,
        64'h203d3e20_434d4d65,
        64'h00000000_000a2978,
        64'h6c257830_2878616d,
        64'h20736465_65637865,
        64'h20786c25_78302072,
        64'h65626d75_6e206b63,
        64'h6f6c6220_3a434d4d,
        64'h00000000_00000a64,
        64'h6d632070_6f747320,
        64'h646e6573_206f7420,
        64'h6c696166_20636d6d,
        64'h00000000_000a7964,
        64'h61657220_64726163,
        64'h20676e69_74696177,
        64'h2074756f_656d6954,
        64'h0000000a_58383025,
        64'h7830203a_726f7272,
        64'h45207375_74617453,
        64'h00000000_65646f6d,
        64'h206e776f_6e6b6e55,
        64'h00000000_00006473,
        64'h5f637369_72776f6c,
        64'h00000078_25782520,
        64'h00000020_3a78250a,
        64'h00000000_0a732574,
        64'h69622d64_25203a68,
        64'h74646957_20737542,
        64'h00000000_0000203a,
        64'h79746963_61706143,
        64'h00000000_00000a73,
        64'h25203a79_74696361,
        64'h70614320_68676948,
        64'h00000a64_25203a64,
        64'h65657053_20737542,
        64'h00000000_00000a20,
        64'h63256325_63256325,
        64'h6325203a_656d614e,
        64'h00000000_00000000,
        64'h0a782520_3a4d454f,
        64'h00000000_0a782520,
        64'h3a444920_72657275,
        64'h74636166_756e614d,
        64'h00000000_000a7325,
        64'h203a6563_69766544,
        64'h00202020_3a434d4d,
        64'h00000000_52444420,
        64'h00000000_00006f4e,
        64'h00000000_00736559,
        64'h0000000a_7825203d,
        64'h2074736f_68202c78,
        64'h25207461_20646574,
        64'h61657263_20636d6d,
        64'h00000000_00000a64,
        64'h25206f74_20646567,
        64'h6e616863_206b7361,
        64'h6d202c64_65747265,
        64'h736e6920_64726143,
        64'h00000000_0000000a,
        64'h6425206f_74206465,
        64'h676e6168_63206b73,
        64'h616d202c_6465766f,
        64'h6d657220_64726143,
        64'h000a7475_6f656d69,
        64'h74207325_203a6473,
        64'h5f637369_72776f6c,
        64'h00726464_615f6573,
        64'h61625f64_73203d3d,
        64'h20657361_625f6473,
        64'h00000000_00000063,
        64'h2e636d6d_5f637369,
        64'h72776f6c_2f637273,
        64'h00000000_00000000,
        64'h66656463_62613938,
        64'h37363534_33323130,
        64'h007f7c5d_5b3f3e3d,
        64'h3c3b3a2e_2c2b2a22,
        64'h00007f7c_5d5b3f3e,
        64'h3d3c3b3a_2c2b2a22,
        64'h0000000a_2e783230,
        64'h253a7832_30253a78,
        64'h3230253a_78323025,
        64'h3a783230_253a7832,
        64'h3025203d_20737365,
        64'h72646461_2043414d,
        64'h00000a78_6c253a78,
        64'h6c25203d_2043414d,
        64'h00000000_00000a78,
        64'h25203d20_5d64255b,
        64'h4d454f20_49505351,
        64'h000a7264_64612043,
        64'h414d2070_75746553,
        64'h0000000a_21747075,
        64'h72726574_6e692064,
        64'h656c646e_61686e75,
        64'h00000000_00000a78,
        64'h25783020_3d206570,
        64'h79745f6f_746f7270,
        64'h00000000_0a297825,
        64'h28206465_74726f70,
        64'h7075736e_75203d20,
        64'h6f746f72_70205049,
        64'h000a5741_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a534c50_4d203d20,
        64'h6f746f72_50205049,
        64'h00000000_000a4554,
        64'h494c5044_55203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505443_53203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a504d4f_43203d20,
        64'h6f746f72_50205049,
        64'h00000000_0000004d,
        64'h00000000_0000000a,
        64'h5041434e_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000a48,
        64'h50544545_42203d20,
        64'h6f746f72_50205049,
        64'h000a5054_4d203d20,
        64'h6f746f72_50205049,
        64'h00000a48_41203d20,
        64'h6f746f72_50205049,
        64'h000a5053_45203d20,
        64'h6f746f72_50205049,
        64'h000a4552_47203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505653_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000036,
        64'h00000000_00000000,
        64'h0a504343_44203d20,
        64'h6f746f72_50205049,
        64'h00000a50_54203d20,
        64'h6f746f72_50205049,
        64'h000a5044_49203d20,
        64'h6f746f72_50205049,
        64'h000a3a73_746e6574,
        64'h6e6f6320_74736574,
        64'h0000000a_3a726564,
        64'h61656820_74736574,
        64'h000a5055_50203d20,
        64'h6f746f72_50205049,
        64'h000a5047_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000054,
        64'h00000000_00000000,
        64'h0a504950_49203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000047,
        64'h00006425_2b544553,
        64'h46464f5f_524c5052,
        64'h00000000_3f3f3f3f,
        64'h00000000_00544553,
        64'h46464f5f_524c5052,
        64'h00000000_00544553,
        64'h46464f5f_44414252,
        64'h00000000_00005445,
        64'h5346464f_5f525352,
        64'h00000000_00544553,
        64'h46464f5f_53434652,
        64'h00544553_46464f5f,
        64'h4c525443_4f49444d,
        64'h00000000_00544553,
        64'h46464f5f_53434654,
        64'h00000000_00544553,
        64'h46464f5f_524c5054,
        64'h00000000_54455346,
        64'h464f5f49_4843414d,
        64'h00000000_54455346,
        64'h464f5f4f_4c43414d,
        64'h00000000_000a3b29,
        64'h78257830_2c302c78,
        64'h25287465_736d656d,
        64'h00000000_0a3b2978,
        64'h2578302c_78257830,
        64'h2c782528_6e666c65,
        64'h00000a70_2520726f,
        64'h72726520_7974696e,
        64'h61732072_64646170,
        64'h00000020_3a5d6425,
        64'h5b6e6f69_74636553,
        64'h000a7325_20202020,
        64'h00786c6c_2a302520,
        64'h00003a78_6c383025,
        64'h00732542_69632520,
        64'h00000000_00732573,
        64'h65747942_20756c25,
        64'h0073257a_48632520,
        64'h00000000_646c252e,
        64'h00000000_00756c25,
        64'h00000000_00000000,
        64'h73257a48_20756c25,
        64'h00000000_00007325,
        64'h00000000_00732520,
        64'h3a646c69_7542202c,
        64'h00000000_73257325,
        64'h00000000_00000a0a,
        64'h00000058_32302520,
        64'h00000000_0000002e,
        64'h00000000_00006325,
        64'h00000000_00000020,
        64'h20202020_20202020,
        64'h000a5245_46464f5f,
        64'h50434844_20726f66,
        64'h20676e69_74696157,
        64'h00000a73_25203a73,
        64'h25206563_69766564,
        64'h206e6f20_59524556,
        64'h4f435349_44205043,
        64'h48442064_6e657320,
        64'h74276e64_6c756f43,
        64'h000a5832_30253a58,
        64'h3230253a_58323025,
        64'h3a583230_253a5832,
        64'h30253a58_32302520,
        64'h3a204341_4d207325,
        64'h00000000_30687465,
        64'h00000000_000a2973,
        64'h2528726f_72726570,
        64'h000a5952_45564f43,
        64'h5349445f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_0000000a,
        64'h64252065_646f6370,
        64'h6f205043_48442064,
        64'h656c646e_61686e55,
        64'h00000000_0a642520,
        64'h6e6f6974_706f2064,
        64'h656c646e_61686e75,
        64'h00000000_0000000a,
        64'h73252072_6f727245,
        64'h00000000_00000a64,
        64'h65737566_65722073,
        64'h73657264_64612064,
        64'h65747365_75716552,
        64'h00000000_0000000a,
        64'h4b414e20_50434844,
        64'h00000000_0a444550,
        64'h50494b53_204b4341,
        64'h000a2273_2522203d,
        64'h20656d61_6e74736f,
        64'h4820746e_65696c43,
        64'h00000a22_73252220,
        64'h3d206e69_616d6f44,
        64'h00000000_0000000a,
        64'h7364253a_6d64253a,
        64'h68642520_3d20656d,
        64'h69742065_7361654c,
        64'h000a6425_2e64252e,
        64'h64252e64_2520203a,
        64'h73736572_64646120,
        64'h6b73616d_2074654e,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h61207265_74756f52,
        64'h00000000_00000000,
        64'h0a64252e_64252e64,
        64'h252e6425_20203a73,
        64'h73657264_64412050,
        64'h49207265_76726553,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h41205049_20746e65,
        64'h696c4320_50434844,
        64'h00000000_0000000a,
        64'h4b434120_50434844,
        64'h0000000a_54534555,
        64'h5145525f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_00000000,
        64'h0a702520_2c726f72,
        64'h7265206c_616e7265,
        64'h746e6920_70636864,
        64'h00000a29_73252c73,
        64'h25287075_6b6f6f6c,
        64'h000a6563_69766564,
        64'h206e776f_6e6b6e75,
        64'h00000000_203a6425,
        64'h20656369_7665440a,
        64'h00203a64_25206563,
        64'h69766564_2073250a,
        64'h00000000_00203a64,
        64'h25206563_69766544,
        64'h00000000_00000000,
        64'h73736572_6464612d,
        64'h63616d2d_6c61636f,
        64'h6c006874_6469772d,
        64'h6f692d67_65720074,
        64'h66696873_2d676572,
        64'h00737470_75727265,
        64'h746e6900_746e6572,
        64'h61702d74_70757272,
        64'h65746e69_00646565,
        64'h70732d74_6e657272,
        64'h75630076_65646e2c,
        64'h76637369_72007974,
        64'h69726f69_72702d78,
        64'h616d2c76_63736972,
        64'h0073656d_616e2d67,
        64'h65720064_65646e65,
        64'h7478652d_73747075,
        64'h72726574_6e690073,
        64'h65676e61_7200656c,
        64'h646e6168_702c7875,
        64'h6e696c00_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h00100000_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_00000064,
        64'h6e727768_2d637369,
        64'h72776f6c_1b000000,
        64'h0e000000_03000000,
        64'h00003030_30303030,
        64'h30344064_6e727768,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h00800000_00000000,
        64'h00000030_00000000,
        64'h67000000_10000000,
        64'h03000000_00007fe3,
        64'h023e1800_47010000,
        64'h06000000_03000000,
        64'h03000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_00636d6d,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_02000000,
        64'h25010000_04000000,
        64'h03000000_02000000,
        64'h14010000_04000000,
        64'h03000000_00000100,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40636d6d,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h04000000_3a010000,
        64'h04000000_03000000,
        64'h02000000_30010000,
        64'h04000000_03000000,
        64'h01000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h00c20100_06010000,
        64'h04000000_03000000,
        64'h80f0fa02_4b000000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000010_00000000,
        64'h67000000_10000000,
        64'h03000000_00303537,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000000,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'hffff0000_01000000,
        64'hca000000_08000000,
        64'h03000000_00333130,
        64'h2d677562_65642c76,
        64'h63736972_1b000000,
        64'h10000000_03000000,
        64'h00003040_72656c6c,
        64'h6f72746e_6f632d67,
        64'h75626564_01000000,
        64'h02000000_02000000,
        64'hbb000000_04000000,
        64'h03000000_02000000,
        64'hb5000000_04000000,
        64'h03000000_03000000,
        64'hfb000000_04000000,
        64'h03000000_07000000,
        64'he8000000_04000000,
        64'h03000000_00000004,
        64'h00000000_0000000c,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h09000000_01000000,
        64'h0b000000_01000000,
        64'hca000000_10000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00000c00,
        64'h00000000_00000002,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_01000000,
        64'h03000000_01000000,
        64'hca000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6e696c63,
        64'h01000000_c3000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000008_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h01000000_bb000000,
        64'h04000000_03000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00007663_73697200,
        64'h656e6169_7261202c,
        64'h7a687465_1b000000,
        64'h13000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha8060000_59010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'he0060000_38000000,
        64'h39080000_edfe0dd0,
        64'h00000000_fffffa0a,
        64'hfffff9d0_fffff9f8,
        64'hfffff9d0_fffff9e6,
        64'hfffff9d2_fffff9be,
        64'h00000000_64726143,
        64'h2d445320_726f6620,
        64'h746f6f62_2d752064,
        64'h6573696d_696e696d,
        64'h20435349_52776f4c,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00020000_00010000,
        64'h0000c000_00008000,
        64'h00006000_00004000,
        64'h00002000_00001000,
        64'h00000800_00000400,
        64'h00000200_00000100,
        64'h00000080_00000040,
        64'h00000020_00000000,
        64'h0bebc200_0c65d400,
        64'h02faf080_05f5e100,
        64'h02faf080_017d7840,
        64'h03197500_03197500,
        64'h02faf080_018cba80,
        64'h017d7840_017d7840,
        64'h00989680_000f4240,
        64'h000186a0_00002710,
        64'h50463c37_322d2823,
        64'h1e19140f_0d0c0a00,
        64'h00000000_00000000,
        64'h00000000_10000000,
        64'h00000001_00000000,
        64'h20000000_00000002,
        64'h00000000_40000000,
        64'h00000005_00000001,
        64'h20000000_00000006,
        64'h00000001_40000000,
        64'h70000000_00000000,
        64'h70000000_00000002,
        64'h70000000_00000004,
        64'h60000000_00000005,
        64'h30000000_00000001,
        64'h30000000_00000003,
        64'h00000000_40050100,
        64'h40050000_40040500,
        64'h40040401_40040400,
        64'h40040300_40040200,
        64'h40040100_40040000,
        64'h00000000_87feb360,
        64'h00000000_87feb348,
        64'h00000000_87feb330,
        64'h00000000_87feb318,
        64'h00000000_87feb300,
        64'h00000000_87feb2e8,
        64'h00000000_87feb2d0,
        64'h00000000_87feb2b8,
        64'h00000000_87feb2a0,
        64'h00000000_87feb288,
        64'h00000000_87feb278,
        64'h00000000_87feb268,
        64'hffffbb7e_ffffbb7e,
        64'hffffbb7e_ffffbb7e,
        64'hffffbb7a_ffffbb76,
        64'hffffbb76_ffffbb50,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_87fe4d04,
        64'h00000000_87fe4aa6,
        64'h00000000_87fe4e98,
        64'h00646374_65675f63,
        64'h6d6d5f64_72616f62,
        64'h00000002_0000ffff,
        64'h004c4b40_004c4b40,
        64'h00300000_20000000,
        64'h00000000_87fe9c88,
        64'h00000000_87feaf50,
        64'h00717269_5f646e65,
        64'h5f617461_645f6473,
        64'h5f637369_72776f6c,
        64'h00000000_00007172,
        64'h695f646d_635f6473,
        64'h5f637369_72776f6c,
        64'h00007172_695f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0067616c,
        64'h665f7470_75727265,
        64'h746e695f_74696177,
        64'h5f637369_72776f6c,
        64'h00000000_646d635f,
        64'h74726174_735f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0000006e,
        64'h655f7172_695f6473,
        64'h00000000_00007475,
        64'h6f656d69_745f6473,
        64'h00000000_0000657a,
        64'h69736b6c_625f6473,
        64'h00000000_00000074,
        64'h6e636b6c_625f6473,
        64'h00000000_00000000,
        64'h74657365_725f6473,
        64'h00000000_74726174,
        64'h735f646d_635f6473,
        64'h00000000_0000676e,
        64'h69747465_735f6473,
        64'h00000000_00007669,
        64'h645f6b6c_635f6473,
        64'h00000000_00000000,
        64'h6e67696c_615f6473,
        64'h00000000_00006465,
        64'h6c5f7465_735f6473,
        64'h5f637369_72776f6c,
        64'h09020b04_0d060f08,
        64'h010a030c_050e0700,
        64'h020f0c09_0603000d,
        64'h0a070401_0e0b0805,
        64'h0c07020d_08030e09,
        64'h040f0a05_000b0601,
        64'heb86d391_2ad7d2bb,
        64'hbd3af235_f7537e82,
        64'h4e0811a1_a3014314,
        64'hfe2ce6e0_6fa87e4f,
        64'h85845dd1_ffeff47d,
        64'h8f0ccc92_655b59c3,
        64'hfc93a039_ab9423a7,
        64'h432aff97_f4292244,
        64'hc4ac5665_1fa27cf8,
        64'he6db99e5_d9d4d039,
        64'h04881d05_d4ef3085,
        64'heaa127fa_289b7ec6,
        64'hbebfbc70_f6bb4b60,
        64'h4bdecfa9_a4beea44,
        64'hfde5380c_6d9d6122,
        64'h8771f681_fffa3942,
        64'h8d2a4c8a_676f02d9,
        64'hfcefa3f8_a9e3e905,
        64'h455a14ed_f4d50d87,
        64'hc33707d6_21e1cde6,
        64'he7d3fbc8_d8a1e681,
        64'h02441453_d62f105d,
        64'he9b6c7aa_265e5a51,
        64'hc040b340_f61e2562,
        64'h49b40821_a679438e,
        64'hfd987193_6b901122,
        64'h895cd7be_ffff5bb1,
        64'h8b44f7af_698098d8,
        64'hfd469501_a8304613,
        64'h4787c62a_f57c0faf,
        64'hc1bdceee_242070db,
        64'he8c7b756_d76aa478,
        64'h02020202_02020202,
        64'h10020202_02020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02010101_01010101,
        64'h10010101_01010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h08101010_10020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02424242_42424210,
        64'h10101010_10010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h01414141_41414110,
        64'h10101010_10100404,
        64'h04040404_04040404,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h08080808_08080808,
        64'h08080808_08080808,
        64'h08082828_28282808,
        64'h08080808_08080808,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_bf5dd0ff,
        64'hf0efef3f_b0ef07e5,
        64'h05130000_2517b7e1,
        64'he14f80ef_f05fb0ef,
        64'h08050513_00002517,
        64'hbfe9c37f_f0eff17f,
        64'hb0ef0825_05130000,
        64'h2517b7f5_edbff0ef,
        64'h8522f2bf_b0ef0865,
        64'h05130000_2517a001,
        64'haa9fe0ef_8522f3ff,
        64'hb0ef08a5_05130000,
        64'h25178782_97ba439c,
        64'h97ba078a_65470713,
        64'h00000717_02f76463,
        64'h47190054_579b0ff4,
        64'h7413fd39_1be3f6ff,
        64'hb0ef2581_8552688c,
        64'h0004b823_f7dfb0ef,
        64'h86222401_25816080,
        64'h608ce09c_09058556,
        64'h0007c783_016907b3,
        64'h49910caa_0a130000,
        64'h2a170baa_8a930000,
        64'h2a974000_04b727eb,
        64'h0b130000_2b174901,
        64'hda0f80ef_fe9416e3,
        64'hfc1fb0ef_0405854a,
        64'h0004059b_6390078e,
        64'h013407b3_44950de9,
        64'h09130000_29170800,
        64'h09b74401_935fe0ef,
        64'h0e050513_00002517,
        64'h90ffe0ef_e05ae456,
        64'he852ec4e_f04af426,
        64'hf822fc06_7139957f,
        64'he06f1a25_05130000,
        64'h2517b4ff_e06f0141,
        64'h60a281af_c06f0141,
        64'hc9050513_00002517,
        64'h40a005b3_60a20005,
        64'h5c63d35f_70eff885,
        64'h05130000_051783ef,
        64'hc0efe406_c9c50513,
        64'h00002517_1141bf6d,
        64'h00fab023_04a19381,
        64'h178200c4_579b2421,
        64'hf51ff0ef_85a68082,
        64'h61616ae2_7a0279a2,
        64'h794274e2_640660a6,
        64'hecbfd0ef_92018526,
        64'h002c1602_4089063b,
        64'hf79ff0ef_002c0334,
        64'h66630144_053b4000,
        64'h0ab7ff86_099b4401,
        64'h89328a2e_84aae486,
        64'hec56f052_f44ef84a,
        64'hfc26e0a2_715d8082,
        64'h61056442_60e2fee7,
        64'h9ae30585_37e100d5,
        64'h802300f5_56b35761,
        64'h03800793_85a2f4ff,
        64'hf0ef454d_46010034,
        64'h4589f5bf_f0efec06,
        64'hc43e454d_45894601,
        64'h0034842e_c62ae822,
        64'h8fd90585_65133007,
        64'h07131101_0085151b,
        64'h67050185_579b9d3d,
        64'h00b007b7_a1ffe06f,
        64'h014160a2_64020004,
        64'h4503943e_20478793,
        64'h00002797_883dfebf,
        64'hf0ef2501_35fd0045,
        64'h551b00b7_d863842a,
        64'h4785e406_e0221141,
        64'hbfe1f710_06912785,
        64'h0006e603_80827388,
        64'h400007b7_ffe537fd,
        64'hc3198b09_7a984000,
        64'h06b73e80_079300b7,
        64'hef634000_07374781,
        64'h2581f788_8d514000,
        64'h07b70106_161b8d5d,
        64'h0085979b_80822501,
        64'h7b884000_07b78082,
        64'h25016b88_0007b823,
        64'h400007b7_80822501,
        64'h63884000_07b78082,
        64'he3884000_07b79101,
        64'h1502bff1_f5dff0ef,
        64'h4541f63f_f0ef4521,
        64'hf69ff0ef_4511f6ff,
        64'hf0ef4509_f75ff0ef,
        64'h4505f7bf_f0ef4501,
        64'he4061141_bf51c000,
        64'h28f3c020_26f3fac7,
        64'h10e39f2f_c06f28e5,
        64'h05130000_251702a7,
        64'h473302a7_67b302b3,
        64'h45bb02c7_47334000,
        64'h059302a6_87334116,
        64'h86b33e80_0513c000,
        64'h26f38e15_c0202673,
        64'h02b71d63_2705fe08,
        64'h13e397aa_387d0007,
        64'h802397aa_00078023,
        64'h97aa0007_802397aa,
        64'h00078023_40000813,
        64'h87f245a9_01f61e13,
        64'h46814881_470100c5,
        64'h131b4605_80828082,
        64'h614569a2_694264e2,
        64'h740270a2_ff2417e3,
        64'he6dff0ef_24050135,
        64'h85334605_46850084,
        64'h95b34979_01f49993,
        64'h4441a92f_c0ef4485,
        64'h03050513_00002517,
        64'haa0fc0ef_2f450513,
        64'h00002517_aacfc0ef,
        64'h2d050513_00002517,
        64'hab8fc0ef_2b450513,
        64'h00002517_04000593,
        64'hc19fe0ef_e44ee84a,
        64'hec26f022_f4062b65,
        64'h05130000_25177179,
        64'hbfa10485_ae4fc0ef,
        64'h08050513_00002517,
        64'hb7e94a89_af4fc0ef,
        64'h2c850513_00002517,
        64'h97828522_85ce6642,
        64'h008a3783_b0cfc0ef,
        64'h2d850513_00002517,
        64'hc58d000a_358302f7,
        64'h49636762_010a2783,
        64'hb28fc0ef_856eed15,
        64'h920ff0ef_852265a2,
        64'hb38fc0ef_856a85e6,
        64'hb40fc0ef_8562b46f,
        64'hc0ef855e_85ca0009,
        64'h0663b52f_c0ef855a,
        64'h85a68082_61497da2,
        64'h7d427ce2_6c066ba6,
        64'h6b466ae6_7a0679a6,
        64'h794674e6_8556640a,
        64'h60aab7af_c0ef3565,
        64'h05130000_25170299,
        64'h7863e72a_0a130000,
        64'h3a17362d_8d930000,
        64'h2d97362d_0d130000,
        64'h2d1735ac_8c930000,
        64'h2c9735ac_0c130000,
        64'h2c1735ab_8b930000,
        64'h2b9735ab_0b130000,
        64'h2b174485_4a81e43e,
        64'h99a20034_d793e83e,
        64'h0014d993_0044d793,
        64'hbd8fc0ef_ec36e506,
        64'hf46ef86a_fc66e0e2,
        64'he4dee8da_ecd6f0d2,
        64'hf4ce3725_05130000,
        64'h251785aa_962a84ae,
        64'h842afca6_e122fff5,
        64'h86138932_f8ca7175,
        64'h80826505_b789547d,
        64'hbf290d85_e73fe0ef,
        64'h0007c503_97ea8b8d,
        64'h00078b1b_001b079b,
        64'he87fe0ef_4521ef91,
        64'h034df7b3_00f69323,
        64'h93c117c2_0064d783,
        64'h00f69223_93c117c2,
        64'h0044d783_00f69123,
        64'h93c117c2_0024d783,
        64'h00f69023_93c117c2,
        64'h0004d783_e38866c2,
        64'h67e2f6a7_bd230000,
        64'h37978d41_91011402,
        64'h15028c51_8d590106,
        64'h161b0105_151b6702,
        64'h6622fdbf_d0efe02a,
        64'hfe1fd0ef_e42afe7f,
        64'hd0ef842a_fedfd0ef,
        64'he836ec3e_b7758c4a,
        64'h8bce4a85_80826149,
        64'h7da27d42_7ce26c06,
        64'h6ba66b46_6ae67a06,
        64'h79a67946_74e6640a,
        64'h60aa8522_cd4fc0ef,
        64'h45050513_00002517,
        64'h020a8863_e579842a,
        64'ha82ff0ef_854a85ce,
        64'h866e059d_956397de,
        64'h00fc06b3_003d9793,
        64'h4d818c4e_8bca7ced,
        64'h0d130000_2d179c4a,
        64'h0a1301a4_84930000,
        64'h34974a81_f73fe0ef,
        64'h4b018cb2_f46ee122,
        64'he506f86a_fc66e0e2,
        64'he4dee8da_ecd6fca6,
        64'h6a050200_051389ae,
        64'h892af0d2_f4cef8ca,
        64'h7175bfa1_547dbf0d,
        64'h0d85fa9f_e0ef0007,
        64'hc50397e6_8b8d0007,
        64'h8a9b001a_879bfbdf,
        64'he0ef4521_ef910ba1,
        64'h033df7b3_ffa795e3,
        64'h00d60023_0ff6f693,
        64'h078500fb_86330006,
        64'hc6830187_86b34781,
        64'he28808a7_b9230000,
        64'h37978d41_66e29101,
        64'h14021502_8c510106,
        64'h161b8d5d_0105151b,
        64'h664267a2_8fcfe0ef,
        64'he42a902f_e0efe82a,
        64'h908fe0ef_842a90ef,
        64'he0efec36_b7758ba6,
        64'h8b4a4a05_80826149,
        64'h7da27d42_7ce26c06,
        64'h6ba66b46_6ae67a06,
        64'h79a67946_74e6640a,
        64'h60aa8522_df4fc0ef,
        64'h57050513_00002517,
        64'h020a0863_ed45842a,
        64'hba2ff0ef_852685ca,
        64'h866e04fd_956396da,
        64'h003d9693_67824d21,
        64'h4d818bca_8b268eec,
        64'h8c930000_3c979c49,
        64'h8993132c_0c130000,
        64'h3c174a01_892ff0ef,
        64'h4a81e032_f46ef86a,
        64'he122e506_fc66e0e2,
        64'he4dee8da_ecd6f0d2,
        64'h69850200_0513892e,
        64'h84aaf4ce_f8cafca6,
        64'h7175b7e9_5b7db749,
        64'h060500b8_3023e30c,
        64'h85d6e111_85e20016,
        64'h75138082_61096de2,
        64'h7d027ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_855a7446,
        64'h70e6ea2f_c0ef5f65,
        64'h05130000_2517fafb,
        64'h90e30400_07932b85,
        64'hfbb41be3_8c562405,
        64'he9318b2a_c5eff0ef,
        64'h854a85ce_6622ecef,
        64'hc0ef856a_85daed6f,
        64'hc0efe432_855206f6,
        64'h1063974e_00e90833,
        64'h00361713_67824601,
        64'hfffc4a93_ef4fc0ef,
        64'h856685da_00848b3b,
        64'hf00fc0ef_85524401,
        64'h003b949b_01779c33,
        64'h47854da1_5fcd0d13,
        64'h00002d17_5f4c8c93,
        64'h00002c97_5eca0a13,
        64'h00002a17_f2cfc0ef,
        64'h4b81e032_89aef862,
        64'he0dae4d6_f4a6f8a2,
        64'hfc86ec6e_f06af466,
        64'hfc5ee8d2_ecce6065,
        64'h05130000_2517892a,
        64'hf0ca7119_bf755dfd,
        64'hbfc585ba_fe081be3,
        64'h85c6b761_0605e10c,
        64'he28c85be_00081363,
        64'h859a008b_ea630016,
        64'h78138082_61096de2,
        64'h7d027ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_856e7446,
        64'h70e6fa2f_c0ef6f65,
        64'h05130000_2517f8f4,
        64'h1be30800_07932405,
        64'hed298daa_d56ff0ef,
        64'h852685ca_6622fc6f,
        64'hc0ef8566_85a2fcef,
        64'hc0efe432_854e0546,
        64'h1c6396ca_00d48533,
        64'h00361693_4601fff7,
        64'hc313fff7_48938fd5,
        64'h008d16b3_00fd17b3,
        64'h0024079b_8f5d00ed,
        64'h173300fd_17b3408b,
        64'h07bb408a_873b80ff,
        64'hc0ef8562_85a2817f,
        64'hc0ef854e_704c8c93,
        64'h00002c97_03f00b93,
        64'h08100b13_4d0507f0,
        64'h0a9370ac_0c130000,
        64'h2c177029_89930000,
        64'h2997843f_c0ef4401,
        64'h8a32892e_ec6efc86,
        64'hf06af466_f862fc5e,
        64'he0dae4d6_e8d2ecce,
        64'hf0caf8a2_71c50513,
        64'h00002517_84aaf4a6,
        64'h7119b7f1_5dfdbfe5,
        64'he19ce31c_bf610605,
        64'he194e314_008c6663,
        64'h80826109_6de27d02,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e67906,
        64'h74a6856e_744670e6,
        64'h8a9fc0ef_7fc50513,
        64'h00002517_fb5417e3,
        64'h2405e139_8daae58f,
        64'hf0ef8526_85ca6622,
        64'h8c9fc0ef_856a85a2,
        64'h8d1fc0ef_e4328552,
        64'h05661a63_974a00e4,
        64'h85b30036_17134601,
        64'hfff6c693_fff7c793,
        64'h008996b3_00f997b3,
        64'h408b87bb_8fdfc0ef,
        64'h856685a2_905fc0ef,
        64'h85520800_0a937f6d,
        64'h0d130000_2d1703f0,
        64'h0c134985_07f00b93,
        64'h7f8c8c93_00002c97,
        64'h7f0a0a13_00002a17,
        64'h931fc0ef_44018b32,
        64'h892eec6e_fc86f06a,
        64'hf466f862_fc5ee0da,
        64'he4d6e8d2_eccef0ca,
        64'hf8a280a5_05130000,
        64'h351784aa_f4a67119,
        64'hb7f15dfd_bfe5e298,
        64'he398bf61_0605e28c,
        64'he38c008c_66638082,
        64'h61096de2_7d027ca2,
        64'h7c427be2_6b066aa6,
        64'h6a4669e6_790674a6,
        64'h856e7446_70e6997f,
        64'hc0ef8ea5_05130000,
        64'h3517fb54_1be32405,
        64'he1398daa_f46ff0ef,
        64'h852685ca_66229b7f,
        64'hc0ef856a_85a29bff,
        64'hc0efe432_85520566,
        64'h1a6397ca_00f486b3,
        64'h00361793_46010089,
        64'h95b300e9_9733408b,
        64'h873b9e3f_c0ef8566,
        64'h85a29ebf_c0ef8552,
        64'h08000a93_8dcd0d13,
        64'h00003d17_03f00c13,
        64'h498507f0_0b938dec,
        64'h8c930000_3c978d6a,
        64'h0a130000_3a17a17f,
        64'hc0ef4401_8b32892e,
        64'hec6efc86_f06af466,
        64'hf862fc5e_e0dae4d6,
        64'he8d2ecce_f0caf8a2,
        64'h8f050513_00003517,
        64'h84aaf4a6_7119bff1,
        64'h59fdb74d_0605e29c,
        64'he31c8082_61256c42,
        64'h6be27b02_7aa27a42,
        64'h79e26906_64a6854e,
        64'h644660e6_a6dfc0ef,
        64'h9c050513_00003517,
        64'hf94c19e3_0c05e91d,
        64'h89aa81df_f0ef8522,
        64'h85a66622_a8dfc0ef,
        64'h855e85ce_a95fc0ef,
        64'he432854a_05561763,
        64'h972600e4_06b30036,
        64'h17134601_8fd9038c,
        64'h17138fd9_030c1713,
        64'h8fd9028c_17138fd9,
        64'h020c1713_8fd9018c,
        64'h17130187_e7b38fd9,
        64'h010c1793_008c1713,
        64'had9fc0ef_855a85ce,
        64'h000c099b_ae5fc0ef,
        64'h854a1000_0a139d6b,
        64'h8b930000_3b979ceb,
        64'h0b130000_3b179c69,
        64'h09130000_3917b07f,
        64'hc0ef4c01_8ab284ae,
        64'hfc4eec86_e862ec5e,
        64'hf05af456_f852e0ca,
        64'he4a69da5_05130000,
        64'h3517842a_e8a2711d,
        64'hb7e15d7d_b7790605,
        64'he198e398_872ac291,
        64'h876a0016_7693bf49,
        64'h000b3d03_80826165,
        64'h6d426ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h694664e6_856a7406,
        64'h70a6b6bf_c0efabe5,
        64'h05130000_3517fb44,
        64'h1ae32405_e5298d2a,
        64'h91bff0ef_852685ca,
        64'h6622b8bf_c0ef8566,
        64'h85a2b93f_c0efe432,
        64'h854e0556_1c6397ca,
        64'h00f485b3_00361793,
        64'hfffd4513_4601baff,
        64'hc0ef8562_85a2000b,
        64'hbd03cba5_00147793,
        64'hbc1fc0ef_854e0400,
        64'h0a13ab2c_8c930000,
        64'h3c97aaac_0c130000,
        64'h3c17db2b_8b930000,
        64'h3b97db2b_0b130000,
        64'h3b17ab29_89930000,
        64'h3997bf3f_c0ef4401,
        64'h8ab2892e_e86af486,
        64'hec66f062_f45ef85a,
        64'hfc56e0d2_e4cee8ca,
        64'hf0a2aca5_05130000,
        64'h351784aa_eca67159,
        64'hbfc154fd_bf590605,
        64'he198e398_8726c291,
        64'h87660016_76938082,
        64'h61656ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h64e66946_85267406,
        64'h70a6c53f_c0efba65,
        64'h05130000_3517fb54,
        64'h1be32405_e12984aa,
        64'ha03ff0ef_854a85ce,
        64'h6622c73f_c0ef8562,
        64'h85a2c7bf_c0efe432,
        64'h85520566_186397ce,
        64'h00f905b3_00361793,
        64'h14fd4601_40900cb3,
        64'hc99fc0ef_8885855e,
        64'h85a2fff4_4493ca7f,
        64'hc0ef8552_04000a93,
        64'hb98c0c13_00003c17,
        64'hb90b8b93_00003b97,
        64'hb88a0a13_00003a17,
        64'hcc9fc0ef_44018b32,
        64'h89aeec66_eca6f486,
        64'hf062f45e_f85afc56,
        64'he0d2e4ce_f0a2b9e5,
        64'h05130000_3517892a,
        64'he8ca7159_bfc90705,
        64'h00a83023_e28800f7,
        64'h0533a9df_f06f6121,
        64'h863a69e2_854e7902,
        64'h74a270e2_744200c7,
        64'h1c6396ae_00d98833,
        64'h00371693_47018fc5,
        64'h90811782_65a26602,
        64'h14828fc1_8cc90109,
        64'h179b0105_151b887f,
        64'he0ef84aa_88dfe0ef,
        64'h892a893f_e0ef842a,
        64'h899fe0ef_89aaec4e,
        64'hf04af426_f822fc06,
        64'he032e42e_7139b7f1,
        64'h00e83023_8f690008,
        64'h3703e314_8ee90785,
        64'h6314b15f_f06f6121,
        64'h863e69e2_854e7902,
        64'h74a270e2_744200c7,
        64'h9c63974e_00e58833,
        64'h00379713_47818d5d,
        64'h91011782_65a26602,
        64'h15028fc1_8d450109,
        64'h179b0105_151b8fff,
        64'he0ef84aa_905fe0ef,
        64'h892a90bf_e0ef842a,
        64'h911fe0ef_89aaec4e,
        64'hf04af426_f822fc06,
        64'he032e42e_7139b7f1,
        64'h00e83023_8f490008,
        64'h3703e314_8ec90785,
        64'h6314b8df_f06f6121,
        64'h863e69e2_854e7902,
        64'h74a270e2_744200c7,
        64'h9c63974e_00e58833,
        64'h00379713_47818d5d,
        64'h91011782_65a26602,
        64'h15028fc1_8d450109,
        64'h179b0105_151b977f,
        64'he0ef84aa_97dfe0ef,
        64'h892a983f_e0ef842a,
        64'h989fe0ef_89aaec4e,
        64'hf04af426_f822fc06,
        64'he032e42e_7139b7d1,
        64'h00e83023_02a75733,
        64'h00083703_e31402a6,
        64'hd6b30785_63144505,
        64'he111c0df_f06f6121,
        64'h863e69e2_854e7902,
        64'h74a270e2_744200c7,
        64'h9c63974e_00e58833,
        64'h00379713_47818d5d,
        64'h91011782_65a26602,
        64'h15028fc1_8d450109,
        64'h179b0105_151b9f7f,
        64'he0ef84aa_9fdfe0ef,
        64'h892aa03f_e0ef842a,
        64'ha09fe0ef_89aaec4e,
        64'hf04af426_f822fc06,
        64'he032e42e_7139b7e1,
        64'h00e83023_02a70733,
        64'h00083703_e31402a6,
        64'h86b30785_6314c89f,
        64'hf06f6121_863e69e2,
        64'h854e7902_74a270e2,
        64'h744200c7_9c63974e,
        64'h00e58833_00379713,
        64'h47818d5d_91011782,
        64'h65a26602_15028fc1,
        64'h8d450109_179b0105,
        64'h151ba73f_e0ef84aa,
        64'ha79fe0ef_892aa7ff,
        64'he0ef842a_a85fe0ef,
        64'h89aaec4e_f04af426,
        64'hf822fc06_e032e42e,
        64'h7139b7f1_00e83023,
        64'h8f090008_3703e314,
        64'h8e890785_6314d01f,
        64'hf06f6121_863e69e2,
        64'h854e7902_74a270e2,
        64'h744200c7_9c63974e,
        64'h00e58833_00379713,
        64'h47818d5d_91011782,
        64'h65a26602_15028fc1,
        64'h8d450109_179b0105,
        64'h151baebf_e0ef84aa,
        64'haf1fe0ef_892aaf7f,
        64'he0ef842a_afdfe0ef,
        64'h89aaec4e_f04af426,
        64'hf822fc06_e032e42e,
        64'h7139b7f1_00e83023,
        64'h8f290008_3703e314,
        64'h8ea90785_6314d79f,
        64'hf06f6121_863e69e2,
        64'h854e7902_74a270e2,
        64'h744200c7_9c63974e,
        64'h00e58833_00379713,
        64'h47818d5d_91011782,
        64'h65a26602_15028fc1,
        64'h8d450109_179b0105,
        64'h151bb63f_e0ef84aa,
        64'hb69fe0ef_892ab6ff,
        64'he0ef842a_b75fe0ef,
        64'h89aaec4e_f04af426,
        64'hf822fc06_e032e42e,
        64'h7139b7ad_0485a9df,
        64'hf0ef0007_c50397e2,
        64'h0039f793_0985aadf,
        64'hf0ef4521_ef8100ad,
        64'hb02300ac_b0238d41,
        64'h91011402_150201a4,
        64'h643300a9_6533010d,
        64'h1d1b0105_151b0344,
        64'hf7b3bcbf_e0ef892a,
        64'hbd1fe0ef_8d2abd7f,
        64'he0ef842a_bddfe0ef,
        64'he33ff06f_61657ae2,
        64'h85567b42_64e685da,
        64'h86266da2_6d426ce2,
        64'h7c027ba2_6a0669a6,
        64'h694670a6_74068bef,
        64'hd0ef03a5_05130000,
        64'h35170374_9b6300fb,
        64'h0cb300fa_8db30034,
        64'h97933a2c_0c130000,
        64'h3c179c4a_0a134981,
        64'hb3fff0ef_44818bb2,
        64'h8b2ee46e_e86aec66,
        64'he8caf0a2_f486f062,
        64'hf45ef85a_e4ceeca6,
        64'h02000513_8aaa6a05,
        64'hfc56e0d2_7159bfa5,
        64'h07a10585_80826125,
        64'h6ca26c42_6be27b02,
        64'h7aa27a42_79e26906,
        64'h64a66446_60e6557d,
        64'h938fd0ef_06c50513,
        64'h00003517_944fd0ef,
        64'h04050513_00003517,
        64'h058e02e6_0d6340e9,
        64'h87330035_9713c689,
        64'h873e8a85_63900085,
        64'h86b3bf5d_07a10485,
        64'h6398e398_40e98733,
        64'h00349713_c689873e,
        64'h8a850084_86b3a889,
        64'h450198af_d0ef0de5,
        64'h05130000_3517fd54,
        64'h17e30405_02b49b63,
        64'h458187ca_9a4fd0ef,
        64'h856285e6_9acfd0ef,
        64'h85520364_98634481,
        64'h87ca9baf_d0ef855e,
        64'h85e60004_0c9b9c6f,
        64'hd0ef8552_4ac10b6c,
        64'h0c130000_3c17fff9,
        64'h49930b2b_8b930000,
        64'h3b970aaa_0a130000,
        64'h3a179eaf_d0ef4401,
        64'h8b2ee466_e4a6ec86,
        64'he862ec5e_f05af456,
        64'hf852fc4e_e8a20be5,
        64'h05130000_3517892a,
        64'he0ca711d_bf5d0785,
        64'ha001a1af_d0ef0be5,
        64'h05130000_351785a2,
        64'h8626a2af_d0ef0a65,
        64'h05130000_35176090,
        64'h600c02e8_03636098,
        64'h00043803_80826105,
        64'h450164a2_644260e2,
        64'h00c79863_00d50433,
        64'h00d584b3_00379693,
        64'h4781e426_e822ec06,
        64'h1101bbbf_f06f8082,
        64'h45018082_45018082,
        64'h80828082_80824509,
        64'h80824509_80824509,
        64'hbff92605_20040413,
        64'h6622e37f_c0efe432,
        64'h852285b2_80826145,
        64'h450164e2_740270a2,
        64'h00961863_00c684bb,
        64'h842ef406_ec26f022,
        64'h71798082_45058082,
        64'h45058082_45058082,
        64'h01418d7d_640260a2,
        64'h95224080_07b3f57f,
        64'hf0efe406_952e842a,
        64'he0221141_a001cbbf,
        64'hf0ef4505_aecfd0ef,
        64'he4061325_05130000,
        64'h351785aa_862e86b2,
        64'h87361141_808202f5,
        64'h553347a9_b0002573,
        64'h80824501_80824501,
        64'h80820141_450160a2,
        64'hee5fc0ef_20000537,
        64'hb28fd0ef_e4061465,
        64'h05130000_35171141,
        64'h80828082_61056442,
        64'h60e28522_944ff0ef,
        64'h45816622_c509842a,
        64'hfd1ff0ef_e4328532,
        64'hec06e822_110102b5,
        64'h06338082_953e055e,
        64'h10d00513_e3089536,
        64'h00178693_00756513,
        64'h157d631c_c1c70713,
        64'h00004717_80824501,
        64'h80822405_0513000f,
        64'h4537a001_d69ff0ef,
        64'he4062501_11419002,
        64'h00000023_ee1ff0ef,
        64'h8522b781_1ac50513,
        64'h00003517_c5112501,
        64'hcb9fa0ef_4501e265,
        64'h85930000_35974605,
        64'hbfb91b25_05130000,
        64'h3517c511_2501b9af,
        64'hb0efa4a5_05130000,
        64'h4517be2f_d06f0141,
        64'h05850513_00003517,
        64'h60a26402_408005b3,
        64'hcf81439c_ca878793,
        64'h00004797_00054863,
        64'h842a90cf_90efca07,
        64'hab230000_4797cc07,
        64'ha1230000_4797e985,
        64'h05130000_0517c26f,
        64'hd0ef0825_05130000,
        64'h3517b7e1_20450513,
        64'h00003517_c5112501,
        64'hd9bfa0ef_ab450513,
        64'h00004517_20c58593,
        64'h00003597_4605c56f,
        64'hd0ef1fa5_05130000,
        64'h3517c62f_d06f0141,
        64'h60a26402_1ec50513,
        64'h00003517_c9112501,
        64'hd79fa0ef_e022e406,
        64'hd3050513_00004517,
        64'hef058593_00003597,
        64'h46051141_83020141,
        64'hbb858593_00002597,
        64'h60a26402_8322f140,
        64'h25730ff0_000f0000,
        64'h100fcb2f_d0efe406,
        64'h20850513_00003517,
        64'h842a85aa_e0221141,
        64'hbf95d687_a9230000,
        64'h47979c25_bf5d3200,
        64'h10ef854e_de7ff0ef,
        64'h00094503_993e0039,
        64'h79132327_87930000,
        64'h37970009_099b00c4,
        64'h591be05f_f0ef4521,
        64'hb775daf7_27230000,
        64'h47174785_d0cfd0ef,
        64'h23850513_00003517,
        64'h85a60496_75634632,
        64'hdca7a623_00004797,
        64'hc50d2501_814fb0ef,
        64'hba050513_00004517,
        64'h85ca8626_0074def7,
        64'h23230000_471757fd,
        64'h80826121_69e27902,
        64'h74a27442_70e2e0a7,
        64'ha1230000_4797c10d,
        64'h2501f3af_b0efbd65,
        64'h05130000_451702b7,
        64'h856384b2_842e892a,
        64'hec4efc06_f04af426,
        64'hf8227139_439ce2e7,
        64'h87930000_47978082,
        64'h610560e2_e9fff0ef,
        64'h00914503_ea7ff0ef,
        64'h00814503_f13ff0ef,
        64'hec06002c_11018082,
        64'h61456942_64e27402,
        64'h70a2fe94_10e3ec9f,
        64'hf0ef0091_4503ed1f,
        64'hf0ef3461_00814503,
        64'hf3fff0ef_0ff57513,
        64'h002c0089_553354e1,
        64'h03800413_892af406,
        64'he84aec26_f0227179,
        64'h80826145_694264e2,
        64'h740270a2_fe9410e3,
        64'hf0bff0ef_00914503,
        64'hf13ff0ef_34610081,
        64'h4503f81f_f0ef0ff5,
        64'h7513002c_0089553b,
        64'h54e14461_892af406,
        64'he84aec26_f0227179,
        64'h80826105_644260e2,
        64'hf43ff0ef_00914503,
        64'hf4bff0ef_00814503,
        64'hfb7ff0ef_0ff47513,
        64'h002cf5df_f0ef0091,
        64'h4503f65f_f0ef0081,
        64'h4503fd1f_f0efec06,
        64'h8121842a_002ce822,
        64'h11018082_00f58023,
        64'h00e580a3_0007c783,
        64'h00074703_97aa973e,
        64'h811100f5_7713d567,
        64'h87930000_2797b7f5,
        64'h0405fa5f_f0ef8082,
        64'h01416402_60a2e509,
        64'h00044503_842ae406,
        64'he0221141_808200e7,
        64'h88230200_071300e7,
        64'h8423fc70_071300e7,
        64'h8623470d_00078223,
        64'h00e78023_476d00e7,
        64'h8623f800_07130007,
        64'h82231000_07b78082,
        64'h00a70023_dfe50207,
        64'hf7930147_47831000,
        64'h07378082_02057513,
        64'h0147c503_100007b7,
        64'h80820005_45038082,
        64'h00b50023_80826105,
        64'h690264a2_644260e2,
        64'hf47dfa1f_f0ef4124,
        64'h0433854a_89260084,
        64'hf3638922_68048493,
        64'h842ae04a_ec06e822,
        64'h009894b7_e4261101,
        64'h80826105_690264a2,
        64'h644260e2_fe856ee3,
        64'hf45ff0ef_0405944a,
        64'h02855433_24040413,
        64'h000f4437_02a48533,
        64'h3e2000ef_892af63f,
        64'hf0ef84aa_e04ae426,
        64'he822ec06_11018082,
        64'h02a7d533_01419101,
        64'h15026402_60a202f4,
        64'h07b32407_8793000f,
        64'h47b74140_00ef842a,
        64'hf95ff0ef_e022e406,
        64'h11418082_610564a2,
        64'h8d0502a7_d5336442,
        64'h60e29101_150202f4,
        64'h07b33e80_07934400,
        64'h00ef842a_fc1ff0ef,
        64'h84aae426_e822ec06,
        64'h11018082_45018082,
        64'h01418d5d_91011782,
        64'h150260a2_1007e783,
        64'h10a7a223_10e1a023,
        64'h27051001_a70300e5,
        64'h7763878e_1041e703,
        64'h504000ef_e4061141,
        64'h8082cf3f_f06fc6e5,
        64'h85930000_45974611,
        64'hcb81e867_d7830000,
        64'h47978082_24010113,
        64'h22013903_22813483,
        64'h23013403_23813083,
        64'hf63ff0ef_8522002c,
        64'hea2ff0ef_e802c44a,
        64'h08282040_061385a6,
        64'he60ff0ef_22113c23,
        64'h00282180_06134581,
        64'h893284ae_842a2321,
        64'h30232291_34232281,
        64'h3823dc01_0113ebff,
        64'hf06f6145_05c170a2,
        64'h41907402_d8bff06f,
        64'h614570a2_65a27402,
        64'h85228a3f_d0efe42e,
        64'h59850513_00003517,
        64'h842a8b3f_d06f6145,
        64'h5c050513_00003517,
        64'h70a27402_02e78a63,
        64'h470d00e7_8e6301e1,
        64'h578300f1_0f230115,
        64'hc78300f1_0fa34709,
        64'h0105c783_f022f406,
        64'h71798082_61056902,
        64'h64a26442_60e2d49f,
        64'hf06f6105_690264a2,
        64'h60e26442_905fd0ef,
        64'h5e050513_00003517,
        64'h0087cf63_278d439c,
        64'hf7078793_00004797,
        64'hf6f71e23_00004717,
        64'h27850007_d783f8a7,
        64'h87930000_47972400,
        64'h00ef0200_0513d1bf,
        64'hf0ef4515_fa05d583,
        64'h00004597_256000ef,
        64'h4535e2bf_f0ef854a,
        64'hda858593_00004597,
        64'hdaa79923_00004797,
        64'h4611cf1f_f0effca5,
        64'h55030000_4517dca7,
        64'h93230000_4797d05f,
        64'hf0ef4511_dabff0ef,
        64'h00448513_ffc4059b,
        64'h06a79a63_25010024,
        64'hd783d21f_f0efffa5,
        64'h55030000_451708a7,
        64'h95632501_0004d783,
        64'hd37ff0ef_84ae450d,
        64'h892a08c7_df638432,
        64'h478de04a_e426ec06,
        64'he8221101_b79102f7,
        64'h15230000_47174785,
        64'heb1ff0ef_854ee2e5,
        64'h85930000_45974611,
        64'he2a79d23_00004797,
        64'hd77ff0ef_4501e4a7,
        64'h93230000_4797d85f,
        64'hf0ef06f7_35230000,
        64'h471706f7_35230000,
        64'h47174511_07e20810,
        64'h0793a1bf_d0ef6d65,
        64'h05130000_3517858a,
        64'h43900827_87930000,
        64'h4797df2f_f0ef850a,
        64'h85a2dfaf_f0ef850a,
        64'h6f058593_00003597,
        64'h00f70963_02f00793,
        64'h01294703_deaff0ef,
        64'h850a4c25_85930000,
        64'h3597863f_f0ef850a,
        64'h45811000_0613b755,
        64'h0cf72423_00004717,
        64'h20000793_80826155,
        64'h69b26952_64f27412,
        64'h70b2a8bf_d0ef71e5,
        64'h05130000_351700a4,
        64'h05b3f24f_f0ef5065,
        64'h05130000_3517842a,
        64'hf32ff0ef_852204a7,
        64'hf2630ff0_07939526,
        64'hf42ff0ef_52450513,
        64'h00003517_84aaf50f,
        64'hf0ef8522_12a7a223,
        64'h00004797_04e7ee63,
        64'h1ff00793_fff5071b,
        64'he93ff0ef_95260505,
        64'hf72ff0ef_852600a4,
        64'h04b30505_f7eff0ef,
        64'h892eea4a_ee26f606,
        64'h852289aa_e64e0125,
        64'h8413f222_71698082,
        64'h45018082_01416402,
        64'h60a2557d_00850363,
        64'h878fa0ef_8432e406,
        64'he0221141_6680006f,
        64'h610564a2_60e26442,
        64'hb39fd06f_61057ae5,
        64'h05130000_351740a0,
        64'h05b364a2_60e26442,
        64'h00055e63_857f90ef,
        64'hef650513_00000517,
        64'hb61fd0ef_7bc50513,
        64'h00003517_b6dfd0ef,
        64'h7b050513_00003517,
        64'h862286aa_608ce63f,
        64'hc0ef85a2_6088b87f,
        64'hd0ef85a2_9c11ec06,
        64'h7b850513_00003517,
        64'h6380e822_60901fe4,
        64'h84930000_4497e426,
        64'h21078793_00004797,
        64'h11018082_610564a2,
        64'h6442e00c_95a660e2,
        64'h600ca15f_f0efec06,
        64'h600885aa_84ae862e,
        64'he42623a4_04130000,
        64'h4417e822_11018082,
        64'h24f73423_00004717,
        64'h24f73423_00004717,
        64'h07e20810_07935000,
        64'h006f0305_05130141,
        64'h60a26402_02a4753b,
        64'h4529fe7f_f0ef357d,
        64'h02b455bb_45a900b7,
        64'hf86347a5_00a04563,
        64'h842ee406_e0221141,
        64'hbff90505_fd07879b,
        64'h9fb902f5_87bb00d6,
        64'h67630ff6_f693fd07,
        64'h069b8082_853ee319,
        64'h00054703_45a94625,
        64'h4781aa5f_f06f95be,
        64'h92011602_91811582,
        64'h639c2c27_87930000,
        64'h47978082_014100e1,
        64'h550300a1_07238121,
        64'h00a107a3_1141fa5f,
        64'hf06f4581_d7dff06f,
        64'h01410505_45814629,
        64'h60a26402_f77d8b11,
        64'h00074703_973e0005,
        64'h4703fea4_7ae3157d,
        64'h80820141_557d6402,
        64'h60a2e719_8b110007,
        64'h4703973e_fff58513,
        64'he3078793_00002797,
        64'hfff5c703_00a405b3,
        64'h95bff0ef_e589842a,
        64'he406e022_1141bfd5,
        64'h0789bff1_052a052a,
        64'hb7e9e01c_078d00e6,
        64'h98630420_07130027,
        64'hc683fce6_9fe3052a,
        64'h06900713_0017c683,
        64'hfed716e3_06b00693,
        64'h02d70763_04d00693,
        64'h80820141_640260a2,
        64'h02d70e63_04700693,
        64'h00e6ea63_02d70463,
        64'h0007c703_04b00693,
        64'h601cf87f_f0ef842e,
        64'he406e022_1141b7e1,
        64'he008b7cd_fc97879b,
        64'h0ff7f793_fe07079b,
        64'hc6098a09_b7d196be,
        64'h050502d5_86b3feb7,
        64'hf4e3fd07_879b0008,
        64'h8b630046_78938082,
        64'h61058536_644260e2,
        64'hec050008_98630446,
        64'h78930006_460300f8,
        64'h06330007_079b0005,
        64'h4703f0a8_08130000,
        64'h28174681_00c16583,
        64'he0fff0ef_c632ec06,
        64'h006c842e_e8221101,
        64'hbfd50789_bff1052a,
        64'h052ab7e9_e01c078d,
        64'h00e69863_04200713,
        64'h0027c683_fce69fe3,
        64'h052a0690_07130017,
        64'hc683fed7_16e306b0,
        64'h069302d7_076304d0,
        64'h06938082_01416402,
        64'h60a202d7_0e630470,
        64'h069300e6_ea6302d7,
        64'h04630007_c70304b0,
        64'h0693601c_f0dff0ef,
        64'h842ee406_e0221141,
        64'h80820141_40a00533,
        64'h60a2f23f_f0efe406,
        64'h05051141_f2dff06f,
        64'h00e68463_02d00713,
        64'h00054683_b7e94501,
        64'he088fcf7_18e347a9,
        64'hfd279be3_07858f81,
        64'hcb010007_c703fe87,
        64'h82e367e2_f5dff0ef,
        64'h8522082c_892a862e,
        64'h80826121_790274a2,
        64'h744270e2_5529e901,
        64'h65a2b0df_f0ef84b2,
        64'h842ae42e_00063023,
        64'hf04afc06_f426f822,
        64'h7139b7e1_e008b7cd,
        64'hfc97879b_0ff7f793,
        64'hfe07079b_c6098a09,
        64'hb7d196be_050502d5,
        64'h86b3feb7_f4e3fd07,
        64'h879b0008_8b630046,
        64'h78938082_61058536,
        64'h644260e2_ec050008,
        64'h98630446_78930006,
        64'h460300f8_06330007,
        64'h079b0005_470305e8,
        64'h08130000_28174681,
        64'h00c16583_f63ff0ef,
        64'hc632ec06_006c842e,
        64'he8221101_bf6d47a9,
        64'hbf7d47a1_80820509,
        64'h00e79363_07800713,
        64'h0ff7f793_0207879b,
        64'hc7098b05_00074703,
        64'h973e0a27_07130000,
        64'h27170015_478302f7,
        64'h16630300_07930005,
        64'h470302f7_1c6347c1,
        64'h4198c19c_47c1c3b1,
        64'h0447f793_0007c783,
        64'h97ba0025_470304d7,
        64'h1b630780_06930ff7,
        64'h77130207_071bc689,
        64'h8a850006_c68300e7,
        64'h86b30f27_87930000,
        64'h27970015_470308f7,
        64'h11630300_07930005,
        64'h4703e7a9_419cb7f1,
        64'h377d87aa_bfa5fef5,
        64'h1be30785_f8b712e3,
        64'h0007c703_00d80a63,
        64'h00878513_0007b803,
        64'hbfcd367d_0785f8b7,
        64'h1fe30007_c703d24d,
        64'h8a1deb11_87aa2701,
        64'h8edd0036_57130207,
        64'h96938fd9_01071793,
        64'h00b7e733_00859793,
        64'h8e1d953e_93810207,
        64'h1793faf5_078536fd,
        64'hfcb81ce3_0007c803,
        64'h87aa0007_069b40e7,
        64'h873b47a1_c31d0075,
        64'h7713b7f5_367d0785,
        64'hfeb71ce3_0007c703,
        64'h8082853e_4781e601,
        64'h87aa2601_00c7ef63,
        64'h0ff5f593_47c1b7ed,
        64'h853efeb7_0be30015,
        64'h07930005_47038082,
        64'h450100c5_14630ff5,
        64'hf593962a_bfe90405,
        64'hd175f8bf_f0ef397d,
        64'h852285ce_86268082,
        64'h614569a2_694264e2,
        64'h740270a2_85224401,
        64'h00995b63_0005091b,
        64'hd13ff0ef_8522c889,
        64'h0005049b_d1fff0ef,
        64'h89aee84a_f406e44e,
        64'hec26852e_842af022,
        64'h7179bfc5_0505feb7,
        64'h8de30005_47838082,
        64'h00c51363_962ab7dd,
        64'h05850505_fbed9f99,
        64'h0005c703_00054783,
        64'h8082853e_478100c5,
        64'h1563962a_b7fd00f6,
        64'h802316fd_0005c783,
        64'h15fdd7e5_00e587b3,
        64'h40b60733_00c506b3,
        64'h95b28082_01416402,
        64'h60a28522_f57ff0ef,
        64'h00a5e963_842ae406,
        64'he0221141_80826145,
        64'h64e26942_85267402,
        64'h70a20004_0023f79f,
        64'hf0ef944a_864a8522,
        64'hfff60913_00c56463,
        64'h6582892a_ce1184aa,
        64'h6622dcdf_f0efe02e,
        64'he84af406_e432ec26,
        64'h852e842a_f0227179,
        64'hbf65fee7_8fa30785,
        64'hfff5c703_0585bfe1,
        64'h469d00c5_08b387aa,
        64'h872ebfc1_00e507b3,
        64'h963e95ba_070e02f7,
        64'h07b357e1_00365713,
        64'hff06e8e3_40f88833,
        64'hff07bc23_07a1ff87,
        64'h38030721_808202c7,
        64'h9e63963e_87aacb9d,
        64'h8b9d00a5_e7b300b5,
        64'h0a63bf6d_feb78fa3,
        64'h0785bfe1_fef73c23,
        64'h0721bfd1_0ff5f693,
        64'h4725bfc1_963a97aa,
        64'h078e02e7_87335761,
        64'h00365793_0106ef63,
        64'h40e88833_469d00c5,
        64'h08b3872a_ff6d377d,
        64'h8fd507a2_808204c7,
        64'h9063963e_87aacb9d,
        64'h00757793_80824501,
        64'hb7e50789_00d780a3,
        64'h00e78023_8082e311,
        64'h0017c703_ce810007,
        64'hc68387aa_cf990005,
        64'h4783c11d_80826105,
        64'h64a28526_644260e2,
        64'he0080505_00050023,
        64'hc501f73f_f0ef8526,
        64'h842ac891_e822ec06,
        64'h6104e426_1101bfd9,
        64'h6aa7b023_00004797,
        64'h05050005_0023c781,
        64'h00054783_c519f9ff,
        64'hf0ef8522_85a68082,
        64'h610564a2_644260e2,
        64'h85224401_6c07b623,
        64'h00004797_ef810004,
        64'h4783942a_f9dff0ef,
        64'h85a68522_cc116380,
        64'h6e878793_00004797,
        64'he519842a_84aeec06,
        64'he426e822_1101bfd5,
        64'h87aeb7e5_0505fafd,
        64'h0007c683_0785fee6,
        64'h8fe38082_4501eb19,
        64'h00054703_bff90785,
        64'hbfd5872e_8082fe08,
        64'h1be30007_48030705,
        64'h00c80a63_8082ea11,
        64'h40d78533_0007c603,
        64'h87aa86aa_bfcd872e,
        64'hb7d50785_fe081be3,
        64'h00074803_0705fed8,
        64'h0fe38082_ea9940c7,
        64'h85330007_c68387aa,
        64'h862ab7fd_07858082,
        64'h40a78533_e7010007,
        64'hc70300b7_856387aa,
        64'h95aa8082_61056442,
        64'h60e24501_fe857be3,
        64'h157d00b7_86630005,
        64'h47830ff5_f5939522,
        64'h65a2fe5f_f0efec06,
        64'h842ae42e_e8221101,
        64'hbfcd0785_808240a7,
        64'h8533e701_0007c703,
        64'h87aabfcd_0505dffd,
        64'h808200b7_93630005,
        64'h47830ff5_f5938082,
        64'h4501bfcd_0505c399,
        64'h808200b7_93630005,
        64'h47830ff5_f5938082,
        64'h853eff79_0505e399,
        64'h4187d79b_0187979b,
        64'h40f707bb_fff5c783,
        64'h00054703_0585a839,
        64'h478100c5_9463962e,
        64'h8082853e_f37d0505,
        64'he3994187_d79b0187,
        64'h979b40f7_07bbfff5,
        64'hc7830005_47030585,
        64'hb7cd87ba_80820007,
        64'h80a300c7_15638082,
        64'he291fed7_0fa30017,
        64'h8713fff5_c6830585,
        64'h963efb7d_00178693,
        64'h0007c703_87b68082,
        64'he21987aa_b7d587b6,
        64'h8082fb75_fee78fa3,
        64'h0785fff5_c7030585,
        64'heb090017_86930007,
        64'hc70387aa_8082fb65,
        64'hfee78fa3_0785fff5,
        64'hc7030585_00c78963,
        64'h87aa962a_8082fb75,
        64'hfee78fa3_0785fff5,
        64'hc7030585_87aa8082,
        64'h01416402_60a28d41,
        64'h15029001_fd1ff0ef,
        64'h14020005_041bfdbf,
        64'hf0efe022_e4061141,
        64'h80820141_25016402,
        64'h60a28d41_0105151b,
        64'hfe9ff0ef_842afeff,
        64'hf0efe022_e4061141,
        64'hfc3ff06f_8ec50513,
        64'h00005517_80822501,
        64'h8d5d00f7_17bb40f0,
        64'h07b300f7_553b93ed,
        64'h836d8f3d_0127d713,
        64'he1189736_00176713,
        64'h02d786b3_65186294,
        64'h611c6b26_86930000,
        64'h46971bc0_106f8082,
        64'h61056902_64a26442,
        64'h60e28522_e99ff0ef,
        64'h10f40023_0247c783,
        64'h85220ea4_2e23681c,
        64'h18f43423_2ae78793,
        64'h00001797_18f43023,
        64'h2be78793_00001797,
        64'h16f43c23_91c78793,
        64'hfffff797_e65ff0ef,
        64'h04052823_03253023,
        64'he90410f5_02a34785,
        64'h0ef52c23_4799c57c,
        64'h57fdcd21_842a2000,
        64'h10ef4505_1c000593,
        64'h84aa892e_c7ad639c,
        64'hc7bd651c_cbad511c,
        64'hcbbd4d5c_cfad4401,
        64'h4d1cc141_4401e04a,
        64'he426ec06_e8221101,
        64'hb7716000_32a010ef,
        64'h79850513_00003517,
        64'h01a98863_da4fe0ef,
        64'h856685e2_00978e63,
        64'h601cdb2f_e0ef855e,
        64'h85ca0009_0663dbef,
        64'he0ef638c_855a0fc4,
        64'h2603681c_89560007,
        64'hc3638952_4c1cc791,
        64'h4901541c_ddcfe06f,
        64'h612537a5_05130000,
        64'h45176d02_6ca26c42,
        64'h6be27b02_7aa27a42,
        64'h79e26906_64a660e6,
        64'h64460294_15634d29,
        64'h810c8c93_00004c97,
        64'h00050c1b_22cb8b93,
        64'h00004b97_22cb0b13,
        64'h00004b17_224a8a93,
        64'h00004a97_234a0a13,
        64'h00004a17_89aae0ca,
        64'hec86e06a_e466e862,
        64'hec5ef05a_f456f852,
        64'hfc4e6080_e8a2a764,
        64'h84930000_5497e4a6,
        64'h711d8082_e308e518,
        64'he11ce788_6798a8e7,
        64'h87930000_5797e508,
        64'h80829207_a5230000,
        64'h5797e79c_e39caa67,
        64'h87930000_5797b7d5,
        64'h6000a9cf_f0ef8522,
        64'hc78119a4_47838082,
        64'h610564a2_644260e2,
        64'h00941763_84beec06,
        64'he4266380_e822ad67,
        64'h87930000_57971101,
        64'h80824388_97478793,
        64'h00005797_80820f85,
        64'h05138082_c3980015,
        64'h071b4388_98c78793,
        64'h00005797_bfd55535,
        64'h80826105_64a26442,
        64'h60e2e080_0f840413,
        64'he501cf0f_f0ef842a,
        64'hcd09f7df_f0ef84ae,
        64'he822ec06_e4261101,
        64'hbfcdf840_0513bfe5,
        64'h45018082_610560e2,
        64'h5535eb3f_e06f6105,
        64'h60e200f7_0c630ff0,
        64'h07930815_470302b7,
        64'h006365a2_10354703,
        64'hc105fbdf_f0efe42e,
        64'hec061101_41488082,
        64'h853ebfd1_87b600a6,
        64'h04630fc7_a6038082,
        64'h0141853e_478160a2,
        64'hf60fe0ef_e4063465,
        64'h05130000_451785aa,
        64'h114102e7_90636394,
        64'h631cba27_07130000,
        64'h57178082_45018082,
        64'h01414501_640260a2,
        64'h0dc000ef_13e000ef,
        64'h02c00513_fc5ff0ef,
        64'h85220005_5563aeef,
        64'he0ef8522_12a000ef,
        64'hbcf72a23_00005717,
        64'h842ae406_e0224785,
        64'h1141ef9d_439cbea7,
        64'h87930000_57978082,
        64'h18b50d23_8082557d,
        64'h8082557d_80824501,
        64'hc56ce54f_f06ffa10,
        64'h0413f0ef_f06f2006,
        64'h061b4001_0637f0a6,
        64'h09634505_f0c54363,
        64'h8ca602e3_45098a3d,
        64'h01a6d61b_f2c51a63,
        64'h40000637_06bba423,
        64'h06eba223_06fba023,
        64'h04dbae23_018ba503,
        64'h45e64756_47c646b6,
        64'hea051163_842a93bf,
        64'he0efc4be_855e0107,
        64'h979b008c_460107cb,
        64'hd783c2be_479d04f1,
        64'h102347a5_06fb9e23,
        64'h04e15783_0007d663,
        64'h018ba783_ec051b63,
        64'h842a96ff_e0efc2be,
        64'h47d5855e_c4be0107,
        64'h979b008c_460107cb,
        64'hd78304f1_1023478d,
        64'h6da000ef_06cb8513,
        64'h00ec4641_bf6d1187,
        64'h2583974e_83790207,
        64'h9713fcfc_65e34581,
        64'hb7c9f521_d31fe0ef,
        64'h855e4585_0b700613,
        64'h0ff6f693_bb91fd31,
        64'h9fdfe0ef_855ecb0f,
        64'hf0ef855e_460118fb,
        64'hae2308bb_a2230017,
        64'hb79317ed_088ba583,
        64'hef8d1afb_a823409c,
        64'he79d0046_f7930089,
        64'h2683f941_808ff0ef,
        64'h855e408c_933fe0ef,
        64'h855e02eb_aa230017,
        64'hb71341b7_87b301a7,
        64'h86634711_00d78963,
        64'h47214000_06b70009,
        64'h2783bb6d_925fe0ef,
        64'h39850513_00004517,
        64'hf7649fe3_04a1fb99,
        64'h11e30931_973fe0ef,
        64'h855e035b_aa2308fb,
        64'ha223180b_ae231a0b,
        64'ha823088b_a783ddbf,
        64'he0ef855e_45850b70,
        64'h06134681_c131debf,
        64'he0ef855e_0fb6f693,
        64'h45850b70_06130089,
        64'h4683c3a1_8ff900fa,
        64'h77b30009_270340dc,
        64'h04f71863_0017b793,
        64'h17ed0049_4703409c,
        64'h10000db7_20000d37,
        64'hf9890913_00003917,
        64'hcbb52781_00fa77b3,
        64'h00fa97bb_409cfeac,
        64'h8c930000_3c974c2d,
        64'hfb8b0b13_00003b17,
        64'h4a85db4f_f0effa64,
        64'h84930000_349700fa,
        64'h7a33855e_4601088b,
        64'ha583044b_a783040b,
        64'haa0304fb_a02300c7,
        64'he793040b_a783c799,
        64'h8b8504eb_a0230107,
        64'h6713040b_a70304eb,
        64'ha0230217_071bc689,
        64'h00c7f693_ce910027,
        64'hf6931adb_a42303f7,
        64'hf6930c46_c78304fb,
        64'ha0230017_079b7000,
        64'h0737bb95_4c450513,
        64'h00004517_e691ecf7,
        64'h6ce31a0b_b6834004,
        64'h07b704fb_a0232785,
        64'h100007b7_b8d102fb,
        64'ha4234785_7e4010ef,
        64'h8526a3ff_e0ef8a3d,
        64'h8abd0146_561b0106,
        64'h569b0624_85135465,
        64'h85930000_4597074b,
        64'ha603a5ff_e0ef04d4,
        64'h851354a5_85930000,
        64'h45972681_0ff77713,
        64'h0ff87813_0ff7f793,
        64'h0188569b_0108571b,
        64'h0088579b_06cbc603,
        64'h077bc883_070ba803,
        64'ha95fe0ef_fef53623,
        64'h02450513_56c58593,
        64'h00004597_84aa06fb,
        64'hc603074b_d68307ab,
        64'hd70302c7_d7b3ed10,
        64'h92010a8b_b783d11c,
        64'h9fb90712_00e03733,
        64'h8f750207_161376c1,
        64'h9fb5068e_00d036b3,
        64'h8ef9f006_8693ff01,
        64'h06b79fb5_068a00d0,
        64'h36b38ef9_0f068693,
        64'hf0f0f6b7_9fb500f0,
        64'h37b30686_00d036b3,
        64'h27818ef9_8ff9ccc6,
        64'h8693aaa7_8793cccc,
        64'hd6b7aaaa_b7b708cb,
        64'ha7030005_06230005,
        64'h15234840_00ef855e,
        64'h08fba823_08fba623,
        64'h20000793_c79919cb,
        64'ha7831afb_aa231b0b,
        64'ha7830adb_a2230afb,
        64'ha02302d6_06bb02f7,
        64'h57bb8a8d_0106d69b,
        64'h02e6073b_3e800613,
        64'hc305c38d_03f77713,
        64'h27810126_d71b8fd1,
        64'h0186d61b_8ff917fd,
        64'h67c100cc_a68308fb,
        64'hae230087_171b1487,
        64'ha78397b6_078a0f66,
        64'h86930000_369704d6,
        64'h1c638003_06b7018b,
        64'ha60300f6_f8638bbd,
        64'h00c7579b_46a5008c,
        64'ha703fdb5_9ee3fefd,
        64'hae238fd9_8ff58f51,
        64'h0087d79b_8e690087,
        64'h961b8f51_0187971b,
        64'h0187d61b_0d91000d,
        64'ha783f006_869300ff,
        64'h0537040d_859366c1,
        64'hb5451187_2583974e,
        64'h83790207_9713eaf7,
        64'h68e34581_472db35d,
        64'h04fba023_00876793,
        64'hda06d9e3_040ba703,
        64'h02e79693_8fd18ff5,
        64'h0087d79b_0087961b,
        64'hf0068693_66c144dc,
        64'hfbe18b85_83a54cdc,
        64'hd0051ce3_d61fe0ef,
        64'hdc3ef84a_f426c556,
        64'h855e010c_04000793,
        64'h1030c33e_47d508f1,
        64'h10234799_020a0863,
        64'h3a7d0905_3ac54a15,
        64'h98811902_01000ab7,
        64'h0ff10493_4905bbc5,
        64'h80030737_de075ee3,
        64'h03079713_00ebac23,
        64'h80020737_b519a007,
        64'h071b8001_1737b61d,
        64'hdf400413_cbdfe0ef,
        64'h73050513_00004517,
        64'he6f49fe3_2a478793,
        64'h00003797_04a1eafa,
        64'h94e347a1_0a918c9f,
        64'hf0ef855e_84058593,
        64'h4601180b_ae23096b,
        64'ha2231afb_a823017d,
        64'h85b74785_f3ed37fd,
        64'h670267a2_0e050c63,
        64'he0dfe0ef_e03ac93a,
        64'he552e16e_e43e855e,
        64'h110c0110_04000713,
        64'h4791d502_d33a0af1,
        64'h102347b5_6702e915,
        64'he35fe0ef_d53ee03a,
        64'hd33a8cee_855e110c,
        64'h0107979b_46014755,
        64'h07cbd783_0af11023,
        64'h03700793_fe07fd93,
        64'h0ff10793_947ff0ef,
        64'h855e4601_18fbae23,
        64'h08bba223_0017b793,
        64'h17ed088b_a5831407,
        64'h9a631afb_a823409c,
        64'h09b79463_8bbd010c,
        64'h4783e941_e91fe0ef,
        64'hc93ee552_e162855e,
        64'h110c0400_07930110,
        64'hd53e00fd_e7b317c1,
        64'h2d818100_07b7d33e,
        64'h47d50af1_10234799,
        64'h4d850ce7_9163470d,
        64'h01a78663_409cdfdf,
        64'he0ef855e_02fbaa23,
        64'h001cb793_40fc8cb3,
        64'h100007b7_00ec8863,
        64'h47912000_073700ec,
        64'h8d6347a1_40000737,
        64'h0e051c63_8daa971f,
        64'hf0ef855e_0015b593,
        64'h40bc85b3_100005b7,
        64'h00fc8863_45912000,
        64'h07b700fc_8d6345a1,
        64'h400007b7_14078163,
        64'h0197f7b3_00f977b3,
        64'h40dc0007_ac8397d6,
        64'h109c840b_0b1b4a81,
        64'h017d8b37_16078563,
        64'h278100f9_77b300e7,
        64'h97bb4785_40980a05,
        64'hfe07fc13_83f97913,
        64'h0ff10793_00f97933,
        64'h42848493_00003497,
        64'h020d1a13_044ba783,
        64'hf0be4d05_040ba903,
        64'h639c03a7_87930000,
        64'h57971ef7_18638001,
        64'h07b7018b_a70304fb,
        64'ha0238fd9_20000737,
        64'h040ba783_00075963,
        64'h02d79713_00ebac23,
        64'h80010737_20d70263,
        64'h46892127_00638b3d,
        64'h0187d71b_04ebac23,
        64'h8f558f71_8ecd0087,
        64'h571b8de9_0087159b,
        64'h8ecd0187_169b0187,
        64'h559b40d8_04fbaa23,
        64'h27818fd5_8ef1f007,
        64'h06138fd1_67410087,
        64'h569b8e69_8fd50087,
        64'h161b0187_179b0187,
        64'h569b00ff_05374098,
        64'hb5558b1d_938100f7,
        64'h571b1782_8fd501e7,
        64'h569b8ff5_0027979b,
        64'h16f16685_b54d08bb,
        64'ha82300b5_15bb89bd,
        64'h0165d59b_bd994003,
        64'h0637a7a9_40020637,
        64'hbb45842a_fe0a16e3,
        64'h3a7dc131_850ff0ef,
        64'hd05aec56_e826855e,
        64'h108c0810_4b210a85,
        64'h4a11d482_06f11023,
        64'h98810209_1a930330,
        64'h07930bf1_04934905,
        64'hd2caed05_880ff0ef,
        64'hd4bed2ca_855e0107,
        64'h979b108c_460107cb,
        64'hd78306f1_10230370,
        64'h079304fb_a0232789,
        64'h100007b7_54075a63,
        64'h018ba703_e0051fe3,
        64'h842affbf_e0ef855e,
        64'h00b54583_0f7000ef,
        64'h855ee205_1ae3842a,
        64'hc9aff0ef_855e08fb,
        64'h80a357fd_08fbaa23,
        64'h4785e405_16e3842a,
        64'h8e4ff0ef_c4bec2ca,
        64'h855e008c_0107979b,
        64'h46014955_07cbd783,
        64'h04f11023_479d902f,
        64'hf0efc282_c4be04e1,
        64'h1023855e_008c4601,
        64'h0107979b_471100e7,
        64'h8e63577d_04cba783,
        64'hc21508fb_a82300e7,
        64'hf4632000_0793090b,
        64'ha70308fb_a6230107,
        64'hd4632000_07930afb,
        64'hb8230e0b_b0230c0b,
        64'hbc230c0b_b8230c0b,
        64'hb4230c0b_b0230a0b,
        64'hbc230307_87b300e7,
        64'h97b30709_07854721,
        64'h93811782_8fd98ff5,
        64'h0107571b_003f06b7,
        64'h0107979b_14068e63,
        64'h02cba683_090ba823,
        64'h1408dc63_090ba623,
        64'h00d5183b_8abd0107,
        64'hd69b08db_a22308db,
        64'ha42304cb_a823180b,
        64'hae231a0b_a8238a05,
        64'h00c7d61b_02d606bb,
        64'h018ba883_45051086,
        64'ha6830f86_460396ce,
        64'h964e068a_8a3d60e9,
        64'h89930000_39978a9d,
        64'h0036d61b_00cbac23,
        64'h4006061b_40010637,
        64'ha0294004_06370ea6,
        64'h1ee34511_1aa60f63,
        64'h450dbf05_06fb9e23,
        64'h478502fb_a6238b85,
        64'h41e7d79b_048ba783,
        64'h00fbac23_400007b7,
        64'hbfe91d70_10ef0640,
        64'h051312a9_6ee31490,
        64'h10ef8526_0007cc63,
        64'h048ba783_f155842a,
        64'hb36ff0ef_855e4585,
        64'h3e800913_90810205,
        64'h149316d0_10ef4501,
        64'hb16ff0ef_855e0407,
        64'hc163180b_8c23048b,
        64'ha7838082_615d6db6,
        64'h6d566cf6_7c167bb6,
        64'h7b567af6_6a1a69ba,
        64'h695a64fa_741a70ba,
        64'h8522d55d_842ad99f,
        64'hf0ef855e_a031020b,
        64'ha423f4fd_34fd1005,
        64'h03e3842a_aa0ff0ef,
        64'h855e008c_46014495,
        64'hcf818b85_1b8ba783,
        64'h120500e3_842aabaf,
        64'hf0efc482_c2be855e,
        64'h008c479d_460104f1,
        64'h10234789_e7b5180b,
        64'h8ca3198b_c783c7b1,
        64'h199bc783_1ff010ef,
        64'h45018baa_e3b54401,
        64'he6eeeaea_eee6f2e2,
        64'hf6defada_fed6e352,
        64'he74eeb4a_ef26f706,
        64'hf3227161_551cb585,
        64'h84aab595_fa100493,
        64'ha10ff0ef_c5450513,
        64'h00005517_d965c1cf,
        64'hf0ef8522_4585bfd1,
        64'h18f40c23_47850007,
        64'hd663443c_ed09c34f,
        64'hf0ef8522_4581c04f,
        64'hf0ef8522_02f51f63,
        64'hf9200793_b55d18f4,
        64'h0ca34785_06041e23,
        64'hd45c8b85_41e7d79b,
        64'hc43ccc18_80010737,
        64'h00e68563_80020737,
        64'h4c14bf45_331010ef,
        64'h3e800513_06090863,
        64'h397d0007_ca6347b2,
        64'hed1db8ef_f0ef8522,
        64'h858a4601_c43e0197,
        64'he7b30187_1563c43e,
        64'h0177f7b3_c25a4bdc,
        64'h01511023_4c18681c,
        64'he13dbb6f_f0efc402,
        64'hc2520131_10238522,
        64'h858a4601_40000cb7,
        64'h80020c37_00ff8bb7,
        64'h4b050290_0a934a55,
        64'h03700993_3e900913,
        64'hcc1c8002_07b700f7,
        64'h15630aa0_079300c1,
        64'h4703e911_bf8ff0ef,
        64'hc23ec43a_8522858a,
        64'h460147d5_0aa00713,
        64'he3991aa0_07138ff9,
        64'h4bdc00ff_8737681c,
        64'h00f11023_47a10005,
        64'h05a345d0_00ef8522,
        64'hf14984aa_cf2ff0ef,
        64'h8522f1df_f0ef8522,
        64'h45814601_b72ff0ef,
        64'h8522d85c_478508f4,
        64'h22231a04_28231804,
        64'h2e230884_2783f945,
        64'h84aa9782_6b9c679c,
        64'h8522681c_421010ef,
        64'h7d000513_ba2ff0ef,
        64'h85220204_2c2302f4,
        64'h08234785_1af42c23,
        64'h478df93f_f0eff3e5,
        64'h4481541c_80826109,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e674a6,
        64'h79068526_744670e6,
        64'hf8500493_bacff0ef,
        64'hdd850513_00005517,
        64'h02042423_eb8d6b9c,
        64'h679c681c_c509f11f,
        64'hf0ef842a_c17c8fd9,
        64'hf466f862_fc5ee0da,
        64'he4d6e8d2_eccef0ca,
        64'hf4a6fc86_f8a2070d,
        64'h4b9c7119_10000737,
        64'h691c8082_8082c2cf,
        64'hf06f02c5_0823dd0c,
        64'h0007059b_00e7f463,
        64'h85be2781_4f1887ae,
        64'h00f5f363_4f5c6918,
        64'hee09b7cd_c402fef4,
        64'h14e34785_80826121,
        64'h790274a2_744270e2,
        64'hd34ff0ef_8526858a,
        64'h4601c43e_478900f4,
        64'h1f634791_c24a00f1,
        64'h10234799_ed19d52f,
        64'hf0efc43e_c24a8526,
        64'h858a4601_0107979b,
        64'h4955842e_07c4d783,
        64'h00f11023_03700793,
        64'h04f59263_55294785,
        64'h00f58663_84aa4791,
        64'hf04af822_fc06f426,
        64'h71398082_01416402,
        64'h60a24505_83020141,
        64'h60a26402_85220003,
        64'h07630187_b303679c,
        64'h681c0005_5e63810f,
        64'hf0ef842a_e406e022,
        64'h1141b32d_dd79842a,
        64'h945ff0ef_854a4585,
        64'h0a700613_86cebb3d,
        64'h842a957f_f0ef854a,
        64'h458509b0_06134685,
        64'h01379b63_0a7a4783,
        64'hd4fb0de3_4785ed19,
        64'h975ff0ef_854a4585,
        64'h09c00613_86defdb4,
        64'h98e30c11_0ff4f493,
        64'h248dffac_90e30ffa,
        64'hfa932ca1_2a85e139,
        64'h99dff0ef_854a0ff6,
        64'hf6930196_d6bb4585,
        64'h8656000c_26834c81,
        64'h8aa609b0_0d934d61,
        64'hffa492e3_2ca10ff4,
        64'hf4932485_e9359cbf,
        64'hf0ef854a_45858626,
        64'h0ff6f693_019ad6bb,
        64'h08f00d13_4c81ffb4,
        64'h92e32d21_0ff4f493,
        64'h2485ed49_9f1ff0ef,
        64'h854a4585_86260ff6,
        64'hf69301ac_d6bb08c0,
        64'h0d934d01_08800493,
        64'h08f92a23_00a7979b,
        64'h0e0a4783_0afa07a3,
        64'h4785e569_a21ff0ef,
        64'h854a4585_0af00613,
        64'h4685e395_8b850afa,
        64'h4783e20b_02e3b51d,
        64'h547ddbaf_f0effc65,
        64'h05130000_5517cb89,
        64'h8b8509ba_4783bfd1,
        64'h00f9f9b3_fff7c793,
        64'hb5913700_20eff965,
        64'h05130000_5517ef89,
        64'h8b850a6a_478302d9,
        64'h8263fcc5_92e3872e,
        64'h0ff9f993_00f9e9b3,
        64'hc70d4189_d99b4187,
        64'hd79b8b05_0189999b,
        64'h0187979b_0027571b,
        64'h00b517bb_02080463,
        64'h00187813_0017581b,
        64'h4b189726_070e0017,
        64'h059b4611_45054701,
        64'h0016e993_c3990fe6,
        64'hf9938b89_c71989b6,
        64'h0017f713_0a7a4683,
        64'h0084c783_b5c1e56f,
        64'hf0effe25_05130000,
        64'h551785ce_01367a63,
        64'h963e09da_47839e3d,
        64'h0087979b_0106161b,
        64'h09ea4783_09fa4603,
        64'hee0519e3_842af94f,
        64'hf0ef854a_85d2fe0a,
        64'h7a1302f1_0a13f006,
        64'h00e3ff25_05130000,
        64'h55178a09_000b8963,
        64'hfbc596e3_87ae0511,
        64'h08210133_09bb0ffb,
        64'hfb9300db_ebb300be,
        64'h96bbcb89_8b850107,
        64'hc78397a6_078e0208,
        64'h80630065_202302e8,
        64'hd33bb7f1_4b814a81,
        64'h4c81b7c1_ee4ff0ef,
        64'h01050513_00005517,
        64'h00030d63_02e8f33b,
        64'h0017859b_00082883,
        64'h4e114e85_478189d6,
        64'h856200c4_88138c0a,
        64'h009c9c9b_e3994b85,
        64'h02eadabb_02c92783,
        64'hbf415429_f24ff0ef,
        64'h01850513_00005517,
        64'hcb8902ec_f7bb0005,
        64'hac83e791_02eaf7bb,
        64'h060a8163_0045aa83,
        64'hdb450125_05130000,
        64'h55170989_27038082,
        64'h2a010113_23813d83,
        64'h24013d03_24813c83,
        64'h25013c03_25813b83,
        64'h26013b03_26813a83,
        64'h27013a03_27813983,
        64'h28013903_28813483,
        64'h29013403_29813083,
        64'h8522f840_0413f96f,
        64'hf0ef03a5_05130000,
        64'h5517e7b9_00167793,
        64'h07e94603_00e7eb63,
        64'h01850513_00005517,
        64'h84ae8b32_892abfe7,
        64'h87933ffc_07b79f3d,
        64'hbff7879b_bffc07b7,
        64'h4d180ac7_e9634789,
        64'h23b13c23_25a13023,
        64'h25913423_25813823,
        64'h25713c23_27613023,
        64'h27513423_27413823,
        64'h27313c23_29213023,
        64'h28913423_28813823,
        64'h28113c23_d6010113,
        64'h80826145_69a26942,
        64'h64e27402_70a28522,
        64'h013505a3_15e010ef,
        64'h8526842a_875ff0ef,
        64'h852685ca_00091c63,
        64'h00f51e63_842a57b5,
        64'hc519cc7f_f0ef84aa,
        64'h45850b30_06138edd,
        64'h892e9be1_0079f693,
        64'h0ff5f993_08154783,
        64'hf022f406_e44ee84a,
        64'hec267179_b74d84aa,
        64'hb75ddf40_0493f7d5,
        64'h0b944783_e51998df,
        64'hf0ef854a_85a29801,
        64'h01f10413_f1e92581,
        64'h99f5ffe4_059bf571,
        64'h84aad1ff_f0ef892a,
        64'h45850b90_0613842e,
        64'h4685fef7_60e34705,
        64'hffc5879b_80822401,
        64'h01132281_34832201,
        64'h39038526_23013403,
        64'h23813083_54a9c585,
        64'h468102b7_e16302f5,
        64'h88634789_23213023,
        64'h22913423_22813823,
        64'h22113c23_dc010113,
        64'hbf455929_bf555951,
        64'hbf651a04_b0235c80,
        64'h20efd169_1a04b503,
        64'h892abf4d_08f4aa23,
        64'h02f707bb_27852705,
        64'h8bfd8b7d_0057d79b,
        64'h00a7d71b_50fc8082,
        64'h25010113_22813983,
        64'h23013903_23813483,
        64'h854a2401_34032481,
        64'h308308f4_80230a74,
        64'h478308d4_ac2302f6,
        64'h86bb00a6_969b0dd4,
        64'h4783f8dc_07a60d44,
        64'h27830009_8663c799,
        64'h54dc08f4_aa2300a6,
        64'h979bc7b9_8b850e04,
        64'h46830af4_47830af4,
        64'h07a34785_ed35e0bf,
        64'hf0ef8526_45850af0,
        64'h06134685_ce81e391,
        64'h8bfd09c4_4783c789,
        64'h8b850a04_4783f4fc,
        64'h07a6c319_f4fc54d8,
        64'h9fb90884_47039fb9,
        64'h0087171b_08944703,
        64'h9fb90107_171b0187,
        64'h979b08a4_470308b4,
        64'h4783f8fc_07ce02e7,
        64'h87b30dd4_478302f7,
        64'h07330e04_470397ba,
        64'h08c44703_9fb90087,
        64'h171b0107_979b4685,
        64'h08d44703_08e44783,
        64'h04098f63_fca714e3,
        64'h0621070d_e21c07ce,
        64'h02b787b3_0dd44783,
        64'h02f585b3_0e044583,
        64'h00098c63_4685c391,
        64'h97aeffe7_45839fad,
        64'h0105959b_0087979b,
        64'h00074583_fff74783,
        64'he0fc07c6_468109d4,
        64'h05130a84_4783fcdc,
        64'h07c60c84_86130914,
        64'h07130e24_478306f4,
        64'h8fa309c4_4783c789,
        64'h8b890a04_47830009,
        64'h8a6308f4_80a30b34,
        64'h4783c789_0e244783,
        64'he7810019_f9938b85,
        64'h06f48f23_09b44983,
        64'h0a044783_f8dc00d7,
        64'h73630147_d69307a6,
        64'h80070713_67050d44,
        64'h278300e7_fd63cc98,
        64'h1ff78793_400407b7,
        64'h53b897ba_078affe7,
        64'h07130000_47171cf7,
        64'h6b634721_0c044783,
        64'h123010ef_85a22000,
        64'h06131e05_03631a04,
        64'hb5031aa4_b0237660,
        64'h20ef2000_0513e799,
        64'h1a04b783_1e051863,
        64'h892ac09f_f0ef84aa,
        64'h85a29801_01f10413,
        64'h1ce7f563_49013ffc,
        64'h07372331_34232291,
        64'h3c232481_30232411,
        64'h34239fb9_23213823,
        64'hbffc07b7_db010113,
        64'h4d18bfcd_fc79347d,
        64'h80826121_74a27442,
        64'h70e2d91f_f0ef8526,
        64'h3e800593_e919c53f,
        64'hf0ef8526_858a4601,
        64'h440dc436_84aafc06,
        64'hf426f822_8ed10106,
        64'h161b8edd_030007b7,
        64'h0086969b_c23e47f5,
        64'h00f11023_47997139,
        64'h80826121_6aa26a42,
        64'h69e274a2_79028526,
        64'h744270e2_fc0999e3,
        64'h9aa20287_84339a22,
        64'h408989b3_08c96783,
        64'hfc851ae3_f01ff0ef,
        64'h854a85d6_865286a2,
        64'h844e0089_f3630207,
        64'he4030109_378389a6,
        64'hf96decdf_f0ef854a,
        64'h08c92583_a0894481,
        64'hbd9ff0ef_41450513,
        64'h00005517_00b67a63,
        64'h014485b3_68100005,
        64'h4d638d3f_a0ef8522,
        64'h00b44583_c11d892a,
        64'h482010ef_8ab684b2,
        64'h8a2e4148_842ace05,
        64'he456e852_ec4ef04a,
        64'hf426f822_fc067139,
        64'hb7c54401_b7d50004,
        64'h841bb74d_02f6063b,
        64'hbf6147c5_80826125,
        64'h690664a6_644660e6,
        64'h8522c43f_f0ef45e5,
        64'h05130000_5517c11d,
        64'hd55ff0ef_d23ed402,
        64'h854a100c_47f54601,
        64'h02f11023_47b10497,
        64'hf0634785_e529842a,
        64'hd75ff0ef_c83eca26,
        64'hd23a854a_100c4785,
        64'h0030cc3e_e42e4755,
        64'hd432cf31_08c92783,
        64'h260102f1_102302c9,
        64'h270347c9_06d7f663,
        64'h84b6892a_4785e8a2,
        64'hec86e0ca_e4a6711d,
        64'h80824501_bfd54501,
        64'h80826121_74a27442,
        64'h70e2f8ed_34fdc901,
        64'hdcdff0ef_8522858a,
        64'h46014495_cb918b89,
        64'h1b842783_c11dde3f,
        64'hf0efc23e_842af426,
        64'hfc06f822_858a4601,
        64'h47d5c42e_00f11023,
        64'h47c17139_e7a919c5,
        64'h2783bf7d_f9200513,
        64'hd09ff0ef_50450513,
        64'h00005517_fc8049e3,
        64'h4501b755_5d8020ef,
        64'h3e800513_00f05763,
        64'h0014079b_347dfe04,
        64'hc6e334fd_80826125,
        64'h7aa27a42_79e26906,
        64'h64a66446_60e6fba0,
        64'h0513d4bf_f0ef52e5,
        64'h05130000_5517c78d,
        64'h0125f7b3_05479363,
        64'h0135f7b3_c7891005,
        64'hf79345b2_ed0de73f,
        64'hf0ef8556_858a4601,
        64'he00a0a13_e0098993,
        64'h08090913_4495c43e,
        64'h842e8aaa_ec86f456,
        64'he4a6e8a2_6a056989,
        64'hfdf94937_0107979b,
        64'hf852fc4e_e0ca07c5,
        64'h5783c23e_47d500f1,
        64'h102347b5_711d8082,
        64'h61457402_70a2c43c,
        64'h47b2e119_ec9ff0ef,
        64'h8522858a_4601c43e,
        64'h8fd98f55_400006b7,
        64'h8f756000_06b78ff5,
        64'h8ff9f807_87934ad4,
        64'h008007b7_45386914,
        64'hc195842a_c402c23e,
        64'hf406f022_478500f1,
        64'h10234785_71798082,
        64'h61457402_70a28522,
        64'h6cc020ef_7d000513,
        64'he509842a_f21ff0ef,
        64'hc202c402_00011023,
        64'h858a4601_85226ea0,
        64'h20eff406_3e800513,
        64'h842af022_7179b761,
        64'hfb600513_d55156f0,
        64'h10ef0d44_85130d44,
        64'h05934611_00f71a63,
        64'h0e044783_0e04c703,
        64'h02f71063_0c044783,
        64'h0c04c703_02f71663,
        64'h0dd44783_0dd4c703,
        64'h02f71c63_0a044783,
        64'h0a04c703_f579f95f,
        64'hf0ef1a05_34832211,
        64'h3c232291_342385a2,
        64'h980101f1_04132281,
        64'h3823dc01_01138082,
        64'h24010113_22813483,
        64'h23013403_23813083,
        64'h45018082_450100e6,
        64'hfe634004_07374d14,
        64'h80826161_60a6fd3f,
        64'hf0efcc3e_d402e486,
        64'h100c2000_07930030,
        64'he83ee42e_07851782,
        64'h4785d23e_47d502f1,
        64'h102347a1_715d8302,
        64'h0007b303_679c691c,
        64'h80826d25_05130000,
        64'h55178082_6108953e,
        64'h81754527_87930000,
        64'h47971502_00a7eb63,
        64'h47ad8082_557d8082,
        64'h01416402_60a24501,
        64'h83020141_60a26402,
        64'h85220003_07630207,
        64'hb303679c_681c0005,
        64'h5e63ff5f_f0ef842a,
        64'he406e022_11418082,
        64'h557d8082_557db7e9,
        64'h659c95aa_058e05e1,
        64'h35f1bfd9_617cbfe9,
        64'h7d5c8082_61054501,
        64'he91c64a2_644260e2,
        64'h02f457b3_93810204,
        64'h97930c50_10ef7540,
        64'hf55c08c5_2483795c,
        64'h878297ba_e426e822,
        64'hec061101_439c97ba,
        64'h83f94ca7_07130000,
        64'h47170205_979304b7,
        64'hee63479d_80824501,
        64'h83020003_03630087,
        64'hb303679c_691c8082,
        64'h61356452_60f28522,
        64'h129020ef_0808842a,
        64'he3fff0ef_e436eec6,
        64'heac2e6be_e2baea22,
        64'hee060808_10000593,
        64'h1234862a_fe36fa32,
        64'hf62e710d_80826161,
        64'h60e2e69f_f0efe436,
        64'he4c6e0c2_fc3ef83a,
        64'hec061000_05931014,
        64'h862ef436_f032715d,
        64'h80826161_60e2e8df,
        64'hf0efe436_e4c6e0c2,
        64'hfc3ef83a_ec061034,
        64'hf436715d_b7f18522,
        64'h02010393_0005059b,
        64'h4db010ef_85220124,
        64'h74336000_00840b13,
        64'hb5fd845a_d93ff0ef,
        64'h00840b13_02010393,
        64'h00044503_a809ddbf,
        64'hf0ef0028_02010393,
        64'h0005059b_e37ff0ef,
        64'h400845a9_46010016,
        64'hb6930038_00840b13,
        64'hf8b50693_a81145c1,
        64'h00163613_46850038,
        64'h00840b13_fa850613,
        64'hf6e510e3_07800713,
        64'h02e50063_07500713,
        64'ha00d4601_46850038,
        64'h00840b13_f6e51ee3,
        64'h07000713_00a76c63,
        64'h06e50e63_07300713,
        64'hb74d048d_0024c503,
        64'h80826109_0007051b,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_744670e6,
        64'hf55d08f5_09630630,
        64'h079304d5_0f630580,
        64'h069302a6_eb6306d5,
        64'h0f630640_06930489,
        64'h0014c503_478100f6,
        64'hf36346a5_0ff7f793,
        64'hfd07879b_cb9d0004,
        64'hc7830355_10634781,
        64'h04890545_0f630014,
        64'hc503bfe1_e7bff0ef,
        64'h02010393_04850135,
        64'h086304d7_ff639381,
        64'h17827682_0017079b,
        64'hc52d8f1d_0004c503,
        64'h77a27742_02095913,
        64'h03000a93_06c00a13,
        64'h02500993_f82af02e,
        64'hf42afc3e_843684b2,
        64'he0dafc86_e4d6e8d2,
        64'heccef4a6_f8a2597d,
        64'h011cf0ca_7119b7f1,
        64'h06850117_80230066,
        64'h80232605_0006c883,
        64'h0007c303_97ba9381,
        64'h178240c8_07bbb7d9,
        64'h2585fea6_8fa30685,
        64'hbf5d00a8_053b8082,
        64'h00b61b63_fff5081b,
        64'h86ba2581_00068023,
        64'h0015559b_40e6853b,
        64'h068500f6_802302d0,
        64'h07930008_876302f5,
        64'he9630300_051340e6,
        64'h85bbfe71_8532fea6,
        64'h8fa30685_0ff57513,
        64'h02b6563b_0305051b,
        64'h046e6763_0ff37513,
        64'h02b6733b_0005061b,
        64'h385986ba_4e250ff6,
        64'hf8130410_0693c219,
        64'h06100693_488540a0,
        64'h053be681_00055663,
        64'h4881bfe9_00d70023,
        64'h07850007_c68300d3,
        64'hb8230017_06938082,
        64'h852e0007_002300b6,
        64'he6630103_b70340a7,
        64'h86bb87aa_9d9dfff7,
        64'h059b00c6_f5638e9d,
        64'hfff70693_0003b703,
        64'h8f999201_02059613,
        64'h0103b783_0083b703,
        64'h80824501_80820007,
        64'h80234505_0103b783,
        64'h00a70023_00f3b823,
        64'h00170793_00d7fe63,
        64'h93811782_278540f7,
        64'h07b30003_b6830083,
        64'hb7830103_b7038082,
        64'h61454501_6a0269a2,
        64'h694264e2_740270a2,
        64'h2e8000ef_08450513,
        64'h00006517_fd249fe3,
        64'h04052fa0_00ef8191,
        64'h00f5f613_2485854e,
        64'h00044583_30c000ef,
        64'h855285a6_e78901f4,
        64'hf7932000_0913ad69,
        64'h89930000_6997ad6a,
        64'h0a130000_6a174481,
        64'hed5ff0ef_84264581,
        64'h852633a0_00efad65,
        64'h05130000_6517dae6,
        64'h06130000_6617e789,
        64'ha5060613_00006617,
        64'h584c19c4_2783dc3f,
        64'hb0ef0fa5_85930000,
        64'h65977448_102030ef,
        64'haf850513_00006517,
        64'h378000ef_aec50513,
        64'h00006517_a7458593,
        64'h00006597_c789a865,
        64'h85930000_6597545c,
        64'h398000ef_afc50513,
        64'h00006517_5c0c3a60,
        64'h00ef2601_0ff6f693,
        64'h0ff7f793_0ff77713,
        64'h0187d61b_0107d69b,
        64'h0087d71b_b0c50513,
        64'h00006517_06c44583,
        64'h583c3d20_00ef91c1,
        64'h15c20085_d59bb165,
        64'h05130000_6517546c,
        64'h3e8000ef_b0c50513,
        64'h00006517_06f44583,
        64'h3f8000ef_638cb0e5,
        64'h05130000_6517681c,
        64'h206010ef_842a4910,
        64'h10ef4501_44b010ef,
        64'h0001b503_1b2030ef,
        64'hb2850513_00006517,
        64'h84aa0aa0_30efe052,
        64'he44ee84a_ec26f022,
        64'hf4062000_05137179,
        64'h7940006f_61054685,
        64'h60e26622_644285a2,
        64'h4d3010ef_e42eec06,
        64'h4501842a_e8221101,
        64'h80820141_640260a2,
        64'h557de391_4505703c,
        64'h170030ef_ac450513,
        64'h00006517_ab458593,
        64'h00006597_34c00613,
        64'h97068693_00005697,
        64'h02f40263_200007b7,
        64'he4066380_e0221141,
        64'h711c8082_25016108,
        64'h953e050e_200007b7,
        64'hf73ff06f_20000537,
        64'h45814609_8082bff9,
        64'h557d18c0_30ef8522,
        64'hb7e5c45c_4785d4fd,
        64'h45018885_80826145,
        64'h69a26942_64e27402,
        64'h70a24501_c45c4789,
        64'hcb990024_f793f404,
        64'h01242423_e01c2000,
        64'h07b70209_8b634fe0,
        64'h00efbd25_05130000,
        64'h65178622_85aa89aa,
        64'h785010ef_9d450513,
        64'h00005517_85a2cc1d,
        64'h5551842a_1a4030ef,
        64'h892e84b2_e44ef406,
        64'he84aec26_f0220480,
        64'h05137179_08b04163,
        64'h5535b7dd_87ca0ca1,
        64'h39a020ef_e43e002c,
        64'h46218566_639c0087,
        64'h8913fa97_8de394be,
        64'h00093c83_01096483,
        64'h97a667a1_bf41b1df,
        64'hf0ef8522_b77100f9,
        64'h2623000c_b783dbd9,
        64'h8b85bd95_641020ef,
        64'h4505d80c_8ee3c47f,
        64'hf0ef8522_484cc85c,
        64'h9bf54c85_485cb4df,
        64'hf0ef8522_ef8d8b85,
        64'h00892783_00090963,
        64'h04043023_2b4030ef,
        64'h855685d2_0ca00613,
        64'ha6868693_00005697,
        64'h01748c63_04043903,
        64'h6004cc9d_4c858889,
        64'hc85c9bf9_485cc85c,
        64'h0027e793_485ccbb5,
        64'h603cfeb6_90e30791,
        64'h872a2685_c3988f51,
        64'h8361ff87_37030106,
        64'h8763c390_0086161b,
        64'hff870513_63104591,
        64'h480d4681_00c90793,
        64'h018c8713_08e69f63,
        64'h0037f693_470d0204,
        64'h3c230049_2783cba9,
        64'h7c1c3320_30ef8556,
        64'h85d209c0_0613ace6,
        64'h86930000_5697017c,
        64'h8c630384_39030004,
        64'h3c83cfb5_0014f793,
        64'h658000ef_d0450513,
        64'h00006517_85cad1ff,
        64'hf0ef85ca_00496913,
        64'hff397913_85220144,
        64'h2903c395_0084f793,
        64'h680000ef_d0450513,
        64'h00006517_85cad47f,
        64'hf0ef85ca_00896913,
        64'hff397913_85220144,
        64'h2903c395_0044f793,
        64'hb27ff0ef_85224581,
        64'hb6fff0ef_85224581,
        64'hcc5cf920_0793c781,
        64'h7c1c00f7_6f630c89,
        64'h37830209_37031204,
        64'h8e632481_8cfd4c81,
        64'h485c0709_34833de0,
        64'h30ef8556_85d20f20,
        64'h061386e2_01790963,
        64'h00043903_b7116f60,
        64'h00efd625_05130000,
        64'h6517b625_85930000,
        64'h5597000b_1d633b7d,
        64'h20000bb7_8b4ebd61,
        64'h00c4e493_bd8541e0,
        64'h30efd725_05130000,
        64'h6517d625_85930000,
        64'h65971490_0613b7e6,
        64'h86930000_5697b765,
        64'h47014781_2585e31c,
        64'h97469381_83751782,
        64'h170200be_873b8fd9,
        64'h8fe90107_67330087,
        64'hd79b01c8_78330087,
        64'h981b0107_67330187,
        64'h971b0187_d81bf2e5,
        64'h00670363_16fd0605,
        64'h27810107_e7b301e8,
        64'h183b0705_00371f1b,
        64'h00064803_ec0689e3,
        64'h6e89f005_051300ff,
        64'h0e374311_47014781,
        64'h45816390_0107e683,
        64'h65410004_3883603c,
        64'hee079be3_8b85449c,
        64'hdf3ff0ef_8522488c,
        64'hdb7ff0ef_e0248522,
        64'h44cc8082_61654501,
        64'h6ce27c02_7ba27b42,
        64'h7ae26a06_69a66946,
        64'h64e67406_70a6efe9,
        64'h485ce42a_8a930000,
        64'h6a976819_8993eb7f,
        64'hf0ef2581_0015e593,
        64'h009899b7_85220d89,
        64'hb583cd1f_f0ef8522,
        64'h4585e93f_f0ef8522,
        64'h24058593_000f45b7,
        64'hd27ff0ef_85224581,
        64'h46054685_4705cf5f,
        64'hf0ef8522_4581cbdf,
        64'hf0ef8522_85a6c81f,
        64'hf0efe82a_0a130000,
        64'h6a178522_00095583,
        64'hc4fff0ef_cdcc0c13,
        64'h00005c17_85220089,
        64'h2583be1f_f0ef8522,
        64'h4581d71f_f0ef8522,
        64'h45814605_46814705,
        64'h0144e493_16078663,
        64'h8b85008a_2783000a,
        64'h09638cdd_03243c23,
        64'h4c1c4485_e391448d,
        64'h8b89c709_0017f713,
        64'h44810049_278316f9,
        64'h9a630404_3a032000,
        64'h07b70004_3983bf5f,
        64'hf0ef4585_60080e04,
        64'h9c636ca0_20ef00c9,
        64'h05134581_4611d01c,
        64'he03084b2_892e0005,
        64'hd7830204_08a3ec66,
        64'hf062f45e_f85afc56,
        64'he0d2e4ce_f486e8ca,
        64'heca67100_f0a27159,
        64'h80826105_690264a2,
        64'h644260e2_c8440499,
        64'h3c236120_30eff665,
        64'h05130000_6517f565,
        64'h85930000_65970760,
        64'h0613d626_86930000,
        64'h569702f9_026384ae,
        64'h842a2000_07b7ec06,
        64'he426e822_00053903,
        64'he04a1101_80826105,
        64'h64a26442_60e2e424,
        64'h658030ef_fac50513,
        64'h00006517_f9c58593,
        64'h00006597_06f00613,
        64'hd9868693_00005697,
        64'h02f40263_84ae2000,
        64'h07b7ec06_e4266100,
        64'he8221101_80826105,
        64'h64a26442_60e2e0a0,
        64'h8c7d17fd_678569e0,
        64'h30efff25_05130000,
        64'h6517fe25_85930000,
        64'h65970680_0613dce6,
        64'h86930000_569702f4,
        64'h8263842e_200007b7,
        64'hec06e822_6104e426,
        64'h11018082_610564a2,
        64'h644260e2_fc809041,
        64'h14426e20_30ef0365,
        64'h05130000_65170265,
        64'h85930000_65970610,
        64'h0613e026_86930000,
        64'h569702f4_8263842e,
        64'h200007b7_ec06e822,
        64'h6104e426_1101d4df,
        64'hf06f0141_458160a2,
        64'h64026008_f23ff0ef,
        64'h46054685_47054581,
        64'h8522ef1f_f0ef4581,
        64'h8522f39f_f0ef842a,
        64'h45810405_30230205,
        64'h3c234605_46814705,
        64'he022e406_11418082,
        64'h01414501_640260a2,
        64'hd97ff0ef_45816008,
        64'hf67ff0ef_45814605,
        64'h46854705_8522f35f,
        64'hf0ef4581_8522f7df,
        64'hf0efe406_45818522,
        64'h46054681_47057100,
        64'he0221141_80826121,
        64'h69e27902_74a202b9,
        64'hb8238dc5_744270e2,
        64'h88a10125_e5b30034,
        64'h949b8dd9_00497913,
        64'h0029191b_8b058989,
        64'h0014159b_67227c60,
        64'h30efe43a_11c50513,
        64'h00006517_10c58593,
        64'h00006597_05a00613,
        64'hed868693_00005697,
        64'h02f98463_84368932,
        64'h84ae2000_07b7fc06,
        64'hf04af426_f8220005,
        64'h3983ec4e_71398082,
        64'h610564a2_644260e2,
        64'hf4040130_30ef1665,
        64'h05130000_65171565,
        64'h85930000_65970530,
        64'h0613f126_86930000,
        64'h569702f4_026384ae,
        64'h200007b7_ec06e426,
        64'h6100e822_11018082,
        64'h610564a2_644260e2,
        64'hf0040530_30ef1a65,
        64'h05130000_65171965,
        64'h85930000_659704c0,
        64'h0613f426_86930000,
        64'h569702f4_026384ae,
        64'h200007b7_ec06e426,
        64'h6100e822_11018082,
        64'h610564a2_644260e2,
        64'hec809001_14020970,
        64'h30ef1ea5_05130000,
        64'h65171da5_85930000,
        64'h65970450_0613e566,
        64'h86930000_769702f4,
        64'h8263842e_200007b7,
        64'hec06e822_6104e426,
        64'h11018082_610564a2,
        64'h644260e2_e8809001,
        64'h14020db0_30ef22e5,
        64'h05130000_651721e5,
        64'h85930000_659703e0,
        64'h0613ea26_86930000,
        64'h769702f4_8263842e,
        64'h200007b7_ec06e822,
        64'h6104e426_11018082,
        64'h610564a2_644260e2,
        64'he40411b0_30ef26e5,
        64'h05130000_651725e5,
        64'h85930000_65970360,
        64'h0613ffa6_86930000,
        64'h569702f4_026384ae,
        64'h200007b7_ec06e426,
        64'h6100e822_11018082,
        64'h610564a2_644260e2,
        64'he00415b0_30ef2ae5,
        64'h05130000_651729e5,
        64'h85930000_659702f0,
        64'h061302a6_86930000,
        64'h569702f4_026384ae,
        64'h200007b7_ec06e426,
        64'h6100e822_11018082,
        64'h610564a2_644260e2,
        64'hfc2419b0_30ef2ee5,
        64'h05130000_65172de5,
        64'h85930000_65970880,
        64'h06130526_86930000,
        64'h569702f5_026384ae,
        64'h842a2000_07b7ec06,
        64'he426e822_11018082,
        64'h556dbfe5_0007ac23,
        64'h80824501_cf980200,
        64'h071300d7_17634691,
        64'h00d70d63_711c46a1,
        64'h59588082_6149640a,
        64'h60aaf83f_f0ef0808,
        64'hf01ff0ef_0808e85f,
        64'hf0ef0808_85a26622,
        64'hf71ff0ef_e42ee506,
        64'h0808842a_e1227175,
        64'h80826105_12450513,
        64'h00007517_60e2fca7,
        64'h1de3fef6_8fa3fec6,
        64'h8f230007_c78397ae,
        64'h00064603_8bbd962e,
        64'h0047d613_07050689,
        64'h0007c783_00e107b3,
        64'h454137a5_85930000,
        64'h65971626_86930000,
        64'h76974701_3bf020ef,
        64'hec06850a_46410505,
        64'h05931101_8082e13c,
        64'hb6c78793_00000797,
        64'hed3c639c_f4478793,
        64'h00007797_e93c0405,
        64'h3423639c_f4c78793,
        64'h00007797_80826145,
        64'h69a26942_64e27402,
        64'h70a2fd24_fde34501,
        64'h97828522_603cfc1c,
        64'h078e643c_0124f563,
        64'h3c9020ef_95224581,
        64'h92011602_0006091b,
        64'h40a9863b_449d0400,
        64'h099300e7_802397a2,
        64'hf8000713_00178513,
        64'he84af406_e44eec26,
        64'h842a03f7_f793f022,
        64'h7179653c_80826161,
        64'h6ba26b42_6ae27a02,
        64'h79a27942_74e26406,
        64'h60a6b7c9_97824401,
        64'h852660bc_01741763,
        64'h99d64159_09334810,
        64'h20ef0144_043b8656,
        64'h00848533_85ce020a,
        64'hda93020a_1a930009,
        64'h0a1b00f9_74639381,
        64'h17820007_8a1b408b,
        64'h07bb0400_0b930400,
        64'h0b13e53c_893289ae,
        64'h84aa97b2_03f7f413,
        64'hec56f052_e486e45e,
        64'he85af44e_f84afc26,
        64'he0a2715d_653c8082,
        64'h61056922_64c2cd70,
        64'hcd34c97c_05052823,
        64'h00c8863b_00d306bb,
        64'h00fe07bb_010e883b,
        64'h6462f3ef_9de300e5,
        64'h87bb0005_869b0003,
        64'h861b0f11_8f5d0157,
        64'h171b00b7_579b9f3d,
        64'h00774733_9fa18f4d,
        64'hfff74713_0007081b,
        64'h00b385bb_40809fa1,
        64'h8dd50115_d59b94aa,
        64'h00f5969b_048a9db5,
        64'hffc2a403_8db902c1,
        64'h0075e5b3_fff7c593,
        64'h023f4483_9ead00c7,
        64'h03bb00c3_e633400c,
        64'h9ead0166_561b00a6,
        64'h139b0082_a5839e2d,
        64'h8e3d8e59_fff6c613,
        64'h9db100f8_073b0107,
        64'h683301a8_581b0003,
        64'ha5839e2d_0068171b,
        64'h0107083b_0042a583,
        64'h9f2d942a_040a418c,
        64'h95aa058a_93aa038a,
        64'h020f4583_9f2d022f,
        64'h4403021f_43830002,
        64'ha70300d7_45b38f5d,
        64'hfff64713_2a428293,
        64'h00005297_f5f592e3,
        64'h00e407bb_0004069b,
        64'h0002861b_0f918f5d,
        64'h0177171b_0097579b,
        64'h9f3d8f21_9fa50057,
        64'h47330007_081b00d2,
        64'h843b8ec1_00092483,
        64'h0106d69b_9fa50106,
        64'h941b992a_9ea1090a,
        64'h0056c6b3_00e7c6b3,
        64'hffc3a483_9c3500c7,
        64'h02bb03c1_00c2e633,
        64'h0156561b_013fc903,
        64'h00b6129b_408000c2,
        64'h863b9ea1_94aa00e2,
        64'hc2b3048a_00f8073b,
        64'h0083a403_9e210107,
        64'h683301c8_581b0048,
        64'h171b012f_c4830107,
        64'h083b4080_9e2194aa,
        64'h048a0043_a4039f21,
        64'h011fc483_9f254000,
        64'h00c2c4b3_942a040a,
        64'h00d7c2b3_0003a703,
        64'h010fc403_32c38393,
        64'h00005397_8ffa3b6f,
        64'h0f130000_5f17f255,
        64'h99e300e4_07bb0004,
        64'h069b0003_861b000f,
        64'h081b8f5d_0147171b,
        64'h00c7579b_9f3d0077,
        64'h473301e7_77330083,
        64'hc7339fb9_00d3843b,
        64'h8ec14098_0126d69b,
        64'h9fb900e6_941b94aa,
        64'h048affcf_a7039eb9,
        64'h0fc101e6_c6b3fff5,
        64'hc4838efd_007f46b3,
        64'h05919f35_00cf03bb,
        64'h00c3e633_40189eb9,
        64'h0176561b_0096139b,
        64'h008fa703_9e398e3d,
        64'h8e7501e7_c6339f31,
        64'h00f80f3b_010f6833,
        64'h0003a703_01b8581b,
        64'h9e390058_1f1b010f,
        64'h083b004f_a70300ef,
        64'h0f3b942a_040a4318,
        64'h972a070a_93aa038a,
        64'h0005c703_00ef0f3b,
        64'h0025c403_0015c383,
        64'h000faf03_01e6c733,
        64'h00cf7f33_00d7cf33,
        64'h4a028293_00005297,
        64'h3d8f8f93_00005f97,
        64'h4a058593_00005597,
        64'hf45f17e3_00e387bb,
        64'h0003869b_0005881b,
        64'h0f418f5d_0167171b,
        64'h00a7579b_9f3d8f2d,
        64'h9fa10077_77338f2d,
        64'h0007061b_00d703bb,
        64'hffcfa403_9fa100d3,
        64'he6b30116_969b00f6,
        64'hd39b0076_86bb8ebd,
        64'h00cf2403_8ef900b7,
        64'hc6b300d3_83bb00c5,
        64'h873b0083_83bb8e59,
        64'h0146561b_00c6171b,
        64'h9e39008f_23838e35,
        64'h8e6d00f6_c6339f31,
        64'h00f805bb_0077073b,
        64'h0105e833_0198581b,
        64'h0078159b_0105883b,
        64'h004f2703_ff4fa383,
        64'h9db90075_85bb0fc1,
        64'h008fa403_000f2583,
        64'h000fa383_00b64733,
        64'h8dfd00c6_c5b345ef,
        64'h8f930000_5f978876,
        64'h87f2869a_86460405,
        64'h02938f2a_e44ae826,
        64'hec221101_05c52883,
        64'h05852303_05452e03,
        64'h05052e83_bf89eaf7,
        64'h1de30e50_07930181,
        64'h4703f8d7_71e30007,
        64'h869b0200_06134729,
        64'h93811782_f4c7e5e3,
        64'h05850685_00e58023,
        64'hf91780e3_b751842a,
        64'hbf1900e7_85a34721,
        64'h6786ae5f_d0ef082c,
        64'h462d6506_b07fd0ef,
        64'h45810200_06136506,
        64'hf4450005_041ba55f,
        64'he0ef1028_dbd50181,
        64'h478302f5_1b634791,
        64'hb7c10005_041b8fef,
        64'he0ef00f5_02234785,
        64'h752200f5_00235795,
        64'ha8850785_00c68023,
        64'h00fe06b3_b7cdffe8,
        64'h1be30608_05630005,
        64'h48030505_bfcdf36d,
        64'h80826125_644660e6,
        64'h85224419_00eef863,
        64'ha8210007_0f1b8e65,
        64'h05130000_75179341,
        64'h17423701_00a36c63,
        64'h91411542_f9f7051b,
        64'h27850006_c70348b1,
        64'h07f00e93_43658e2e,
        64'h4781082c_feb706e3,
        64'h00074703_97369301,
        64'h02079713_fff6079b,
        64'hbf45863e_b74d2605,
        64'ha06100e7_8ca30007,
        64'h8ba30007_8b230460,
        64'h071300e7_8c230210,
        64'h07136786_bc7fd0ef,
        64'h082c462d_c3dd6506,
        64'h01814783_e1792501,
        64'habbfe0ef_10284585,
        64'he8410005_041bbd6f,
        64'he0efda02_10284581,
        64'hea290200_0593eba1,
        64'h0007c783_97b69381,
        64'h02061793_46010001,
        64'h0c2366a2_ec550005,
        64'h041bee3f_d0efec86,
        64'he8a21028_002c4605,
        64'he42a711d_b7d5842a,
        64'hbf550004_802300f5,
        64'h15634791_80826125,
        64'h690664a6_644660e6,
        64'h852200a9_2023c29f,
        64'hd0ef953e_03478793,
        64'h02700793_00e68463,
        64'h00054683_04300793,
        64'h470d6562_e0150005,
        64'h041be69f_d0ef510c,
        64'h65620209_0a63fec7,
        64'h83e3177d_0007c783,
        64'h97a69381_17820007,
        64'h869bfff6_879bce89,
        64'h00070023_02000613,
        64'h46ad00b4_8713ca1f,
        64'hd0ef8526_462d75c2,
        64'he93d2501_b8ffe0ef,
        64'h08284585_e5592501,
        64'hca8fe0ef_d2020828,
        64'h4581c4b9_e0510005,
        64'h041bf9bf_d0efec86,
        64'he8a20828_4601002c,
        64'h893284ae_e42ae0ca,
        64'he4a6711d_80826125,
        64'h644660e6_2501ad6f,
        64'he0ef00f5_02234785,
        64'h00e78ca3_0087571b,
        64'h00e78c23_00445703,
        64'h00e78ba3_0087571b,
        64'h00e78b23_75220064,
        64'h5703cb85_6786eb95,
        64'h0207f793_00b7c783,
        64'h451967a6_e1292501,
        64'h9abfe0ef_e4be1028,
        64'h083c65a2_e9292501,
        64'h810fe0ef_ec861028,
        64'h002c4605_842ee42a,
        64'he8a2711d_bfcd47a1,
        64'h8082614d_853e64ea,
        64'h740a70aa_0005079b,
        64'hb50fe0ef_6506e791,
        64'h0005079b_e24fe0ef,
        64'h008800f7_022306d7,
        64'h07a34785_06f704a3,
        64'h0086d69b_0106d69b,
        64'h0087d79b_0107d79b,
        64'h0107979b_06f70423,
        64'h27810107_d79b06f7,
        64'h07230107_969b57d6,
        64'h02f69d63_05574683,
        64'h02e00793_6706efb1,
        64'h0005079b_fc3fd0ef,
        64'h8522c5a5_47890005,
        64'h059bcaef_e0ef8522,
        64'h0005059b_f2dfd0ef,
        64'h85a60004_450306f7,
        64'h086357d6_4736cbbd,
        64'h8bc100b4_c78300f4,
        64'h02234785_00f485a3,
        64'h0207e793_64060281,
        64'h4783e0df_d0ef00d4,
        64'h851302a1_0593464d,
        64'h648aefc5_0005079b,
        64'hdc5fe0ef_10a80ce7,
        64'h93634711_cbf90005,
        64'h079baadf_e0ef10a8,
        64'h65820c05_4d6347ad,
        64'hf05fd0ef_850ae49f,
        64'hd0ef10a8_008c0280,
        64'h0613e55f_d0ef1028,
        64'h05ad4655_0e058e63,
        64'h479165e6_10071263,
        64'h02077713_479900b7,
        64'hc7037786_10079a63,
        64'h0005079b_af7fe0ef,
        64'hf0be083c_f4be0088,
        64'h65a26786_12079663,
        64'h0005079b_964fe0ef,
        64'hed26f122_f5060088,
        64'h002c4605_e02ee42a,
        64'h71718082_616564e6,
        64'h740670a6_2501c9ef,
        64'he0ef00f5_02234785,
        64'h008705a3_8c3d0274,
        64'h74138c65_8cbd7522,
        64'h00b74783_c30d6706,
        64'he39d0207_f79300b7,
        64'hc7834519_67a6e915,
        64'h2501b65f_e0efe4be,
        64'h1028083c_65a2e131,
        64'h25019caf_e0eff486,
        64'h10284605_002c8432,
        64'h84aee42a_eca6f0a2,
        64'h7159b7c5_44218082,
        64'h614d6d46_6ce67c06,
        64'h7ba67b46_7ae66a0a,
        64'h69aa694a_64ea740a,
        64'h70aa8522_f25fe0ef,
        64'h85ca7522_441db749,
        64'h8c6a0ffb_fb93f61f,
        64'hd0ef3bfd_85524581,
        64'h20000613_ec090005,
        64'h041b8dcf_e0ef0195,
        64'h02230385_2823001c,
        64'h0d1b7522_a82d0005,
        64'h041bd5af_e0ef00f5,
        64'h02234785_00978aa3,
        64'h01678a23_01378da3,
        64'h01578d23_00e78ca3,
        64'h00078ba3_00078b23,
        64'h04600713_00e78c23,
        64'h02100713_00e785a3,
        64'h75224741_6786e835,
        64'h0005041b_f59fe0ef,
        64'h1028040b_99634c85,
        64'h00274b83_06f404a3,
        64'h06d407a3_0087d79b,
        64'h0086d69b_0107d79b,
        64'h0106d69b_0107979b,
        64'h06f40423_27810107,
        64'hd79b0107_969b06f4,
        64'h07234781_00f69363,
        64'h571400d6_166357d2,
        64'h00074603_468d0574,
        64'h0aa37722_80efe0ef,
        64'h05440513_85d20494,
        64'h04a30564_04230534,
        64'h07a30554_07230404,
        64'h05a30404_05230374,
        64'h0a230200_061304f4,
        64'h06a30084_d49b0089,
        64'hd99b0460_07930ff9,
        64'h7a9304f4_062302e0,
        64'h0b930104_d49b0210,
        64'h07930109_d99b02f4,
        64'h0fa30104_949b0109,
        64'h199b0ff4_fb1347c1,
        64'h248188cf_e0ef8552,
        64'h02000593_462d898f,
        64'he0ef8552_00050c1b,
        64'h45812000_06130344,
        64'h0a13f6ef_e0ef8522,
        64'h0109549b_85ca7422,
        64'h16041463_0005041b,
        64'ha98fe0ef_752216f9,
        64'h0b634405_57fd16f9,
        64'h0f634409_47851809,
        64'h02630005_091bb45f,
        64'he0ef4581_75221807,
        64'h9f630207_f79300b7,
        64'hc7834419_67a61af4,
        64'h17634791_1c040963,
        64'h0005041b_d67fe0ef,
        64'he4be1028_083c65a2,
        64'h1c041463_0005041b,
        64'hbd0fe0ef_e8eaece6,
        64'hf0e2f4de_f8dafcd6,
        64'he152e54e_e94aed26,
        64'hf506f122_1028002c,
        64'h4605e42a_7171b769,
        64'hd5752501_91cff0ef,
        64'h85a27502_bf612501,
        64'hf20fe0ef_7502e411,
        64'hf1552501_9f5fe0ef,
        64'h1008faf5_18e34791,
        64'hd94d2501_836ff0ef,
        64'h00a84581_f1612501,
        64'h951fe0ef_caa200a8,
        64'h458996cf_e0ef00a8,
        64'h100c0280_0613fc87,
        64'h8de30149_2783c89d,
        64'h88c1cc0d_0005041b,
        64'had8fe0ef_00094503,
        64'h79028082_61497946,
        64'h74e6640a_60aa451d,
        64'hcb810014_f79300b5,
        64'hc483c599_75e2eb89,
        64'h0207f793_00b7c783,
        64'h45196786_e1052501,
        64'he3bfe0ef_e0be1008,
        64'h081c65a2_e9052501,
        64'hca0fe0ef_f8cafca6,
        64'he122e506_1008002c,
        64'h4605e42a_7175b7b1,
        64'h00f40523_fbf7f793,
        64'h00a44783_f55d2501,
        64'h6ec040ef_03040593,
        64'h0017c503_46854c50,
        64'h601cdba5_0407f793,
        64'h00a44783_fcf96ae3,
        64'h4d1c6008_fcf900e3,
        64'h45094785_b769449d,
        64'hb7e12501_a1cff0ef,
        64'h85ca6008_f9792501,
        64'hb37fe0ef_167d1000,
        64'h06374c0c_b7dd4505,
        64'h02f91463_57fd0005,
        64'h091b94df_e0ef4c0c,
        64'hbf7d84aa_00a405a3,
        64'hc5390004_2a232501,
        64'ha58ff0ef_484cef01,
        64'h600800f4_0523c818,
        64'h0207e793_fed772e3,
        64'h48144458_cf390027,
        64'hf71300a4_47838082,
        64'h610564a2_69028526,
        64'h644260e2_0007849b,
        64'hcb9100b4_4783e491,
        64'h0005049b_bc4fe0ef,
        64'h842ae04a_ec06e426,
        64'he8221101_bfad8a2a,
        64'hbfbd4a09_b7494a05,
        64'hb7c539f1_09112485,
        64'he1116582_01557533,
        64'h2501abcf_e0efe02e,
        64'h854ab745_fc0c94e3,
        64'h3cfd39f9_09092485,
        64'he3918fd9_0087979b,
        64'h00094703_00194783,
        64'h038b9163_20000993,
        64'h03440913_85cee921,
        64'h2501d10f_e0ef0015,
        64'h899b8522_00099e63,
        64'h1afd4c09_44814981,
        64'h49011000_0ab7504c,
        64'hb74d009b_202300f4,
        64'h02a30017_e793c804,
        64'h00544783_fef963e3,
        64'h29054c1c_2485e111,
        64'h09550863_09350863,
        64'h2501a55f_e0ef8522,
        64'h85ca4a85_59fd4481,
        64'h490902fb_9f634785,
        64'h00044b83_80826165,
        64'h6ce27c02_7ba27b42,
        64'h7ae26a06_69a66946,
        64'h64e68552_740670a6,
        64'h00fb2023_02f76263,
        64'hffec871b_481c0184,
        64'h2c836000_000a1c63,
        64'h00050a1b_e7cfe0ef,
        64'hec66f062_f45efc56,
        64'he4cee8ca_eca6f486,
        64'he0d28522_002c4601,
        64'h8b2ee42a_f85a8432,
        64'hf0a27159_bfcd4419,
        64'h80826165_64e67406,
        64'h70a68522_c10fe0ef,
        64'h102885a6_c489cf81,
        64'h6786e801_0005041b,
        64'h872ff0ef_e4be1028,
        64'h083c65a2_e00d0005,
        64'h041bedaf_e0eff486,
        64'hf0a21028_002c4601,
        64'h84aee42a_eca67159,
        64'hbf6584aa_d16dbf7d,
        64'h00042a23_00f51663,
        64'h47912501_f8bfe0ef,
        64'h85224581_c68fe0ef,
        64'h852285ca_00042a23,
        64'h02f51363_47912501,
        64'hb32ff0ef_85224581,
        64'h02243023_80826145,
        64'h64e26942_85267402,
        64'h70a20005_049bc5ff,
        64'he0ef8522_45810009,
        64'h1f63e889_0005049b,
        64'hd98fe0ef_892e842a,
        64'hf406e84a_ec26f022,
        64'h71798082_01416402,
        64'h60a20004_3023e119,
        64'h2501dbaf_e0ef842a,
        64'he406e022_1141b7c1,
        64'hfcf501e3_4791bfdd,
        64'h45258082_61217442,
        64'h70e2f971_fcf50be3,
        64'h47912501_cbdfe0ef,
        64'h00f41423_0067d783,
        64'h85224581_67e2c448,
        64'he30fe0ef_0007c503,
        64'h67e2a02d_00043023,
        64'h4515e789_8bc100b5,
        64'hc783cd99_6c0ce529,
        64'h250197cf_f0eff01c,
        64'h101ce01c_852265a2,
        64'h67e2e115_2501fe6f,
        64'he0ef0828_002c4601,
        64'h842ac52d_e42ef822,
        64'hfc067139_b7bdc45c,
        64'h013787bb_413484bb,
        64'hcc0c445c_faf5fae3,
        64'h4f9c601c_fabafee3,
        64'hfd4588e3_0005059b,
        64'hc4bfe0ef_bf6984ce,
        64'he5990005_059bfddf,
        64'he0efcb81_8b896008,
        64'h00a44783_b765cc0c,
        64'hc84cb5ed_490500f4,
        64'h05a34785_00f59763,
        64'h57fdbded_490900f4,
        64'h05a34789_00f59763,
        64'h47850005_059b814f,
        64'hf0efe595_484cbfb1,
        64'h9ca90094_d49bcd11,
        64'h2501c87f_e0ef6008,
        64'hd7b51ff4_f793c45c,
        64'h9fa5445c_0499ea63,
        64'h4a855a7d_d1c19c9d,
        64'hc45c2781_4c0c8ff9,
        64'h413007bb_02c6ed63,
        64'h0337563b_0336d6bb,
        64'hfff4869b_377dc729,
        64'h0097999b_00254783,
        64'h6008bf59_cc44ed35,
        64'h25012bd0_40ef85ce,
        64'h0017c503_86264685,
        64'h601c00f4_0523fbf7,
        64'hf79300a4_4783ed51,
        64'h250130f0_40ef0017,
        64'hc50385ce_4685601c,
        64'hc3850407_f7930304,
        64'h099300a4_4783fc96,
        64'h0ee34c50_d3e51ff7,
        64'hf793445c_4481bf7d,
        64'h00f40523_0207e793,
        64'h00a44783_c81cfcf7,
        64'h78e34818_445ce4bd,
        64'h00042623_445884ba,
        64'he3918b89_00a44783,
        64'h00977763_48188082,
        64'h61216aa2_6a4269e2,
        64'h790274a2_854a7442,
        64'h70e20007_891bcf89,
        64'h00b44783_00091763,
        64'h0005091b_fb4fe0ef,
        64'h84ae842a_e456e852,
        64'hec4efc06_f04af426,
        64'hf8227139_b709fe94,
        64'h65e3fee7_8fa32405,
        64'h07850007_47039736,
        64'h92810204_16936722,
        64'h0789bddd_4545b7e9,
        64'h00c68023_377dfc96,
        64'h4603962a_10889201,
        64'h02071613_b7c12785,
        64'hb7319c3d_01368023,
        64'hfff7c793_01271a63,
        64'h96b29201_66a20206,
        64'h961300e5_86bb40f4,
        64'h05bbfff7_871b04e4,
        64'h62630037_871beb05,
        64'hfc974703_97361094,
        64'h93010207_97134781,
        64'hf5cfe0ef_1828100c,
        64'hb7594509_f8e516e3,
        64'h67a24711_dd612501,
        64'ha9eff0ef_18284581,
        64'h01450e63_25018a7f,
        64'he0ef0007_c50365c6,
        64'h77e2e105_2501e48f,
        64'hf0ef1828_4581f949,
        64'h2501f63f_e0ef1828,
        64'h4581c2aa_8cdfe0ef,
        64'h0007c503_65c677e2,
        64'hf5552501_e6eff0ef,
        64'h18284581_fd452501,
        64'hf89fe0ef_18284585,
        64'h80826149_7a0679a6,
        64'h794674e6_640a60aa,
        64'h00078023_078d00e7,
        64'h812302f0_07130e94,
        64'h186300e7_80a303a0,
        64'h071300e7_80230307,
        64'h071b3427_47030000,
        64'h8717e505_67a24501,
        64'h040a1263_4a16c2be,
        64'h02f00993_4bdc597d,
        64'h842677e2_ecbe081c,
        64'he5292501_acdfe0ef,
        64'h1828002c_460184ae,
        64'h00050023_f0d2f4ce,
        64'hf8cae122_e506e42a,
        64'hfca67175_bfd94415,
        64'hfcf41ee3_4791b7c5,
        64'hc8c897bf_e0ef0004,
        64'hc50374a2_cb998bc1,
        64'h00b5c783_80826165,
        64'h64e67406_70a68522,
        64'hcbd85752_77a2e991,
        64'h6586e41d_0005041b,
        64'hcd2ff0ef_e4be1028,
        64'h083c65a2_ec190005,
        64'h041bb3bf_e0efeca6,
        64'hf486f0a2_1028002c,
        64'h4601e42a_7159bfe5,
        64'h452d8082_610560e2,
        64'h45013ea7_8d230000,
        64'h87970005_4a6395bf,
        64'he0efec06_0028e42a,
        64'h11018082_01416402,
        64'h60a20004_3023e119,
        64'h25019cbf_e0ef8522,
        64'he9012501_effff0ef,
        64'h842ae406_e0221141,
        64'h80820141_640260a2,
        64'h4505ebbf_e06f0141,
        64'h60a26402_00f50223,
        64'h478500f4_0523fdf7,
        64'hf7936008_00a44783,
        64'h000789a3_00078923,
        64'h00e78ca3_00d78da3,
        64'h04600713_0086d69b,
        64'h00e78c23_02100713,
        64'h0106d69b_00e78aa3,
        64'h0087571b_0107571b,
        64'h0107171b_00e78a23,
        64'h27010107_571b0107,
        64'h169b00e7_8d230007,
        64'h8ba30007_8b234858,
        64'h00e78fa3_00d78f23,
        64'h0187571b_0107569b,
        64'h00d78ea3_00e78e23,
        64'h0086d69b_0106d69b,
        64'h0107169b_481800e7,
        64'h85a30207_671300b7,
        64'hc703741c_e15d2501,
        64'hb77fe0ef_6008500c,
        64'h00f40523_fbf7f793,
        64'h00a44783_ed552501,
        64'h685040ef_03040593,
        64'h0017c503_46854c50,
        64'h601cc395_0407f793,
        64'hcf690207_f71300a4,
        64'h4783e175_2501acff,
        64'he0ef842a_e406e022,
        64'h1141bd2d_499db5f9,
        64'hc81cbf41_00f40523,
        64'h0407e793_00a44783,
        64'h9dbfe0ef_952285d2,
        64'h86260305_05130007,
        64'h849b0127_f46340ab,
        64'h87bb1ff5_75130009,
        64'h049b4448_01a42e23,
        64'hfd092501_6c7040ef,
        64'h85da4685_001dc503,
        64'h00e7fa63_445c4818,
        64'h00c78e63_4c5cbdd1,
        64'h00faa023_9fa5000a,
        64'ha783c45c_9fa54099,
        64'h093b445c_9a3e9381,
        64'h02049793_0094949b,
        64'h00f40523_fbf7f793,
        64'h00a44783_a4ffe0ef,
        64'h855a95d2_20000613,
        64'h91811582_0097959b,
        64'h0297f263_41a587bb,
        64'h4c4cf151_25017630,
        64'h40ef85d2_86a6001d,
        64'hc5034197_04bb00f7,
        64'h74639fb5_002dc703,
        64'hc4b58d32_0007849b,
        64'h00a6863b_0099579b,
        64'h000c869b_d1592501,
        64'h97cff0ef_856e4c0c,
        64'h00043d83_00f40523,
        64'hfbf7f793_00a44783,
        64'hf9692501_7b1040ef,
        64'h85da0017_c5034685,
        64'h4c50601c_c38d0407,
        64'hf79300a4_4783c85c,
        64'he311cc1c_4858bf99,
        64'h498500f4_05a34785,
        64'h01879763_b79500f4,
        64'h05230207_e79300a4,
        64'h478312f7_6a634818,
        64'h445cf3fd_0005079b,
        64'hd86ff0ef_4c0cb759,
        64'h498900f4_05a34789,
        64'h02e79863_4705cb91,
        64'h4581485c_ef01040c,
        64'h9a630ffc_fc930197,
        64'hfcb337fd_00254783,
        64'h00975c9b_60081407,
        64'h93631ff7_77930409,
        64'h04634458_5c7d0304,
        64'h0b132000_0b9304f7,
        64'h6c630127_873b445c,
        64'h18078f63_8b8900a4,
        64'h47838082_61656da2,
        64'h6d426ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h694664e6_854e7406,
        64'h70a60007_899bc39d,
        64'h00b44783_00099763,
        64'h0005099b_cb5fe0ef,
        64'h8ab68932_8a2e842a,
        64'h0006a023_e46ee86a,
        64'hec66f062_f45ef85a,
        64'heca6f486_fc56e0d2,
        64'he4cee8ca_f0a27159,
        64'hb59d499d_bf9dbd1f,
        64'he0ef8552_95a28626,
        64'h03058593_0007849b,
        64'h0127f463_40bb87bb,
        64'h1ff5f593_0009049b,
        64'h444c01a4_2e23f115,
        64'h25010bc0_50ef85da,
        64'h0017c503_863a4685,
        64'h601c00f4_0523fbf7,
        64'hf7936722_00a44783,
        64'hf1392501_110050ef,
        64'he43a85da_4685001d,
        64'hc503c38d_0407f793,
        64'h00a44783_04e60163,
        64'h4c50b705_00faa023,
        64'h9fa5000a_a783c45c,
        64'h9fa54099_093b445c,
        64'h9a3e9381_02049793,
        64'h0094949b_c5ffe0ef,
        64'h955285da_20000613,
        64'h91011502_0097951b,
        64'h0097fc63_41a507bb,
        64'h4c48c385_0407f793,
        64'h00a44783_f94d2501,
        64'h14a050ef_85d2863a,
        64'h86a6001d_c5034196,
        64'h84bb00f6_f4639fb1,
        64'h002dc683_c4b58d3a,
        64'h0007849b_00a6073b,
        64'h0099579b_000c861b,
        64'hd5792501_b98ff0ef,
        64'h856e4c0c_00043d83,
        64'hcc08b7a5_498500f4,
        64'h05a34785_01851763,
        64'hb7e52501_bd6ff0ef,
        64'h4c0cb741_498900f4,
        64'h05a34789_00a7ec63,
        64'h47854848_eb11020c,
        64'h99630ffc_fc930197,
        64'hfcb337fd_00254783,
        64'h00975c9b_60081207,
        64'h90631ff7_77934458,
        64'hfa090ce3_5c7d0304,
        64'h0b132000_0b930006,
        64'h091b00f6_7463893e,
        64'h40f907bb_445c0104,
        64'h29031607_89638b85,
        64'h00a44783_80826109,
        64'h6de27d02_7ca27c42,
        64'h7be26b06_6aa66a46,
        64'h69e67906_74a6854e,
        64'h744670e6_0007899b,
        64'hc39d6622_00b44783,
        64'h00099863_0005099b,
        64'he91fe0ef_8ab6e432,
        64'h8a2e842a_0006a023,
        64'hec6ef06a_f466f862,
        64'hfc5ee0da_f0caf4a6,
        64'hfc86e4d6_e8d2ecce,
        64'hf8a27119_b7d5491d,
        64'hb7e54911_80826149,
        64'h6b466ae6_7a0679a6,
        64'h794674e6_854a640a,
        64'h60aa00f4_94230134,
        64'hb0230004_ae230004,
        64'ha623c888_0069d783,
        64'hdbbfe0ef_01c40513,
        64'hc8c8f33f_e0ef0009,
        64'hc5030004_85a3d09c,
        64'h01448523_f4800309,
        64'ha78385a2_79a2020a,
        64'h6a13c399_008a7793,
        64'he3ad8b85_00098463,
        64'h0029f993_e72d0107,
        64'hf71300b4_4783f565,
        64'ha0854921_f60981e3,
        64'h0049f993_e3d98bc5,
        64'h00b44783_a895892a,
        64'hc90d2501_83aff0ef,
        64'h01352623_85da39fd,
        64'h7522e911_2501e3ff,
        64'hf0ef030a_ab038556,
        64'h85ce0409_8b6300fa,
        64'h82230005_099b0004,
        64'h0aa30004_0a230004,
        64'h0da30004_0d234785,
        64'hfc9fe0ef_85a2000a,
        64'hc5030004_0fa30004,
        64'h0f230004_0ea30004,
        64'h0e230004_05a300e4,
        64'h0c230004_0ba30004,
        64'h0b2300e4_08230004,
        64'h07a30004_072300f4,
        64'h0ca300f4_08a30210,
        64'h07130460_07937aa2,
        64'hcfcd008a_77936406,
        64'he949008a_6a132501,
        64'he75ff0ef_102800f5,
        64'h16634791_c54dc3e1,
        64'h01f9fa13_01c9f793,
        64'h4519e011_e1196406,
        64'h2501b6df_f0efe4be,
        64'h1028083c_65a21409,
        64'h10630005_091b9d6f,
        64'hf0ef1028_002c8a79,
        64'h84aa89b2_00053023,
        64'h14050d63_4925e42e,
        64'he8daecd6_f0d2f4ce,
        64'hfca6e122_e506f8ca,
        64'h7175bfe5_452d8082,
        64'h612170e2_2501a0ef,
        64'hf0ef0828_080c4601,
        64'h00f61863_4785cb11,
        64'h4501e398_97aa0007,
        64'h0023c319_67620007,
        64'h0023c319_66226318,
        64'h00a78733_050eace7,
        64'h87930000_97970405,
        64'h426383ef_f0eff42e,
        64'he432e82e_fc061028,
        64'hec2a7139_b7594505,
        64'hbf5d0009_049b00f4,
        64'h02a30017_e7930054,
        64'h4783c81c_27850137,
        64'h8a63481c_f15d2501,
        64'h8afff0ef_852285a6,
        64'h46010339_0763fb49,
        64'h0ce3bf75_45010009,
        64'h14630005_091bec8f,
        64'hf0ef8522_85a600f4,
        64'hfa634c1c_59fd4a05,
        64'hfcf5fde3_84ae842a,
        64'he052e44e_e84af406,
        64'hec26f022_71794d1c,
        64'h80826145_6a0269a2,
        64'h694264e2_740270a2,
        64'h45098082_450900b7,
        64'hed634785_80826105,
        64'h64a28526_644260e2,
        64'h00e78223_4705601c,
        64'h82aff0ef_462d6c08,
        64'h700c84cf_f0ef4581,
        64'h02000613_6c08e085,
        64'h0005049b_a42ff0ef,
        64'h6008484c_e49d0005,
        64'h049bfa9f_f0ef842a,
        64'hec06e426_e8221101,
        64'h80826105_64a26442,
        64'h60e2451d_00f51363,
        64'h4791dd79_2501bcdf,
        64'hf0ef8522_4585cb99,
        64'h00978d63_0007c783,
        64'h6c1ced09_2501a8cf,
        64'hf0ef6008_484c0e50,
        64'h0493e50d_250188ff,
        64'hf0ef842a_e426ec06,
        64'he8224581_1101bfe5,
        64'h4511b7cd_00042a23,
        64'hd9452501_c13ff0ef,
        64'h85224581_80826145,
        64'h69a26942_64e27402,
        64'h70a24501_00979a63,
        64'h0017b793_17e18bfd,
        64'h03378063_03270263,
        64'h03f7f793_00b7c783,
        64'hc3210007_c7036c1c,
        64'he1292501_afaff0ef,
        64'h6008a0b1_c90de199,
        64'h484c49bd_0e500913,
        64'h451184ae_f406842a,
        64'he44ee84a_ec26f022,
        64'h7179bdf9_0ff77713,
        64'h0017e793_3701eea8,
        64'h66e30ff5_7513f9f7,
        64'h051beea8_7ae30ff5,
        64'h7513fbf7_051bbd6d,
        64'h4519f117_10e30008,
        64'h86630005_4883ece5,
        64'h05130000_85170005,
        64'h4c634185_551b0187,
        64'h151b02b6_f263fd37,
        64'h0ae3f957_04e3f947,
        64'h06e3f4e3_74e30007,
        64'h47039722_93011702,
        64'h0017061b_873245ad,
        64'h46a10ff7_f7930027,
        64'h979b0565_9a63bdb9,
        64'hc4c8af2f_f0ef0007,
        64'hc503609c_dbe58bc1,
        64'h00b5c783_6c8cfbf5,
        64'h8b91b73d_4515fb0d,
        64'hbf154501_e80703e3,
        64'h0004bc23_0004a623,
        64'hcb890207_f7930047,
        64'hf713f4e5_18e34711,
        64'hc50500b7_c783709c,
        64'h4511bf65_4701bdfd,
        64'h00e905a3_94329201,
        64'h16020087_671300d7,
        64'h94634691_8bb10107,
        64'h671300b6_94634585,
        64'h0037f693_0ff7f793,
        64'h0027979b_01659663,
        64'h00d90023_469500d5,
        64'h15630e50_06930009,
        64'h4503c6ed_4711a06d,
        64'h268500e5_0023954a,
        64'h91010206_95130027,
        64'he793a8dd_0505a0d1,
        64'h48650200_03134781,
        64'h45a14701_4681b7ad,
        64'h02400793_943a12f6,
        64'he0630200_0693f757,
        64'h8be3bf95_4709bf1d,
        64'h04058082_61216b02,
        64'h6aa26a42_69e27902,
        64'h74a27442_70e20004,
        64'hbc232501_a85ff0ef,
        64'h85264581_b791c55c,
        64'h4bdc611c_bf75dfdf,
        64'hf0ef8526_4581fed6,
        64'h08e3fff7_c683fff7,
        64'h46030785_07050cb7,
        64'h8d6300b7_8593709c,
        64'hef918ba1_00b74783,
        64'hc7e50007_47836c98,
        64'he96d2501_cdaff0ef,
        64'h608848cc_10051063,
        64'h2501adbf_f0ef8526,
        64'h458100f9_05a30200,
        64'h0793943a_09479763,
        64'h470d1b37_8e630024,
        64'h478300f9_00a302e0,
        64'h07930b37_90630014,
        64'h47830139_00230d37,
        64'h92630004_4783b40f,
        64'hf0ef854a_02000593,
        64'h462d0204_b9030d57,
        64'h80630d47_82630004,
        64'h47834b21_02e00993,
        64'h05c00a93_02f00a13,
        64'h0ae7fc63_47fd0004,
        64'h47030004_a6230405,
        64'h0ce79063_05c00713,
        64'h00e78663_842e84aa,
        64'h02f00713_0005c783,
        64'he05ae456_e852ec4e,
        64'hf04afc06_f426f822,
        64'h7139b7e9_db1c2785,
        64'h5b1c2a85_6018f141,
        64'h2501d1cf_f0ef0145,
        64'h0223b7b9_c848a83f,
        64'hf0ef85a6_c8046008,
        64'hd91c4157_87bb591c,
        64'h00faed63_00254783,
        64'h60084a05_02aa2823,
        64'haa5ff0ef_855285a6,
        64'h00043a03_beeff0ef,
        64'h03450513_45812000,
        64'h06136008_f5792501,
        64'hdd8ff0ef_6008fcf4,
        64'h8de357fd_fcf48be3,
        64'h4785d4bd_451d0005,
        64'h049be81f_f0ef480c,
        64'hf60a0ee3_06f4e063,
        64'h4d1c6008_b7614505,
        64'h00f49463_57fdbf49,
        64'h45090097_e4634785,
        64'h0005049b_b27ff0ef,
        64'hfc0a9fe3_0157fab3,
        64'h37fd0049_5a9b0025,
        64'h4783bf5d_4501ec1c,
        64'h97ce0347_87930124,
        64'h15230996_601cfcf7,
        64'h75e30009_071b0085,
        64'h5783e18d_c85c6108,
        64'h2785480c_00099d63,
        64'h842a8a2e_00f97993,
        64'hd7ed495c_80826121,
        64'h6aa26a42_69e27902,
        64'h74a27442_70e24511,
        64'heb9993c1_e456e852,
        64'hec4ef426_03091793,
        64'h2905f822_fc0600a5,
        64'h5903f04a_7139bfad,
        64'h4405f6f5_0fe34785,
        64'hdd612501_dbbff0ef,
        64'h852685ce_8622bf49,
        64'h00f482a3_0017e793,
        64'h0054c783_c89c37fd,
        64'hfae783e3_577dc4c0,
        64'h489c0209_9063e905,
        64'h2501de9f_f0ef8526,
        64'h85a2167d_10000637,
        64'hb76dfb24_11e30545,
        64'h0863fd55_07e3c901,
        64'h2501c05f_f0ef8526,
        64'h85a24409_bf554905,
        64'hb7d5faf4_7ee3894e,
        64'h4c9c8082_61216aa2,
        64'h6a4269e2_790274a2,
        64'h744270e2_8522547d,
        64'h00f41d63_57fd0887,
        64'hf8634785_0005041b,
        64'hc43ff0ef_a8214401,
        64'h052a6063_04f46363,
        64'h24054c9c_5afd4a05,
        64'h844a04f9_77634d1c,
        64'h04090a63_00c52903,
        64'he19d89ae_84aae456,
        64'he852f04a_f822fc06,
        64'hec4ef426_7139bf3d,
        64'h4989b745_012a81a3,
        64'h00fa8123_0189591b,
        64'h0109579b_00fa80a3,
        64'h0087d79b_03240a23,
        64'h0107d79b_94260109,
        64'h179b0125_69338d71,
        64'hf0000637_2501da0f,
        64'hf0ef8556_9aa60344,
        64'h0a931fc4_74130024,
        64'h141bf809_96e30005,
        64'h099bfd8f_f0ef9dbd,
        64'h0075d59b_515cbf79,
        64'h01448223_03240aa3,
        64'h0089591b_0109591b,
        64'h0109191b_03240a23,
        64'h94261fe4_74130014,
        64'h141bfc09_92e30005,
        64'h099b811f_f0ef9dbd,
        64'h0085d59b_515cb7e9,
        64'h0127e933_9bc100f9,
        64'h79130089_591b0347,
        64'hc7830154_87b38082,
        64'h61216aa2_6a4269e2,
        64'h790274a2_854e7442,
        64'h70e200f4_82234785,
        64'h032a8a23_9aa60ff9,
        64'h79130049_591bc40d,
        64'h1ffafa93_00099f63,
        64'h0005099b_86bff0ef,
        64'h9dbd8526_009ad59b,
        64'h50dc00f4_82234785,
        64'h02fa0a23_9a260ff7,
        64'hf7938fd9_8ff50049,
        64'h179b00f7_f71316c1,
        64'h66850347_c7830144,
        64'h87b3cc19_1ffa7a13,
        64'h0ff97793_001a0a9b,
        64'h88050609_96630005,
        64'h099b8b9f_f0ef9dbd,
        64'h009a559b_00ba0a3b,
        64'h515c0015_da1b1547,
        64'h94630ee7_8863470d,
        64'h0ae78f63_842e8932,
        64'h47090005_47830af5,
        64'hf0634989_84aa4d1c,
        64'h16ba7563_4a05e456,
        64'hec4ef04a_f426f822,
        64'hfc06e852_71398082,
        64'h610564a2_85266442,
        64'h60e200e7_82234705,
        64'h601c00e7_80235715,
        64'h6c1cf3cf_f0ef4581,
        64'h02000613_6c08ec99,
        64'h0005049b_933ff0ef,
        64'h6008484c_e4950005,
        64'h049bf33f_f0ef842a,
        64'hec06e426_e8221101,
        64'h00a55583_b78d4505,
        64'hbfc14134_84bbf6f4,
        64'h76e34f9c_00093783,
        64'hf68afbe3_01440c63,
        64'h0005041b_e6fff0ef,
        64'hbf752501_e59ff0ef,
        64'h0134f663_85a20009,
        64'h35034a85_09925a7d,
        64'h843a0027_c9838722,
        64'hb75d4501_00993c23,
        64'h00a92a23_94be0347,
        64'h87930496_88bd0009,
        64'h37839d3d_0044d79b,
        64'hd1710089_28235788,
        64'hfce4f7e3_0087d703,
        64'heb155798_00e69463,
        64'h470d0007_c683e021,
        64'h84aefee4_74e34f98,
        64'h611c8082_61216aa2,
        64'h6a4269e2_790274a2,
        64'h744270e2_450900f4,
        64'h1c63892a_478500b5,
        64'h1523e456_e852ec4e,
        64'hf426fc06_f04a4540,
        64'hf8227139_8082853e,
        64'h4785b765_17fd2501,
        64'h100007b7_807ff0ef,
        64'h954a0345_05131fc5,
        64'h75130024_151bf935,
        64'h2501a39f_f0ef9dbd,
        64'h0075d59b_515cb759,
        64'h8fc90087_979b0349,
        64'h45030359_47839922,
        64'h1fe47413_0014141b,
        64'hfd592501_a63ff0ef,
        64'h9dbd0085_d59b515c,
        64'hbf458fe9_157d6505,
        64'hbf658391_c0198fc5,
        64'h0087979b_88050349,
        64'h4783994e_1ff9f993,
        64'hf5792501_a93ff0ef,
        64'h0344c483_854a9dbd,
        64'h94ca1ff4_f4930099,
        64'hd59b0014_899b0249,
        64'h27838082_6145853e,
        64'h69a26942_64e27402,
        64'h70a257fd_c9112501,
        64'hac7ff0ef_9dbd0094,
        64'hd59b9cad_515c0015,
        64'hd49b00f7_1e6308d7,
        64'h0e63468d_06d70c63,
        64'h842e4689_00054703,
        64'h02e5f963_892ae44e,
        64'hec26f022_f406e84a,
        64'h71794d18_0eb7f763,
        64'h47858082_45018082,
        64'h9d2d02d5_85bb5548,
        64'h00254583_00f6f963,
        64'h37f9ffe5_869b4d1c,
        64'h80826105_64a26442,
        64'h60e200a0_35332501,
        64'h631050ef_45814601,
        64'h00144503_000402a3,
        64'h63d050ef_85a64685,
        64'hd81022f4_01a322e4,
        64'h012320d4_0ca320d4,
        64'h0c230187_d79b0107,
        64'hd71b2605_22e400a3,
        64'h22f40023_07200693,
        64'h00144503_0087571b,
        64'h0107571b_0107971b,
        64'h501020e4_0f23445c,
        64'h20f40fa3_0187d79b,
        64'h0107d71b_20e40ea3,
        64'h20f40e23_0087571b,
        64'h0107571b_0107971b,
        64'h20e40d23_02e40ba3,
        64'h04100713_481c20f4,
        64'h0da302f4_0b230610,
        64'h079302f4_0aa302f4,
        64'h0a230520_079322f4,
        64'h09a3faa0_079322f4,
        64'h09230550_0793a01f,
        64'hf0ef8526_45812000,
        64'h06130344_04930af7,
        64'h1b634785_00544703,
        64'h0cf71063_478d0004,
        64'h4703ed69_2501bfff,
        64'hf0ef842a_e426ec06,
        64'he8221101_bdc59cbd,
        64'h0017d79b_88850297,
        64'h87bb478d_b7010014,
        64'h949b00f9_15634789,
        64'hd41c9fb5_e00a05e3,
        64'hb545a25f_f0ef0544,
        64'h0513b5b9_0005099b,
        64'ha33ff0ef_05840513,
        64'hb3514781_00042a23,
        64'h01240023_00f41323,
        64'h5cf71d23_00009717,
        64'h93c117c2_27855e87,
        64'hd7830000_9797c448,
        64'ha63ff0ef_22040513,
        64'hc808a6df_f0ef21c4,
        64'h051300f5_1c632727,
        64'h87932501_614177b7,
        64'ha83ff0ef_21840513,
        64'h02f51763_25278793,
        64'h25014161_57b7a99f,
        64'hf0ef0344_051304f7,
        64'h1263a557_07134107,
        64'hd79b776d_0107979b,
        64'h8fd90087_979b0004,
        64'h02a32324_47032334,
        64'h4783e13d_2501ce5f,
        64'hf0ef8522_001a859b,
        64'h06f71b63_47054107,
        64'hd79b0107_979b8fd9,
        64'h0087979b_06444703,
        64'h06544783_08f91963,
        64'h478d00f4_02a3f800,
        64'h0793c45c_c81c57fd,
        64'hee99e7e3_24810094,
        64'hd49b1ff4_849b0024,
        64'h949bd408_b17ff0ef,
        64'h06040513_f00a15e3,
        64'h10e91263_470dd05c,
        64'h03542023_cc04d458,
        64'h015787bb_248900ea,
        64'h873b490d_00b67363,
        64'h09051655_00b93933,
        64'h66411955_6905dd8d,
        64'h84ae0364_d5bb40c5,
        64'h04bbf4c5_64e38732,
        64'h00d7063b_9f3d004a,
        64'h571b2781_033906bb,
        64'hdfb18fd9_0087979b,
        64'h25010424_47030434,
        64'h47831405_0e638d45,
        64'h0085151b_04744483,
        64'h04844503_f3c100fa,
        64'h77930144_142300fa,
        64'h6a33008a_1a1b0454,
        64'h47830464_4a03ffc9,
        64'h00fb77b3_fffb079b,
        64'hfa0b03e3_01640123,
        64'h04144b03_faf769e3,
        64'h0ff7f793_012401a3,
        64'hfff9079b_47050134,
        64'h2e230444_49032981,
        64'h1a098663_00f9e9b3,
        64'h0089999b_04a44783,
        64'h04b44983_fef711e3,
        64'h20000713_4107d79b,
        64'h0107979b_8fd90087,
        64'h979b03f4_47030404,
        64'h4783bfb9_47b5c119,
        64'h4a81f6e5_04e34785,
        64'h470db7bd_00e51963,
        64'h4785470d_fe9915e3,
        64'h0491c10d_e9dff0ef,
        64'h852285d6_000a8763,
        64'h45090004_aa830104,
        64'h8913ff2a_14e30991,
        64'h094100a9_a0232501,
        64'hc5bff0ef_854ac789,
        64'h4501ffc9_478389a6,
        64'h23a40a13_1fa40913,
        64'h848a04f5_1a634785,
        64'hee1ff0ef_85224581,
        64'hf5698911_00090463,
        64'hfb71478d_00157713,
        64'h0f4060ef_00a400a3,
        64'h00040023_0ff4f513,
        64'h80826161_853e6b42,
        64'h6ae27a02_79a27942,
        64'h74e26406_60a647a9,
        64'hc1118911_00090563,
        64'he38d0015_77931e20,
        64'h60ef0014_4503cb85,
        64'h00044783_0089b023,
        64'hc01547b1_84aa6380,
        64'h97ba8627_87930000,
        64'ha7970035_17130205,
        64'h4e6347ad_dd9ff0ef,
        64'h8932852e_89aa0005,
        64'h3023e85a_ec56f052,
        64'hfc26e0a2_e486f44e,
        64'hf84a715d_bfcd450d,
        64'h80826105_690264a2,
        64'h644260e2_00a03533,
        64'h8d050125_75332501,
        64'hd33ff0ef_08640513,
        64'h00978c63_45010127,
        64'hf7b31465_04930054,
        64'h4537fff5_09130100,
        64'h05370005_079bd59f,
        64'hf0ef06a4_051302f7,
        64'h1f63a557_07134107,
        64'hd79b776d_0107979b,
        64'h8fd90087_979b4509,
        64'h23244703_23344783,
        64'he52d2501_fa3ff0ef,
        64'h842ad91c_00050223,
        64'h57fde04a_e426ec06,
        64'he8221101_80826105,
        64'h690264a2_644260e2,
        64'h85220324_a823597d,
        64'h4405c119_25012980,
        64'h60ef0344_8593864a,
        64'h46850014_c503ec19,
        64'h0005041b_fddff0ef,
        64'h892e84aa_02b78763,
        64'h4401e04a_e426ec06,
        64'he8221101_591c8082,
        64'h4501f8df_f06fc399,
        64'h00454783_b7f94505,
        64'hb7e5397d_310060ef,
        64'h85ce8626_9cbd4685,
        64'h00144503_4c5cff2a,
        64'h74e34a05_00344903,
        64'h80826145_6a0269a2,
        64'h694264e2_740270a2,
        64'h450100e7_eb6340f4,
        64'h87bb0004_02234c58,
        64'h505ce131_25013520,
        64'h60ef85ce_86264685,
        64'h00154503_842a0345,
        64'h0993e052_e84af406,
        64'h5904e44e_ec26f022,
        64'h71798082_853e2781,
        64'h8fd90107_979b8fd5,
        64'h0087979b_0145c683,
        64'h0155c783_00d51d63,
        64'h0007079b_8f5d0087,
        64'h979b468d_01a5c703,
        64'h01b5c783_80824525,
        64'h80820141_60a24525,
        64'hc3914501_00157793,
        64'h3c4060ef_0017c503,
        64'he4061141_02e69063,
        64'h00855703_0067d683,
        64'hc70d0007_c703cb85,
        64'h611cc915_bfd5a5e7,
        64'h47030000_a7178082,
        64'h853ae11c_0006871b,
        64'h078900b6_66630ff6,
        64'hf593fd06_869b577d,
        64'h46050007_c683b7dd,
        64'h0705a00d_577d00d7,
        64'h06630017_869300c6,
        64'h986302d5_fc630007,
        64'h468303a0_06130200,
        64'h0593cf99_873e611c,
        64'h80826105_690264a2,
        64'h644260e2_00040023,
        64'h00f49323_8fd90087,
        64'h979b0169_47030179,
        64'h478300f4_92238fd9,
        64'h0087979b_01894703,
        64'h01994783_c088f59f,
        64'hf0ef00f5_842384ae,
        64'h01c90513_00b94783,
        64'hfcc79ee3_06850405,
        64'h00e40023_04050064,
        64'h00230117_95630e50,
        64'h07130107_146300a7,
        64'h0e632785_0006c703,
        64'h462d02e0_031348a5,
        64'h481586ca_02000513,
        64'h47810185_3903cfa5,
        64'h00958413_e04ae426,
        64'hec06e822_1101495c,
        64'hbfcd0505_00b50023,
        64'h808200f6_1363367d,
        64'h57fdb7f5_fee50fa3,
        64'h05850505_0005c703,
        64'h808200f6_1363367d,
        64'h57fd8082_25018d5d,
        64'h05628fd9_07c20035,
        64'h45030025_47838f5d,
        64'h07a20005_47030015,
        64'h4783b7d9_14fdb7e9,
        64'hba9ff0ef_bfc1710a,
        64'h849377d0_50ef4501,
        64'hdff154fd_000a2783,
        64'hbfc5bc3f_f0effc07,
        64'h5de30337_97138309,
        64'h37830207_45630337,
        64'h97138309_37835a0b,
        64'h0493ee5f_e0ef8522,
        64'he78d0009_a783e4a9,
        64'hb807ac23_0000a797,
        64'hba07a223_0000a797,
        64'hba07a823_0000a797,
        64'hba07a423_0000a797,
        64'hba079a23_0000a797,
        64'hbcf70ea3_0000a717,
        64'h00544783_bef70423,
        64'h0000a717_00444783,
        64'hbef709a3_0000a717,
        64'h00344783_bef70f23,
        64'h0000a717_30001937,
        64'h00262b37_00244783,
        64'hc0f708a3_0000a717,
        64'h6a89c02a_0a130000,
        64'haa170014_4783c2f7,
        64'h03230000_a717c0e9,
        64'h89930000_a9974481,
        64'h00044783_c3440413,
        64'h0000a417_07d030ef,
        64'he5050513_00009517,
        64'hc485c583_0000a597,
        64'hc5164603_0000a617,
        64'hc5a6c683_0000a697,
        64'hc6584803_0000a817,
        64'hc6c7c783_0000a797,
        64'hc7374703_0000a717,
        64'h0b9030ef_e7c50513,
        64'h00009517_80e7b423,
        64'he05ae456_e852ec4e,
        64'hf04af426_f822fc06,
        64'h8f4d91c1_15c20080,
        64'h07377139_8087b583,
        64'h8007b603_300017b7,
        64'hbf91ff34_10e30f70,
        64'h30effec4_8fa30ff6,
        64'h761300c9_56330286,
        64'h061b0485_24058552,
        64'h85a2028a_863b4999,
        64'hec0a0a13_00009a17,
        64'h5ae14401_ce448493,
        64'h0000a497_80826161,
        64'h6ae27a02_79a27942,
        64'h74e282f6_b42347a1,
        64'h640660a6_8086b783,
        64'h8006b783_80f6b423,
        64'h93c180a6_b02317c2,
        64'h91013000_16b78fd9,
        64'h15020ff7_77138ff1,
        64'h83210087_179bf006,
        64'h06130100_06374722,
        64'hf39ff0ef_45127d00,
        64'h50ef0028_d4458593,
        64'h0000a597_46097e00,
        64'h50ef0048_d5658593,
        64'h0000a597_4611d6a7,
        64'h81a30000_a797fe05,
        64'h6513893d_003070ef,
        64'hd6f70a23_0000a717,
        64'h5791d6f7_0ea30000,
        64'ha717578d_d8f70323,
        64'h0000a717_5789d8f7,
        64'h07a30000_a7175785,
        64'hd8f70c23_0000a717,
        64'h57b90a09_1d631e70,
        64'h30eff825_05130000,
        64'h9517892a_06d070ef,
        64'hc63eec56_f052f44e,
        64'hfc26e0a2_e486f84a,
        64'h04b00513_45854601,
        64'h00740207_879b0700,
        64'h07b7715d_80822501,
        64'h8d5d8d79_00ff0737,
        64'h0085151b_8fd98f75,
        64'h0085571b_f0068693,
        64'h8fd966c1_0185579b,
        64'h0185171b_80829141,
        64'h15428d5d_05220085,
        64'h579b8082_614564e2,
        64'h740270a2_85228d4f,
        64'hf0efe225_05130000,
        64'ha5170450_0693e1a7,
        64'h57030000_a717e168,
        64'h88930000_a89785a6,
        64'h862247b2_0007a803,
        64'he3078793_0000a797,
        64'h0e3050ef_f4060068,
        64'he7858593_0000a597,
        64'h461184ae_8432ec26,
        64'hf0227179_bfc14785,
        64'heb9ff0ef_80826105,
        64'h64a26442_60e2c3c0,
        64'h0c2007b7_2c5030ef,
        64'h04850513_00009517,
        64'he7990206_c1630337,
        64'h16938304_b7033000,
        64'h14b74781_2401ec06,
        64'he42643c0_e8220c20,
        64'h07b71101_b7e1ff06,
        64'hbc2306a1_26050008,
        64'h380300d7_88338082,
        64'h61010113_5f813483,
        64'h85266001_34036081,
        64'h30838287_b8233000,
        64'h17b70405_aa1ff0ef,
        64'h862602e6_446397c2,
        64'h85b63000_08378f95,
        64'h868a83f5_02d7473b,
        64'h17822705_46a10077,
        64'h67139fad_377d8005,
        64'h859b6585_02d51a63,
        64'h80668693_6685c691,
        64'h8005069b_00015503,
        64'h00d10023_0086d69b,
        64'h0106d69b_0106969b,
        64'h00d100a3_872646d4,
        64'h96aa068e_9ebd8006,
        64'h869b7007_f7930084,
        64'h179bea25_4390f4e7,
        64'h87930000_a797cfb5,
        64'h27818ff1_fff7c793,
        64'h00c5963b_10100593,
        64'h8a1d08b8_696335b9,
        64'h5f200813_ffc5849b,
        64'h25816011_34235e91,
        64'h3c23630c_8387b783,
        64'h972a3000_05379f2d,
        64'h8406871b_03877593,
        64'h66850034_171b00f6,
        64'h74132601_60813023,
        64'h9f010113_8307b603,
        64'h300017b7_bba54601,
        64'h401030ef_16c50513,
        64'h00009517_85aab369,
        64'h00f41623_60800793,
        64'h00f41f23_0024d783,
        64'h00f41e23_0004d783,
        64'h02f41423_01e45783,
        64'h02f41323_02a00613,
        64'h01c45783_28f050ef,
        64'h852285ca_46192990,
        64'h50ef0064_05130165,
        64'h85930000_a5974619,
        64'h2ab050ef_854e0265,
        64'h85930000_a5974619,
        64'h2bb050ef_854a85ce,
        64'h461900f5_9a230165,
        64'h89930205_89132000,
        64'h0793eaf7_19e30687,
        64'hd7830000_a7970285,
        64'hd703ecf7_11e30764,
        64'h84930000_a49707e7,
        64'hd7830000_a7970265,
        64'hd703b1e1_1e450513,
        64'h00009517_b9c91d65,
        64'h05130000_9517b9f1,
        64'h1b050513_00009517,
        64'hb1dd19a5_05130000,
        64'h9517b9c5_18c50513,
        64'h00009517_b9ed16e5,
        64'h05130000_9517b311,
        64'h16850513_00009517,
        64'hb3391525_05130000,
        64'h9517bb21_14450513,
        64'h00009517_b30d12e5,
        64'h05130000_9517b335,
        64'h12850513_00009517,
        64'hb79936d0_50ef0868,
        64'h10058593_0000a597,
        64'h4611f4f7_0de30204,
        64'h5703f6f7_01e317fd,
        64'h67c101e4_5703f6e7,
        64'h87e35fe0_0713bf95,
        64'hcc6ff0ef_02a40513,
        64'h85ca5530_30ef14e5,
        64'h05130000_9517cdcf,
        64'hf0ef8522_85a65670,
        64'h30ef1525_05130000,
        64'h951702e7_98634d20,
        64'h0713b765_d6dfe0ef,
        64'h02a40513_14458593,
        64'h0000a597_14060613,
        64'h0000a617_14468693,
        64'h0000a697_f7e9439c,
        64'h15078793_0000a797,
        64'hc799439c_16078793,
        64'h0000a797_14f72e23,
        64'h0000a717_47e204e6,
        64'h94630430_07138082,
        64'h616179a2_794274e2,
        64'h640660a6_552060ef,
        64'h450102a4_0593ff89,
        64'h061b1727_87930000,
        64'ha79766a2_47624410,
        64'h50efe436_18f72e23,
        64'h0000a717_19c50513,
        64'h0000a517_19458593,
        64'h0000a597_461947e2,
        64'h1ad79e23_0000a797,
        64'h04e79b63_01c15683,
        64'h04500713_00e10e23,
        64'h02344703_00e10ea3,
        64'h01c11903_02244703,
        64'h00e10e23_27810274,
        64'h470300e1_0ea301c1,
        64'h178300f1_0e230254,
        64'h478300f1_0ea30264,
        64'h47030244_4783bdb5,
        64'h23850513_00009517,
        64'hb55922a5_05130000,
        64'h9517bd41_21c50513,
        64'h00009517_a06ddcbf,
        64'he0ef4501_85a202f4,
        64'h12238626_01c15783,
        64'h00a10e23_812100a1,
        64'h0ea3db9f_f0ef00f4,
        64'h1e230029_d78300f4,
        64'h1d230009_d78302f4,
        64'h10230224_0513fde4,
        64'h859b01c4_578300f4,
        64'h1f230204_12230204,
        64'h012301a4_57835210,
        64'h50ef854a_29c58593,
        64'h0000a597_46195310,
        64'h50ef8522_85ca4619,
        64'h10f71c63_2ce7d783,
        64'h0000a797_02045703,
        64'h12f71463_2dc98993,
        64'h0000a997_2e47d783,
        64'h0000a797_01e45703,
        64'hb73d41a5_05130000,
        64'h9517f0f5_9ce30880,
        64'h079326f5_89630ff0,
        64'h079326f5_88630890,
        64'h0793b73d_f4f58ae3,
        64'h41050513_00009517,
        64'h06c00793_26f58b63,
        64'h06700793_00b7ef63,
        64'h28f58663_08400793,
        64'hbf91f6f5_8de33fe5,
        64'h05130000_951705e0,
        64'h079328f5_846305c0,
        64'h0793b7bd_f8f58ae3,
        64'h3e850513_00009517,
        64'h03200793_28f58763,
        64'h02f00793_00b7ef63,
        64'h2af58263_03300793,
        64'h04b7e263_2cf58263,
        64'h06200793_b7c93e65,
        64'h05130000_9517faf5,
        64'h96e30290_07932af5,
        64'h86630210_0793bf6d,
        64'hfef580e3_3cc50513,
        64'h00009517_47d916f5,
        64'h8a6347c5_00b7ed63,
        64'h2cf58263_47f5a431,
        64'h7e1030ef_fef591e3,
        64'h3b050513_00009517,
        64'h47a118f5_82634799,
        64'ha41d7fb0_30ef5465,
        64'h05130000_951702f5,
        64'h83633aa5_05130000,
        64'h95174789_10f58463,
        64'h478502b7_e3631af5,
        64'h83634791_04b7e563,
        64'h1cf58263_47b108b7,
        64'he76332f5_896302e0,
        64'h07930174_45836910,
        64'h50ef3d25_05130000,
        64'ha5174619_85ca0064,
        64'h09136a50_50ef4611,
        64'h082884b2_05e94407,
        64'h9a638005_079b0af5,
        64'h0e636dd7_879367a1,
        64'h3cf50563_842e8067,
        64'h8793f44e_f84afc26,
        64'he486e0a2_6785715d,
        64'hbf55943e_00e15783,
        64'h00f10723_00d14783,
        64'h00f107a3_34f90909,
        64'h00c14783_6f7050ef,
        64'h00684609_85ca8082,
        64'h61459141_694264e2,
        64'h1542fff5_45137402,
        64'h70a29522_01045513,
        64'h942a9041_14420104,
        64'h55130290_44634401,
        64'h84ae892a_f406e84a,
        64'hec26f022_71798082,
        64'h42050513_00009517,
        64'hbf7546a5_05130000,
        64'h95178407_8793fce6,
        64'h08e346a5_05130000,
        64'h95178387_8713bfe9,
        64'h45850513_00009517,
        64'h82878793_00c74963,
        64'hfee609e3_47c50513,
        64'h00009517_83078713,
        64'h8082faf6_12e345e5,
        64'h05130000_95178187,
        64'h879300e6_0a6345e5,
        64'h05130000_95178107,
        64'h87138082_01414ce5,
        64'h05130000_a51760a2,
        64'h13c040ef_e4064de5,
        64'h05130000_a5174fe5,
        64'h85930000_95979e3d,
        64'h11417c07_879b77fd,
        64'h04c7c963_50c50513,
        64'h00009517_87f78793,
        64'h6785c3ad_48c50513,
        64'h00009517_8006079b,
        64'h04c74963_06e60b63,
        64'h4b050513_00009517,
        64'h80878713_08a74463,
        64'h862a0ce5_07638207,
        64'h87136785_8082953e,
        64'h057e4505_97aa2000,
        64'h0537e308_95360017,
        64'h86930075_6513157d,
        64'h631c57a7_07130000,
        64'ha7178082_40000537,
        64'h8082057e_4505bfb1,
        64'h24057fb0_50ef854a,
        64'h45818626_204040ef,
        64'h855e85ca_993e8626,
        64'h8c9d7902_0097ff63,
        64'h77a274c2_99828526,
        64'h0009061b_45c22260,
        64'h40ef856a_86ca85a6,
        64'h66428082_612d6d0a,
        64'h6caa6c4a_6bea7b0a,
        64'h7aaa7a4a_79ea690e,
        64'h64ae644e_60ee5575,
        64'h250040ef_50450513,
        64'h00009517_85a60397,
        64'he8630184_87b37482,
        64'h04090863_792226e0,
        64'h40ef855a_85a2cfbd,
        64'h77c20957_926347a2,
        64'h99829dbd_00280380,
        64'h06137786_028a05bb,
        64'ha0916566_00f46463,
        64'h07815783_564d0d13,
        64'h00009d17_08000cb7,
        64'h80000c37_58cb8b93,
        64'h00009b97_554b0b13,
        64'h00009b17_4a850380,
        64'h0a134401_06e79d63,
        64'h55796318_47470713,
        64'h0000a717_8ff98361,
        64'h577d6786_9982e16a,
        64'he566e962_ed5ef15a,
        64'hf556f952_e1cae5a6,
        64'he9a2ed86_00884581,
        64'h89aa0400_0613fd4e,
        64'h7115bfd5_8f8d2505,
        64'h8082e21c_00b7f463,
        64'h45019181_87aa1582,
        64'hbf390705_01070023,
        64'h0005d463_4185d59b,
        64'h0185959b_c5190975,
        64'h75130005_450300bc,
        64'h05330007_4583bfdd,
        64'h4701bf1d_3cfdfe97,
        64'h6ae32705_67220e40,
        64'h70efe43a_855eb75d,
        64'h00c58023_0ff67613,
        64'h00ea85b3_0006c603,
        64'hbf6500c5_90239241,
        64'h164295d6_00171593,
        64'h0006d603_006d1c63,
        64'hbfc1e190_95d60037,
        64'h15936290_011d1863,
        64'hbf856862_78820705,
        64'h96d27322_674266a2,
        64'h3a0040ef_e436e83a,
        64'hec42f046_f41a855a,
        64'h65829201_1602c190,
        64'h260195d6_00271593,
        64'h4290030d_1b63b795,
        64'h557dd135_0b8070ef,
        64'h99369281_168241b4,
        64'h043b66a2_3dc040ef,
        64'hfa060c23_e43667e5,
        64'h05130000_951785d6,
        64'h963e011c_0ac5ed63,
        64'h415705bb_0006861b,
        64'h02e00813_875603bd,
        64'h06bb0d9d_e66399ba,
        64'h03470733_9301020d,
        64'h971305b6_6c630007,
        64'h061b4309_48a14811,
        64'h470186ce_000c8d9b,
        64'h008cf463_00040d9b,
        64'h438040ef_6c450513,
        64'h00009517_85ca8082,
        64'h616d6daa_6d4a6cea,
        64'h7c0a7baa_7b4a7aea,
        64'h6a0e69ae_694e64ee,
        64'h740e70ae_4501e00d,
        64'h5d8c0c13_00008c17,
        64'h670b8b93_00009b97,
        64'h708b0b13_00009b17,
        64'h03810a93_020a5a13,
        64'h0017849b_e03e020d,
        64'h1a13001d_179b03ac,
        64'hdcbb4cc1_000c9563,
        64'h02ccdcbb_04000c93,
        64'h00e7f663_84368d32,
        64'h89ae892a_04000793,
        64'he56ef162_f55ef95a,
        64'hfd56e1d2_eda6f586,
        64'he96ae5ce_e9caf1a2,
        64'h02c7073b_8cbaed66,
        64'h71514da0_406f6105,
        64'h76050513_00009517,
        64'h64a26902_85a6864a,
        64'h60e26442_4f4040ef,
        64'h75850513_00009517,
        64'h85a2c801_504040ef,
        64'h89327625_05130000,
        64'h95170585_14590087,
        64'hf46300e4_5433942a,
        64'h47a500d4_14334405,
        64'h03b6869b_02f50533,
        64'h47a9c10d_44018d7d,
        64'hfff7c793_00e797b3,
        64'h57fdb7f5_7b450513,
        64'h00009517_85aafb07,
        64'h9de32785_5540406f,
        64'h61057ca5_05130000,
        64'h951785aa_690264a2,
        64'h60e26442_e495e04a,
        64'he822ec06_0007c483,
        64'he42697c2_11017f68,
        64'h08130000_a8179381,
        64'h1782cd85_00e555b3,
        64'h03c6871b_02f886bb,
        64'h481958d9_4781862e,
        64'hb78d7ea5_05130000,
        64'h951785aa_5ac0406f,
        64'h610581a5_05130000,
        64'ha5176902_64a285ca,
        64'h862660e2_64425c60,
        64'h40ef82a5_05130000,
        64'ha51785a2_c8015d60,
        64'h40ef84b2_83450513,
        64'h0000a517_f86102f4,
        64'h5433bfc1_02e45433,
        64'ha039943e_00144413,
        64'h03243413_02e47433,
        64'h02f457b3_06400713,
        64'h02877463_06300713,
        64'hc70502f4_773347a9,
        64'h0287e663_47293e80,
        64'h0793c021_02f555b3,
        64'h02f57433_bf7d2407,
        64'h87934685_b7d9a007,
        64'h87934681_63c0406f,
        64'h610588a5_05130000,
        64'ha51785aa_690264a2,
        64'h60e26442_02091663,
        64'he426e822_ec060007,
        64'h4903e04a_97361101,
        64'h8e870713_0000b717,
        64'h3e800793_46890ca7,
        64'hf7633e70_079304a7,
        64'h676323f7_8713000f,
        64'h47b704a7_6963862e,
        64'h9ff78713_3b9ad7b7,
        64'h8082612d_450160ee,
        64'h6a0040ef_8e450513,
        64'h0000a517_002cfebf,
        64'hf0efed86_45050c80,
        64'h0613002c_7115f73f,
        64'hf06f4581_862e86b2,
        64'h80826145_69a26942,
        64'h64e2854a_740270a2,
        64'h26e060ef_8fc58593,
        64'h0000a597_00890533,
        64'hffd4841b_00f44463,
        64'hffe4879b_9c296b60,
        64'h40ef954a_92c60613,
        64'h0000a617_86ce40a4,
        64'h85bb0095_5d630009,
        64'h8f63842a_6d4040ef,
        64'h854a85a6_94460613,
        64'h0000a617_dfc70713,
        64'h00009717_94c68693,
        64'h0000a697_c50919e6,
        64'h86930000_a6978932,
        64'h89ae84b6_f022f406,
        64'he44ee84a_ec267179,
        64'hbfdd7520_40ef8562,
        64'hb7e90905_75c040ef,
        64'h856600fb_e7630ff7,
        64'hf793fe05_879b0007,
        64'hc583012a_07b3b781,
        64'h04852405_77c040ef,
        64'h51850513_0000a517,
        64'h00f45b63_0009079b,
        64'hff047913_794040ef,
        64'h855aff2d_cce32d85,
        64'h7a0040ef_8556a029,
        64'h00f97913_4d81fffd,
        64'h4913028d_1d637b60,
        64'h40ef9d25_05130000,
        64'ha5170104_c583dbe5,
        64'hb7c57ca0_40ef8562,
        64'ha0317d20_40ef8556,
        64'h7d8040ef_57450513,
        64'h0000a517_ffb912e3,
        64'h09057ea0_40ef8566,
        64'h02fbe263_0ff7f793,
        64'hfe05879b_0007c583,
        64'h012487b3_4dc14901,
        64'h009040ef_855ae7a9,
        64'hc42900f4_77938082,
        64'h61656da2_6d426ce2,
        64'h7c027ba2_7b427ae2,
        64'h6a0669a6_694664e6,
        64'h740670a6_03344163,
        64'hfff58d1b_a44c8c93,
        64'h0000ac97_a54c0c13,
        64'h0000ac17_06000b93,
        64'ha48b0b13_0000ab17,
        64'h718a8a93_0000aa97,
        64'h4401ff05_049389ae,
        64'h8a2ae46e_e8caf486,
        64'he86aec66_f062f45e,
        64'hf85afc56_e0d2e4ce,
        64'heca6f0a2_7159b7cd,
        64'h089040ef_be07ae23,
        64'h0000b797_a7450513,
        64'h0000a517_80826151,
        64'h641260b2_85220a70,
        64'h40efa5a5_05130000,
        64'ha517a325_85930000,
        64'ha597860a_c10d842a,
        64'hdedff0ef_85220c70,
        64'h40efa525_05130000,
        64'ha517a525_85930000,
        64'ha597842a_00054603,
        64'h00154683_00254703,
        64'h00354783_00454803,
        64'h00554883_e222e606,
        64'h716d8082_7f010113,
        64'h7c813983_7d013903,
        64'h7d813483_7e013403,
        64'h45017e81_30836165,
        64'h8cfff0ef_86c685a6,
        64'h18085632_6882fbaf,
        64'hf0ef03e1_0513863e,
        64'h86c285a2_67c26822,
        64'hf8aff0ef_d64e0521,
        64'h051385a2_864a86ba,
        64'h943e7fc4_04136762,
        64'h747d97ba_81078793,
        64'h10186785_7ae060ef,
        64'hd602e83e_ec3ae442,
        64'h893689b2_e04605a1,
        64'h051384aa_71597d31,
        64'h34237d21_38237c91,
        64'h3c237e81_30237e11,
        64'h34238101_011318f0,
        64'h406fb025_05130000,
        64'ha51785aa_80826125,
        64'h7aa27a42_79e26906,
        64'h64a66446_450160e6,
        64'h911a6305_96bff0ef,
        64'h85ce86a6_10084652,
        64'h855ff0ef_460156fd,
        64'h02e10513_85a2821f,
        64'hf0ef0440_06130430,
        64'h06930421_051385a2,
        64'h943e1451_978a020a,
        64'h879312f1_1c233537,
        64'h87936799_12f11b23,
        64'h26378793_77e10510,
        64'h60ef04f1_06230661,
        64'h05134641_479985ce,
        64'h04f11523_10100793,
        64'h019060ef_ca3e04a1,
        64'h05134581_0f000613,
        64'h0fc00793_07f060ef,
        64'h000107a3_15410223,
        64'h14f101a3_14510513,
        64'h460585ca_57fd0990,
        64'h60ef13f1_05134611,
        64'h95beff04_0593978a,
        64'h020a8793_12f10f23,
        64'h479112f1_0ea30370,
        64'h07930bd0_60ef0141,
        64'h07a31a68_460585ca,
        64'h993e978a_020a8793,
        64'h12f11d23_13500793,
        64'hc83e4a05_fef40913,
        64'h439cd027_87930000,
        64'hb79709b0_60ef8526,
        64'h55fd4619_94beff84,
        64'h0493978a_020a8793,
        64'h747d2b30_40efca02,
        64'h6a85c125_05130000,
        64'ha517911a_89aaf456,
        64'hf852fc4e_e0cae4a6,
        64'he8a2ec86_711d737d,
        64'hb35d2db0_40efbfe5,
        64'h05130000_a517bf45,
        64'hbf850513_0000a517,
        64'h95be978a_d0040593,
        64'h35078793_67852ff0,
        64'h40efbf25_05130000,
        64'ha51730b0_40efbee5,
        64'h05130000_a51700fa,
        64'h20234785_de0796e3,
        64'h000a2783_bbcd3270,
        64'h40efbfa5_05130000,
        64'ha517b501_335040ef,
        64'hbf050513_0000a517,
        64'h95be978a_f0040593,
        64'h35048793_34d040ef,
        64'hbf850513_0000a517,
        64'h95bee004_0593978a,
        64'h35048793_365040ef,
        64'h02f5d5bb_e107879b,
        64'h678502f6_763b02f5,
        64'hf6bb02f5_d63b03c0,
        64'h0793f4f7_1e230000,
        64'hb7170121_5783f6f7,
        64'h13230000_b717c1e5,
        64'h05130000_a51755c2,
        64'h01015783_3a5040ef,
        64'hc1050513_0000a517,
        64'h01014583_01114603,
        64'h01214683_01314703,
        64'h3c1040ef_c0c50513,
        64'h0000a517_01814583,
        64'h01914603_01a14683,
        64'h01b14703_3dd040ef,
        64'h00b14703_fcf71323,
        64'h0000b717_c0c50513,
        64'h0000a517_00814583,
        64'h35215783_fcf71e23,
        64'h0000b717_00914603,
        64'h00a14683_35015783,
        64'h411040ef_c0c50513,
        64'h0000a517_35014583,
        64'h35114603_35214683,
        64'h35314703_27f060ef,
        64'h01490593_4611953e,
        64'hcb840513_978a3504,
        64'h87936485_297060ef,
        64'h0e880109_05934611,
        64'h451040ef_c3c50513,
        64'h0000a517_00fa2023,
        64'h47851207_9a63000a,
        64'h2783b311_d00d0023,
        64'h2c3060ef_9d228562,
        64'h866ab759_cc048513,
        64'hbb29cef4_2023401c,
        64'h00f40023_ce344783,
        64'h00f400a3_ce244783,
        64'h00f40123_ce144783,
        64'h00f401a3_ce044783,
        64'h2fb060ef_4611953e,
        64'hce048513_978a3507,
        64'h87936785_bfdd855a,
        64'h4611bbb1_317060ef,
        64'h85564611_b39df00d,
        64'h00233250_60ef9d22,
        64'h953e866a_f0048513,
        64'h978a3507_87936785,
        64'ha00d953e_978a3507,
        64'h87936785_4611cd04,
        64'h85138082_3b010113,
        64'h35013d03_35813c83,
        64'h36013c03_36813b83,
        64'h37013b03_37813a83,
        64'h38013a03_38813983,
        64'h39013903_39813483,
        64'h3a013403_3a813083,
        64'h911a6305_cebff0ef,
        64'h0e8885de_86ca5672,
        64'hbd5ff0ef_35e10513,
        64'h85a24601_56fdba1f,
        64'hf0ef3721_051385a2,
        64'h04400613_04300693,
        64'h943ecec4_0413978a,
        64'h350a8793_46f11423,
        64'h35378793_679946f1,
        64'h13232637_879377e1,
        64'h3d3060ef_36f10e23,
        64'h39610513_85de4799,
        64'h464136f1_1d231010,
        64'h079339b0_60efde3e,
        64'h37a10513_45810f00,
        64'h06131020_07934010,
        64'h60ef4731_0d230001,
        64'h03a346f1_0ca347b1,
        64'h051385a6_460557fd,
        64'h41b060ef_47410a23,
        64'h47510513_461195be,
        64'hcf440593_978a350a,
        64'h879346f1_09a30360,
        64'h079343d0_60ef4741,
        64'h072346f1_05134611,
        64'h4a1195be_cf040593,
        64'h978a350a_879346f1,
        64'h06a30320_07934610,
        64'h60efc0d2_46c10513,
        64'h85a64605_94becb74,
        64'h0493c2a6_978a350a,
        64'h879346f1_15231350,
        64'h079300f1_03a3478d,
        64'h439060ef_854a55fd,
        64'h4619993e_cf840913,
        64'h978a350a_879364f0,
        64'h40efde02_54e25a52,
        64'he2850513_0000a517,
        64'h4b3060ef_953e4611,
        64'h01490593_ce840513,
        64'h978a350a_87934c90,
        64'h60ef013c_a023953e,
        64'h46110109_0593ce44,
        64'h05134985_978a350a,
        64'h87936a85_16079263,
        64'h000ca783_3ae79d63,
        64'h470938e7_81634719,
        64'h24e78163_0007859b,
        64'h747d4715_00614783,
        64'hf8e79ce3_0ff00713,
        64'h24e78563_03800713,
        64'haad94605_cb648513,
        64'hfae798e3_03500713,
        64'h22e78063_03300713,
        64'h00f76e63_22e78363,
        64'h03600713_b759e00d,
        64'h00235450_60ef9d22,
        64'h953e866a_e0048513,
        64'h978a3507_87936785,
        64'hfee794e3_473d22e7,
        64'h85634731_b77d7170,
        64'h40ef0525_05130000,
        64'ha51785b6_22e78963,
        64'hcc848513_470d2ae7,
        64'h89634705_02f76263,
        64'h24e78163_471904f7,
        64'h6b6326e7_8d630007,
        64'h869b01a9_89bb0589,
        64'h02a00713_29890f07,
        64'hc7830015_cd030139,
        64'h07b395ca_0f098593,
        64'h9c3a9b3a_49818a36,
        64'h8cb28bae_d0048c13,
        64'hcb848b13_970a3507,
        64'h87139aba_cd848a93,
        64'h970a3507_871374fd,
        64'h678526f7_11634789,
        64'h00054703_a00179f0,
        64'h40eff525_05130000,
        64'ha51785aa_00e7ea63,
        64'h892a5800_073797aa,
        64'hd0040023_f0040023,
        64'he0040023_ca040b23,
        64'hce042023_d00007b7,
        64'h943e747d_978a911a,
        64'h35078793_35a13823,
        64'h35913c23_37813023,
        64'h37713423_37613823,
        64'h37513c23_39413023,
        64'h39313423_38913c23,
        64'h3a113423_39213823,
        64'h3a813023_6785737d,
        64'hc5010113_fadff06f,
        64'h614564e2_00e4859b,
        64'h70a27402_852200f4,
        64'h162347a1_67f060ef,
        64'h85b64619_852266a2,
        64'h68b060ef_e436f406,
        64'h46190519_84b2842a,
        64'hec26f022_71798082,
        64'h01416402_60a28522,
        64'hfa5ff0ef_e4064501,
        64'h85aa8622_0005841b,
        64'he0221141_bff105a1,
        64'h25050116_b02396ba,
        64'h010686bb_0035169b,
        64'h0005b883_808280c7,
        64'h3823973e_678500f5,
        64'h47636805_450102d7,
        64'hc7bb2785_0077e793,
        64'hfff6079b_8007bc23,
        64'h97ba46a1_67856398,
        64'h33878793_0000b797,
        64'h80826145_740270a2,
        64'h00f41523_fff7c793,
        64'h9fb94107_d71b9fb9,
        64'h93411742_4107579b,
        64'hfed79ce3_9f31ffe7,
        64'hd6030789_470187a2,
        64'h01440693_73f060ef,
        64'h01040513_002c4611,
        64'h74b060ef_00c40513,
        64'h00041523_006c4611,
        64'h00f404a3_47c57610,
        64'h60efec3e_00840513,
        64'h00041323_082c4621,
        64'h47c17750_60ef0044,
        64'h05130161_05934609,
        64'h783060ef_00f11b23,
        64'hc4360509_084c57fd,
        64'h460900f1_1a238fd9,
        64'h0087979b_0ff77713,
        64'h0087d713_c632842a,
        64'h419c00f5_10230457,
        64'h879b6785_c19c27d1,
        64'hf022f406_7179419c,
        64'h80820005_132300f5,
        64'h122300d5_112300c5,
        64'h10238fd9_0087979b,
        64'h0ff77713_c19c0087,
        64'hd7138ed9_06a20086,
        64'hd71b8e59_27a10622,
        64'h0086571b_419cc19c,
        64'h2785c319_0017f713,
        64'h419cbfcd_fda00513,
        64'h80826121_74a27442,
        64'h70e29782_85a66562,
        64'h701ce509_c39ff0ef,
        64'h842a0830_65a2c105,
        64'hc7dff0ef_84b2e42e,
        64'hf822fc06_f4267139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2655c,
        64'h862686ca_6562e519,
        64'hc75ff0ef_083065a2,
        64'hc115cb7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2615c,
        64'h862686ca_6562e519,
        64'hcb5ff0ef_083065a2,
        64'hc115cf7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hb7e16522_f569cdbf,
        64'hf0ef8526_85ce0030,
        64'hbfc90284_8493c501,
        64'h695060ef_854a608c,
        64'h288050ef_855285ca,
        64'h60908082_61216a42,
        64'h69e27902_74a27442,
        64'h70e24501_00849b63,
        64'h942602f4_043324ea,
        64'h0a130000_aa1789ae,
        64'h892afc06_e852ec4e,
        64'hf04a0280_079302f4,
        64'h043b840d_8c055a24,
        64'h84930000_b4975aa4,
        64'h04130000_b417f426,
        64'hf822639c_48478793,
        64'h0000b797_7139bfdd,
        64'h45018082_61056442,
        64'h60e2fda0_05138302,
        64'h610560e2_65a26442,
        64'h85220003_0e630205,
        64'h3303c919_db9ff0ef,
        64'he42eec06_4108842a,
        64'he8221101_bfc56562,
        64'hf96dd97f_f0ef0830,
        64'h80826145_70a24501,
        64'he50965a2_de1ff0ef,
        64'hf406e42e_7179bfc1,
        64'h5479fcf7_1be30ff0,
        64'h079300c7_c70367a2,
        64'h0e4080ef_6522f565,
        64'h842adcff_f0ef85a6,
        64'h00308522_80826145,
        64'h64e27402_70a28522,
        64'h54351100_80ef30e5,
        64'h05130000_a51700f4,
        64'hcf63445c_38c050ef,
        64'h31050513_0000a517,
        64'h85a6842a_c11dfda0,
        64'h0413e47f_f0ef84ae,
        64'hf406ec26_f0227179,
        64'h80826145_694264e2,
        64'h740270a2_852214a0,
        64'h80ef6522_3c4050ef,
        64'h33850513_0000a517,
        64'h864a608c_ed01842a,
        64'he45ff0ef_84aa85ca,
        64'h0030c11d_fda00413,
        64'he8dff0ef_892eec26,
        64'hf406e84a_f0227179,
        64'hb7d92405_188080ef,
        64'h65224020_50ef854e,
        64'h85a20127_896300c7,
        64'hc78367a2_ed09e83f,
        64'hf0ef8526_85a20030,
        64'h80826121_69e27902,
        64'h74a27442_70e200f4,
        64'h496344dc_39498993,
        64'h0000a997_0ff00913,
        64'h440184aa_cd01eebf,
        64'hf0efec4e_f04af426,
        64'hf822fc06_7139bfd5,
        64'h54798082_61457402,
        64'h70a28522_1ee080ef,
        64'h00f70963_00c54703,
        64'h0ff00793_6562e911,
        64'h842aee7f_f0ef0830,
        64'h65a2c105_fda00413,
        64'hf2dff0ef_e42ef406,
        64'hf0227179_b7c1fda0,
        64'h0513bf65_24052280,
        64'h80ef4981_65224a60,
        64'h50ef8552_00099563,
        64'h2485cb99_0087c783,
        64'h67a2ed19_f29ff0ef,
        64'h854a85a2_00308082,
        64'h61216a42_69e27902,
        64'h74a27442_70e24501,
        64'hc0915535_00f44d63,
        64'h00c92783_27ca0a13,
        64'h0000ba17_44014481,
        64'h4985892a_cd31f9bf,
        64'hf0efe852_ec4ef04a,
        64'hf426f822_fc067139,
        64'hbfe54501_80820141,
        64'h60a26108_c509fbbf,
        64'hf0efe406_1141b7f5,
        64'h02870713_fea68de3,
        64'h47148082_853a4701,
        64'h00e79563_97ba02d7,
        64'h87b30280_069302d7,
        64'h87bb878d_8f9981a7,
        64'h87930000_c7976294,
        64'h82470713_0000c717,
        64'h6f868693_0000b697,
        64'hb7edfda0_07138302,
        64'h853e85b2_00030563,
        64'h01853303_8082853a,
        64'he21c97b6_470102a7,
        64'h87b30a00_051300b7,
        64'hd963454c_0005cc63,
        64'h5735c285_87ae6914,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h000a2e2e_2e746e65,
        64'h6d6f6d20_61207469,
        64'h61772065_7361656c,
        64'h50202165_6e616972,
        64'h41206d6f_7266206f,
        64'h6c6c6548_ffdff06f,
        64'h10500073_34102373,
        64'h342022f3_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_69a090ef,
        64'hfec5c6e3_02058593,
        64'h0005bc23_0005b823,
        64'h0005b423_0005b023,
        64'h1c860613_0000c617,
        64'ha3058593_0000c597,
        64'h30579073_09078793,
        64'h00000797_00078067,
        64'h40b787b3_00d787b3,
        64'h01478793_00000797,
        64'hfcc5cce3_02068693,
        64'h02058593_00e6bc23,
        64'h0185b703_00e6b823,
        64'h0105b703_00e6b423,
        64'h0085b703_00e6b023,
        64'h0005b703_0006b703,
        64'hff810113_01b11113,
        64'h0110011b_fe0e9ae3,
        64'h0085b703_fffe8e93,
        64'h0005b703_240e8e9b,
        64'h000f4eb7_01169693,
        64'h3ff6869b_000046b7,
        64'ha1c60613_0000c617,
        64'hfc058593_00000597,
        64'h000280e7_13050513,
        64'h00000517_0b828293,
        64'h00008297_000280e7,
        64'h09228293_00008297,
        64'h01111113_3ff1011b,
        64'h00004137_11249463,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
