/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'h01111113fff1011b0000613711249463, /*    1 */
128'h00008297000280e70542829300008297, /*    2 */
128'h000280e7130505130000051707a28293, /*    3 */
128'h81c606130000c617fc05859300000597, /*    4 */
128'h000f4eb701169693fff6869b000066b7, /*    5 */
128'h0085b703fffe8e930005b703240e8e9b, /*    6 */
128'hff81011301b111130110011bfe0e9ae3, /*    7 */
128'h0085b70300e6b0230005b7030006b703, /*    8 */
128'h0185b70300e6b8230105b70300e6b423, /*    9 */
128'hfcc5cce3020686930205859300e6bc23, /*   10 */
128'h40b787b300d787b30147879300000797, /*   11 */
128'h30579073090787930000079700078067, /*   12 */
128'hd90606130000c617830585930000c597, /*   13 */
128'h0005bc230005b8230005b4230005b023, /*   14 */
128'h020004b745e090effec5c6e302058593, /*   15 */
128'h02000937004484930124a02300100913, /*   16 */
128'h3440297310500073ff24c6e34009091b, /*   17 */
128'hf1402973020004b7fe090ae300897913, /*   18 */
128'h0004a903000920230099093300291913, /*   19 */
128'h4009091b0200093700448493fe091ee3, /*   20 */
128'h1050007334102373342022f3ff24c6e3, /*   21 */
128'h41206d6f7266206f6c6c6548ffdff06f, /*   22 */
128'h617720657361656c502021656e616972, /*   23 */
128'h000a2e2e2e746e656d6f6d2061207469, /*   24 */
128'h00000000000000000000000000000000, /*   25 */
128'h00000000000000000000000000000000, /*   26 */
128'h00000000000000000000000000000000, /*   27 */
128'h00000000000000000000000000000000, /*   28 */
128'h00000000000000000000000000000000, /*   29 */
128'h00000000000000000000000000000000, /*   30 */
128'h00000000000000000000000000000000, /*   31 */
128'hd963454c0005cc635735c28587ae6914, /*   32 */
128'he21c97b6470102a787b30a00051300b7, /*   33 */
128'h853e85b200030563018533038082853a, /*   34 */
128'h4d8686930000b697b7edfda007138302, /*   35 */
128'h87930000b7976294624707130000b717, /*   36 */
128'h87b30280069302d787bb878d8f9961a7, /*   37 */
128'h47148082853a470100e7956397ba02d7, /*   38 */
128'hf0efe4061141b7f502870713fea68de3, /*   39 */
128'hbfe545018082014160a26108c509fbbf, /*   40 */
128'hf0efe852ec4ef04af426f822fc067139, /*   41 */
128'h0000ba17440144814985892acd31f9bf, /*   42 */
128'hc091553500f44d6300c9278300ca0a13, /*   43 */
128'h61216a4269e2790274a2744270e24501, /*   44 */
128'h67a2ed19f29ff0ef854a85a200308082, /*   45 */
128'h50ef8552000995632485cb990087c783, /*   46 */
128'h0513bf652405178080ef4981652249a0, /*   47 */
128'hf2dff0efe42ef406f0227179b7c1fda0, /*   48 */
128'h842aee7ff0ef083065a2c105fda00413, /*   49 */
128'h00f7096300c547030ff007936562e911, /*   50 */
128'h547980826145740270a2852213e080ef, /*   51 */
128'hf0efec4ef04af426f822fc067139bfd5, /*   52 */
128'h0000a9970ff00913440184aacd01eebf, /*   53 */
128'h74a2744270e200f4496344dc17498993, /*   54 */
128'hf0ef852685a200308082612169e27902, /*   55 */
128'h85a20127896300c7c78367a2ed09e83f, /*   56 */
128'hb7d924050d8080ef65223f6050ef854e, /*   57 */
128'he8dff0ef892eec26f406e84af0227179, /*   58 */
128'he45ff0ef84aa85ca0030c11dfda00413, /*   59 */
128'h118505130000a517864a608ced01842a, /*   60 */
128'h740270a2852209a080ef65223b8050ef, /*   61 */
128'hf406ec26f022717980826145694264e2, /*   62 */
128'h85a6842ac11dfda00413e47ff0ef84ae, /*   63 */
128'hcf63445c380050ef0f0505130000a517, /*   64 */
128'h5435060080ef0ee505130000a51700f4, /*   65 */
128'h003085228082614564e2740270a28522, /*   66 */
128'h034080ef6522f565842adcfff0ef85a6, /*   67 */
128'h5479fcf71be30ff0079300c7c70367a2, /*   68 */
128'he50965a2de1ff0eff406e42e7179bfc1, /*   69 */
128'hf96dd97ff0ef08308082614570a24501, /*   70 */
128'he42eec064108842ae8221101bfc56562, /*   71 */
128'h852200030e6302053303c919db9ff0ef, /*   72 */
128'h60e2fda005138302610560e265a26442, /*   73 */
128'h0000b7977139bfdd4501808261056442, /*   74 */
128'h04130000b417f426f822639c26478793, /*   75 */
128'h043b840d8c053a2484930000b4973aa4, /*   76 */
128'h892afc06e852ec4ef04a0280079302f4, /*   77 */
128'h942602f4043302ea0a130000aa1789ae, /*   78 */
128'h69e2790274a2744270e2450100849b63, /*   79 */
128'h27c050ef855285ca6090808261216a42, /*   80 */
128'hbfc902848493c501689060ef854a608c, /*   81 */
128'hb7e16522f569cdbff0ef852685ce0030, /*   82 */
128'h84b68432e42efc06f04af426f8227139, /*   83 */
128'hcb5ff0ef083065a2c115cf7ff0ef893a, /*   84 */
128'h70e2978285a2615c862686ca6562e519, /*   85 */
128'hbfc5fda0051380826121790274a27442, /*   86 */
128'h84b68432e42efc06f04af426f8227139, /*   87 */
128'hc75ff0ef083065a2c115cb7ff0ef893a, /*   88 */
128'h70e2978285a2655c862686ca6562e519, /*   89 */
128'hbfc5fda0051380826121790274a27442, /*   90 */
128'hc7dff0ef84b2e42ef822fc06f4267139, /*   91 */
128'h701ce509c39ff0ef842a083065a2c105, /*   92 */
128'h8082612174a2744270e2978285a66562, /*   93 */
128'h2785c3190017f713419cbfcdfda00513, /*   94 */
128'hd71b8e5927a106220086571b419cc19c, /*   95 */
128'h0ff77713c19c0087d7138ed906a20086, /*   96 */
128'h122300d5112300c510238fd90087979b, /*   97 */
128'hf022f4067179419c80820005132300f5, /*   98 */
128'h419c00f510230457879b6785c19c27d1, /*   99 */
128'h0087979b0ff777130087d713c632842a, /*  100 */
128'hc4360509084c57fd460900f11a238fd9, /*  101 */
128'h0513016105934609777060ef00f11b23, /*  102 */
128'h00041323082c462147c1769060ef0044, /*  103 */
128'h00f404a347c5755060efec3e00840513, /*  104 */
128'h73f060ef00c4051300041523006c4611, /*  105 */
128'h01440693733060ef01040513002c4611, /*  106 */
128'hfed79ce39f31ffe7d6030789470187a2, /*  107 */
128'h9fb94107d71b9fb9934117424107579b, /*  108 */
128'h80826145740270a200f41523fff7c793, /*  109 */
128'h97ba46a167856398138787930000b797, /*  110 */
128'hc7bb27850077e793fff6079b8007bc23, /*  111 */
128'h3823973e678500f547636805450102d7, /*  112 */
128'h010686bb0035169b0005b883808280c7, /*  113 */
128'he0221141bff105a125050116b02396ba, /*  114 */
128'hfa5ff0efe406450185aa86220005841b, /*  115 */
128'hec26f022717980820141640260a28522, /*  116 */
128'h67f060efe436f4064619051984b2842a, /*  117 */
128'h162347a1673060ef85b64619852266a2, /*  118 */
128'h614564e200e4859b70a27402852200f4, /*  119 */
128'h3a8130236785737dc5010113fadff06f, /*  120 */
128'h3931342338913c233a11342339213823, /*  121 */
128'h377134233761382337513c2339413023, /*  122 */
128'h3507879335a1382335913c2337813023, /*  123 */
128'hce042023d00007b7943e747d978a911a, /*  124 */
128'hd0040023f0040023e0040023ca040b23, /*  125 */
128'ha51785aa00e7ea63892a5800073797aa, /*  126 */
128'h00054703a001793040efd32505130000, /*  127 */
128'h970a3507871374fd678526f711634789, /*  128 */
128'hcb848b13970a350787139abacd848a93, /*  129 */
128'h9c3a9b3a49818a368cb28baed0048c13, /*  130 */
128'hc7830015cd03013907b395ca0f098593, /*  131 */
128'h869b01a989bb058902a0071329890f07, /*  132 */
128'h24e78163471904f76b6326e78d630007, /*  133 */
128'hcc848513470d2ae78963470502f76263, /*  134 */
128'h40efe22505130000a51785b622e78963, /*  135 */
128'hfee794e3473d22e785634731b77d70b0, /*  136 */
128'h953e866ae0048513978a350787936785, /*  137 */
128'h03600713b759e00d0023539060ef9d22, /*  138 */
128'h22e780630330071300f76e6322e78363, /*  139 */
128'haad94605cb648513fae798e303500713, /*  140 */
128'hf8e79ce30ff0071324e7856303800713, /*  141 */
128'h24e781630007859b747d471500614783, /*  142 */
128'h000ca7833ae79063470936e784634719, /*  143 */
128'h05134985978a350a87936a8516079263, /*  144 */
128'h60ef013ca023953e461101090593ce44, /*  145 */
128'h01490593ce840513978a350a87934bd0, /*  146 */
128'hc08505130000a5174a7060ef953e4611, /*  147 */
128'h978a350a8793643040efde0254e25a52, /*  148 */
128'h42d060ef854a55fd4619993ecf840913, /*  149 */
128'h879346f115231350079300f103a3478d, /*  150 */
128'h85a6460594becb740493c2a6978a350a, /*  151 */
128'h06a303200793455060efc0d246c10513, /*  152 */
128'h4a1195becf040593978a350a879346f1, /*  153 */
128'h0793431060ef4741072346f105134611, /*  154 */
128'hcf440593978a350a879346f109a30360, /*  155 */
128'h40f060ef47410a2347510513461195be, /*  156 */
128'h03a346f10ca347b1051385a6460557fd, /*  157 */
128'h0613102007933f5060ef47310d230001, /*  158 */
128'h079338f060efde3e37a1051345810f00, /*  159 */
128'h3961051385de4799464136f11d231010, /*  160 */
128'h13232637879377e13c7060ef36f10e23, /*  161 */
128'h350a879346f1142335378793679946f1, /*  162 */
128'h0440061304300693943ecec40413978a, /*  163 */
128'h85a2460156fdba1ff0ef3721051385a2, /*  164 */
128'h0e8885de86ca5672bd5ff0ef35e10513, /*  165 */
128'h3a0134033a813083911a6305cebff0ef, /*  166 */
128'h38013a03388139833901390339813483, /*  167 */
128'h36013c0336813b8337013b0337813a83, /*  168 */
128'h851380823b01011335013d0335813c83, /*  169 */
128'ha00d953e978a3507879367854611cd04, /*  170 */
128'h953e866af0048513978a350787936785, /*  171 */
128'h85564611b39df00d0023319060ef9d22, /*  172 */
128'h87936785bfdd855a4611bbb130b060ef, /*  173 */
128'h2ef060ef4611953ece048513978a3507, /*  174 */
128'h00f40123ce14478300f401a3ce044783, /*  175 */
128'h00f40023ce34478300f400a3ce244783, /*  176 */
128'h866ab759cc048513bb29cef42023401c, /*  177 */
128'h2783b311d00d00232b7060ef9d228562, /*  178 */
128'h0000a51700fa2023478510079d63000a, /*  179 */
128'h0e88010905934611445040efa1c50513, /*  180 */
128'hcb840513978a35048793648528b060ef, /*  181 */
128'h35314703273060ef014905934611953e, /*  182 */
128'h0000a517350145833511460335214683, /*  183 */
128'h00a1468335015783405040ef9ec50513, /*  184 */
128'h35215783dcf71e230000b71700914603, /*  185 */
128'h0000b7179ec505130000a51700814583, /*  186 */
128'h01b147033d1040ef00b14703dcf71323, /*  187 */
128'h0000a517018145830191460301a14683, /*  188 */
128'h01214683013147033b5040ef9ec50513, /*  189 */
128'h9f0505130000a5170101458301114603, /*  190 */
128'h05130000a51755c201015783399040ef, /*  191 */
128'hb71701215783d6f713230000b7179fe5, /*  192 */
128'h978a35048793373040efd4f71e230000, /*  193 */
128'h40ef9ea505130000a51795bee0040593, /*  194 */
128'ha51795be978af00405933504879335b0, /*  195 */
128'h0000a517bd29343040ef9e2505130000, /*  196 */
128'h93e3000a2783b531335040ef9e450513, /*  197 */
128'h9d8505130000a51700fa20234785e007, /*  198 */
128'h30d040ef9dc505130000a517319040ef, /*  199 */
128'ha51795be978ad0040593350787936785, /*  200 */
128'h9e8505130000a517bf459e2505130000, /*  201 */
128'he4a6e8a2ec86711d737db3c12e9040ef, /*  202 */
128'h0000a517911a89aaf456f852fc4ee0ca, /*  203 */
128'h8793747d2c1040efca026a859fc50513, /*  204 */
128'h852655fd461994beff840493978a020a, /*  205 */
128'h0913439cb1c787930000b7970a9060ef, /*  206 */
128'h879312f11d2313500793c83e4a05fef4, /*  207 */
128'h014107a31a68460585ca993e978a020a, /*  208 */
128'h0f23479112f10ea3037007930cb060ef, /*  209 */
128'h461195beff040593978a020a879312f1, /*  210 */
128'h0513460585ca57fd0a7060ef13f10513, /*  211 */
128'h60ef000107a31541022314f101a31451, /*  212 */
128'h04a1051345810f0006130fc0079308d0, /*  213 */
128'h85ce04f1152310100793027060efca3e, /*  214 */
128'h05f060ef04f106230661051346414799, /*  215 */
128'h35378793679912f11b232637879377e1, /*  216 */
128'h85a2943e1451978a020a879312f11c23, /*  217 */
128'h83bff0ef044006130430069304210513, /*  218 */
128'h465286fff0ef460156fd02e1051385a2, /*  219 */
128'h60e6911a6305985ff0ef85ce86a61008, /*  220 */
128'h61257aa27a4279e2690664a664464501, /*  221 */
128'h19d0406f8ec505130000a51785aa8082, /*  222 */
128'h7c913c237e8130237e11342381010113, /*  223 */
128'h05a1051384aa71597d3134237d213823, /*  224 */
128'h60efd602e83eec3ae442893689b2e046, /*  225 */
128'h6762747d97ba81078793101867857bc0, /*  226 */
128'h0521051385a2864a86ba943e7fc40413, /*  227 */
128'h863e86c285a267c26822fa4ff0efd64e, /*  228 */
128'h85a6180856326882fd4ff0ef03e10513, /*  229 */
128'h340345017e81308361658e9ff0ef86c6, /*  230 */
128'h01137c8139837d0139037d8134837e01, /*  231 */
128'h480300554883e222e606716d80827f01, /*  232 */
128'h46030015468300254703003547830045, /*  233 */
128'h0000a51783c585930000a597842a0005, /*  234 */
128'h842adedff0ef85220d5040ef83c50513, /*  235 */
128'h0000a51781c585930000a597860ac10d, /*  236 */
128'h6151641260b285220b5040ef84450513, /*  237 */
128'hab230000b79785e505130000a5178082, /*  238 */
128'he4ceeca6f0a27159b7cd097040efa007, /*  239 */
128'hf486e86aec66f062f45ef85afc56e0d2, /*  240 */
128'haa974401ff05049389ae8a2ae46ee8ca, /*  241 */
128'h0b93832b0b130000ab1754aa8a930000, /*  242 */
128'h8c930000ac9783ec0c130000ac170600, /*  243 */
128'h64e6740670a603344163fff58d1b82ec, /*  244 */
128'h6ce27c027ba27b427ae26a0669a66946, /*  245 */
128'he7a9c42900f47793808261656da26d42, /*  246 */
128'hc583012487b34dc14901017040ef855a, /*  247 */
128'h856602fbe2630ff7f793fe05879b0007, /*  248 */
128'h05130000a517ffb912e309057f8040ef, /*  249 */
128'h8562a0317e0040ef85567e6040ef31e5, /*  250 */
128'h000095170104c583dbe5b7c57d8040ef, /*  251 */
128'hfffd4913028d1d637c4040ef7bc50513, /*  252 */
128'h2d857ae040ef8556a02900f979134d81, /*  253 */
128'h079bff0479137a2040ef855aff2dcce3, /*  254 */
128'h40ef2c2505130000a51700f45b630009, /*  255 */
128'h0007c583012a07b3b7810485240578a0, /*  256 */
128'h40ef856600fbe7630ff7f793fe05879b, /*  257 */
128'h7179bfdd760040ef8562b7e9090576a0, /*  258 */
128'h893289ae84b6f022f406e44ee84aec26, /*  259 */
128'h869300009697c509fd8686930000a697, /*  260 */
128'h061300009617c1670713000097177366, /*  261 */
128'h00098f63842a6e2040ef854a85a672e6, /*  262 */
128'h06130000961786ce40a485bb00955d63, /*  263 */
128'h4463ffe4879b9c296c4040ef954a7166, /*  264 */
128'h85930000959700890533ffd4841b00f4, /*  265 */
128'h694264e2854a740270a227c060ef6e65, /*  266 */
128'hf73ff06f4581862e86b28082614569a2, /*  267 */
128'hfebff0efed8645050c800613002c7115, /*  268 */
128'h60ee6ae040ef6ce5051300009517002c, /*  269 */
128'h862e9ff787133b9ad7b78082612d4501, /*  270 */
128'h04a7676323f78713000f47b704a76963, /*  271 */
128'ha7173e80079346890ca7f7633e700793, /*  272 */
128'h00074903e04a97361101702707130000, /*  273 */
128'h64a260e2644202091663e426e822ec06, /*  274 */
128'h406f6105674505130000951785aa6902, /*  275 */
128'h240787934685b7d9a0078793468164a0, /*  276 */
128'h3e800793c02102f555b302f57433bf7d, /*  277 */
128'h0713c70502f4773347a90287e6634729, /*  278 */
128'h743302f457b306400713028774630630, /*  279 */
128'h5433a039943e001444130324341302e4, /*  280 */
128'h051300009517f86102f45433bfc102e4, /*  281 */
128'h0000951785a2c8015e4040ef84b261e5, /*  282 */
128'h85ca862660e264425d4040ef61450513, /*  283 */
128'h406f61056045051300009517690264a2, /*  284 */
128'h862eb78d5d4505130000951785aa5ba0, /*  285 */
128'h55b303c6871b02f886bb481958d94781, /*  286 */
128'h610808130000a81793811782cd8500e5, /*  287 */
128'he04ae822ec060007c483e42697c21101, /*  288 */
128'h0000951785aa690264a260e26442e495, /*  289 */
128'hfb079de327855620406f61055b450513, /*  290 */
128'h97b357fdb7f559e505130000951785aa, /*  291 */
128'h053347a9c10d44018d7dfff7c79300e7, /*  292 */
128'h942a47a500d41433440503b6869b02f5, /*  293 */
128'h00009517058514590087f46300e45433, /*  294 */
128'h951785a2c801512040ef893254c50513, /*  295 */
128'h864a60e26442502040ef542505130000, /*  296 */
128'h610554a505130000951764a2690285a6, /*  297 */
128'hf1a202c7073b8cbaed6671514e80406f, /*  298 */
128'hf95afd56e1d2eda6f586e96ae5cee9ca, /*  299 */
128'h8d3289ae892a04000793e56ef162f55e, /*  300 */
128'h956302ccdcbb04000c9300e7f6638436, /*  301 */
128'h020d1a13001d179b03acdcbb4cc1000c, /*  302 */
128'h9b1703810a93020a5a130017849be03e, /*  303 */
128'h8c1745ab8b9300009b974f2b0b130000, /*  304 */
128'h64ee740e70ae4501e00d3f2c0c130000, /*  305 */
128'h6cea7c0a7baa7b4a7aea6a0e69ae694e, /*  306 */
128'h05130000951785ca8082616d6daa6d4a, /*  307 */
128'h8d9b008cf46300040d9b446040ef4ae5, /*  308 */
128'h0007061b430948a14811470186ce000c, /*  309 */
128'h99ba034707339301020d971305b66c63, /*  310 */
128'h861b02e00813875603bd06bb0d9de663, /*  311 */
128'h85d6963e011c0ac5ed63415705bb0006, /*  312 */
128'h40effa060c23e4364685051300009517, /*  313 */
128'h70ef99369281168241b4043b66a23ea0, /*  314 */
128'h15934290030d1b63b795557dd1350220, /*  315 */
128'h855a658292011602c190260195d60027, /*  316 */
128'h66a23ae040efe436e83aec42f046f41a, /*  317 */
128'h1863bf8568627882070596d273226742, /*  318 */
128'h1c63bfc1e19095d6003715936290011d, /*  319 */
128'h9241164295d6001715930006d603006d, /*  320 */
128'h761300ea85b30006c603bf6500c59023, /*  321 */
128'h04e070efe43a855eb75d00c580230ff6, /*  322 */
128'hbfdd4701bf1d3cfdfe976ae327056722, /*  323 */
128'h097575130005450300bc053300074583, /*  324 */
128'h00230005d4634185d59b0185959bc519, /*  325 */
128'hf4634501918187aa1582bf3907050107, /*  326 */
128'h04000793bfd58f8d25058082e21c00b7, /*  327 */
128'h57f70713464c47370005668312b7f463, /*  328 */
128'h10e6976347090045468310e69c634789, /*  329 */
128'hf0a202f7073371590380079303855703, /*  330 */
128'he4cee8caeca6f48602059a93fc567100, /*  331 */
128'hda93e46ee86aec66f062f45ef85ae0d2, /*  332 */
128'h942a84aa892e06eae663478d9722020a, /*  333 */
128'h00009c1731cb8b9300009b974b054a01, /*  334 */
128'h0384d78333cc8c9300009c9735cc0c13, /*  335 */
128'h741c09679b63401ca835478100fa6463, /*  336 */
128'h8d6302043983272040ef855e85d2cbc1, /*  337 */
128'hfa6395ce00b48db301843d03640c0409, /*  338 */
128'h24c040ef2dc5051300009517864a02ba, /*  339 */
128'h7ae26a0669a6694664e6740670a6478d, /*  340 */
128'h6165853e6da26d426ce27c027ba27b42, /*  341 */
128'h864e21e040ef856686ce85ea866e8082, /*  342 */
128'hf163701c02843983066060ef856a85ee, /*  343 */
128'h85ea9d3e864e40f989b301843d030337, /*  344 */
128'h7ed050ef856a4581864e1f6040ef8562, /*  345 */
128'h45058082853e4785bf99038404132a05, /*  346 */
128'h07130000a7178082400005378082057e, /*  347 */
128'h95360017869300756513157d631c36e7, /*  348 */
128'h8082953e057e450597aa20000537e308, /*  349 */
128'h08a74463862a0ce50763820787136785, /*  350 */
128'h06e60b6327c505130000951780878713, /*  351 */
128'h25850513000095178006079b04c74963, /*  352 */
128'h2d8505130000951787f787936785c3ad, /*  353 */
128'h95979e3d11417c07879b77fd04c7c963, /*  354 */
128'he4062d2505130000a5172ca585930000, /*  355 */
128'h01412c2505130000a51760a2124040ef, /*  356 */
128'h0a6322a5051300009517810787138082, /*  357 */
128'h12e322a50513000095178187879300e6, /*  358 */
128'h2485051300009517830787138082faf6, /*  359 */
128'h000095178287879300c74963fee609e3, /*  360 */
128'h05130000951783878713bfe922450513, /*  361 */
128'h05130000951784078793fce608e32365, /*  362 */
128'h717980821ec5051300009517bf752365, /*  363 */
128'h4463440184ae892af406e84aec26f022, /*  364 */
128'h01045513942a90411442010455130290, /*  365 */
128'h694264e21542fff54513740270a29522, /*  366 */
128'h6df050ef0068460985ca808261459141, /*  367 */
128'h00d1478300f107a334f9090900c14783, /*  368 */
128'h6785715dbf55943e00e1578300f10723, /*  369 */
128'h842e80678793f44ef84afc26e486e0a2, /*  370 */
128'h079b0af50e636dd7879367a13cf50563, /*  371 */
128'h50ef4611082884b205e944079a638005, /*  372 */
128'h05130000a517461985ca0064091368d0, /*  373 */
128'h896302e0079301744583679050ef1c65, /*  374 */
128'h04b7e5631cf5826347b108b7e76332f5, /*  375 */
128'h10f58463478502b7e3631af583634791, /*  376 */
128'h951702f5836317650513000095174789, /*  377 */
128'h82634799a41d7e3030ef312505130000, /*  378 */
128'hfef591e317c505130000951747a118f5, /*  379 */
128'h00b7ed632cf5826347f5a4317c9030ef, /*  380 */
128'h198505130000951747d916f58a6347c5, /*  381 */
128'h07932af5866302100793bf6dfef580e3, /*  382 */
128'hb7c91b25051300009517faf596e30290, /*  383 */
128'h0330079304b7e2632cf5826306200793, /*  384 */
128'h28f5876302f0079300b7ef632af58263, /*  385 */
128'hf8f58ae31b4505130000951703200793, /*  386 */
128'h951705e0079328f5846305c00793b7bd, /*  387 */
128'h08400793bf91f6f58de31ca505130000, /*  388 */
128'h26f58b630670079300b7ef6328f58663, /*  389 */
128'hf4f58ae31dc505130000951706c00793, /*  390 */
128'h89630ff0079326f5886308900793b73d, /*  391 */
128'h051300009517f0f59ce30880079326f5, /*  392 */
128'h0d87d7830000a79701e45703b73d1e65, /*  393 */
128'h0204570312f714630d0989930000a997, /*  394 */
128'h85ca461910f71c630c27d7830000a797, /*  395 */
128'h090585930000a5974619519050ef8522, /*  396 */
128'h12230204012301a45783509050ef854a, /*  397 */
128'h0513fde4859b01c4578300f41f230204, /*  398 */
128'hd78300f41d230009d78302f410230224, /*  399 */
128'h812100a10ea3db9ff0ef00f41e230029, /*  400 */
128'h85a202f41223862601c1578300a10e23, /*  401 */
128'hfe85051300009517a06ddbffe0ef4501, /*  402 */
128'h00009517b559ff65051300009517bd41, /*  403 */
128'h0ea30264470302444783bdb500450513, /*  404 */
128'h0ea301c1178300f10e230254478300f1, /*  405 */
128'h0224470300e10e2327810274470300e1, /*  406 */
128'h00e10e230234470300e10ea301c11903, /*  407 */
128'h0000a79704e79b6301c1568304500713, /*  408 */
128'hf88585930000a597461947e2fad79823, /*  409 */
128'hf8f728230000a717f90505130000a517, /*  410 */
128'h87930000a79766a24762429050efe436, /*  411 */
128'h508060ef450102a40593ff89061bf667, /*  412 */
128'h07138082616179a2794274e2640660a6, /*  413 */
128'hf4f728230000a71747e204e694630430, /*  414 */
128'h0000a797c799439cf54787930000a797, /*  415 */
128'hf38686930000a697f7e9439cf4478793, /*  416 */
128'hf38585930000a597f34606130000a617, /*  417 */
128'h98634d200713b765d61fe0ef02a40513, /*  418 */
128'h85a654f030eff1e505130000951702e7, /*  419 */
128'h30eff1a5051300009517cb6ff0ef8522, /*  420 */
128'h0713bf95ca0ff0ef02a4051385ca53b0, /*  421 */
128'h01e317fd67c101e45703f6e787e35fe0, /*  422 */
128'h0000a5974611f4f70de302045703f6f7, /*  423 */
128'h00009517b799355050ef0868ef458593, /*  424 */
128'hb30defa5051300009517b335ef450513, /*  425 */
128'h051300009517bb21f105051300009517, /*  426 */
128'h9517b311f345051300009517b339f1e5, /*  427 */
128'hf585051300009517b9edf3a505130000, /*  428 */
128'h00009517b1ddf665051300009517b9c5, /*  429 */
128'hb9c9fa25051300009517b9f1f7c50513, /*  430 */
128'ha7970265d703b1e1fb05051300009517, /*  431 */
128'h11e3e6a484930000a497e727d7830000, /*  432 */
128'h19e3e5c7d7830000a7970285d703ecf7, /*  433 */
128'h9a23016589930205891320000793eaf7, /*  434 */
128'ha59746192a3050ef854a85ce461900f5, /*  435 */
128'ha5974619293050ef854ee1a585930000, /*  436 */
128'h4619281050ef00640513e0a585930000, /*  437 */
128'h02a0061301c45783277050ef852285ca, /*  438 */
128'h0004d78302f4142301e4578302f41323, /*  439 */
128'h6080079300f41f230024d78300f41e23, /*  440 */
128'hf38505130000951785aab36900f41623, /*  441 */
128'h8307b603300017b7bba546013e9030ef, /*  442 */
128'h171b00f674132601608130239f010113, /*  443 */
128'h05379f2d8406871b0387759366850034, /*  444 */
128'h34235e913c23630c8387b783972a3000, /*  445 */
128'h696335b95f200813ffc5849b25816011, /*  446 */
128'hfff7c79300c5963b101005938a1d08b8, /*  447 */
128'h4390d42787930000a797cfb527818ff1, /*  448 */
128'h9ebd8006869b7007f7930084179bea25, /*  449 */
128'h0106969b00d100a3872646d496aa068e, /*  450 */
128'h0001550300d100230086d69b0106d69b, /*  451 */
128'h02d51a63806686936685c6918005069b, /*  452 */
128'h46a1007767139fad377d8005859b6585, /*  453 */
128'h08378f95868a83f502d7473b17822705, /*  454 */
128'haa1ff0ef862602e6446397c285b63000, /*  455 */
128'h3403608130838287b823300017b70405, /*  456 */
128'h88338082610101135f81348385266001, /*  457 */
128'hb7e1ff06bc2306a126050008380300d7, /*  458 */
128'h2401ec06e42643c0e8220c2007b71101, /*  459 */
128'hc163033716938304b703300014b74781, /*  460 */
128'h2ad030efe145051300009517e7990206, /*  461 */
128'h8082610564a2644260e2c3c00c2007b7, /*  462 */
128'h8432ec26f0227179bfc14785eb9ff0ef, /*  463 */
128'hf4060068c6c585930000a597461184ae, /*  464 */
128'h0007a803c24787930000a7970cb050ef, /*  465 */
128'ha717c0a888930000a89785a6862247b2, /*  466 */
128'h05130000a51704500693c0e757030000, /*  467 */
128'h614564e2740270a285228aeff0efc165, /*  468 */
128'h8082914115428d5d05220085579b8082, /*  469 */
128'hf00686938fd966c10185579b0185171b, /*  470 */
128'h00ff07370085151b8fd98f750085571b, /*  471 */
128'h051300009517715d808225018d5d8d79, /*  472 */
128'hec56f052f44ef84afc26e0a2e486d765, /*  473 */
128'h47e1ba0785230000a7971e7030efe85a, /*  474 */
128'h0000a71703e00793baf700a30000a717, /*  475 */
128'h578db8f706a30000a7174789b8f70b23, /*  476 */
128'ha59707f007934611b8f702230000a717, /*  477 */
128'hb68404130000a4170028b74585930000, /*  478 */
128'h85a246097e2050efb6f702a30000a717, /*  479 */
128'h89930000a997448145227d8050ef0068, /*  480 */
128'hf00606130100063746b2f4fff0efb2e9, /*  481 */
128'h15028f558f710ff6f69382a10086971b, /*  482 */
128'hb423934180a7b02317429101300017b7, /*  483 */
128'h0513000095178087b7038007b70380e7, /*  484 */
128'h8087b5838007b60382e7b4234721cc65, /*  485 */
128'h91c115c2adca0a130000aa1700800737, /*  486 */
128'h47030000a717113030ef80e7b4238f4d, /*  487 */
128'h48030000a817ad27c7830000a797ad97, /*  488 */
128'h46030000a617ac06c6830000a697acb8, /*  489 */
128'h051300009517aae5c5830000a597ab76, /*  490 */
128'h00989b376a89000447830d7030efc765, /*  491 */
128'h3000193700144783a8f70c230000a717, /*  492 */
128'h0000a71700244783a8f704a30000a717, /*  493 */
128'ha6f709a30000a71700344783a6f70f23, /*  494 */
128'h00544783a6f704230000a71700444783, /*  495 */
128'ha2079a230000a797a4f70ea30000a717, /*  496 */
128'ha207a8230000a797a207a4230000a797, /*  497 */
128'ha007ac230000a797a207a2230000a797, /*  498 */
128'h0493f4bfe0ef8522e78d0009a783e4a9, /*  499 */
128'h3783020745630337971383093783680b, /*  500 */
128'hbfc5c4fff0effc075de3033797138309, /*  501 */
128'h84937bf050ef4501dff154fd000a2783, /*  502 */
128'h17b7b7d914fdb7e9c35ff0efbfc1710a, /*  503 */
128'he40616fd1141ff8006b78087b7033000, /*  504 */
128'h82e7b823f0070713670580e7b4238f75, /*  505 */
128'h7dc030efbac50513000095178307b583, /*  506 */
128'h300027f37d0030efbc85051300009517, /*  507 */
128'h07fe4785300790738fd9880707136709, /*  508 */
128'h7ac030efbc4505130000951734179073, /*  509 */
128'h014160a2302000730ff0000f0000100f, /*  510 */
128'h47838f5d07a200054703001547838082, /*  511 */
128'h25018d5d05628fd907c2003545030025, /*  512 */
128'h0005c703808200f61363367d57fd8082, /*  513 */
128'h1363367d57fdb7f5fee50fa305850505, /*  514 */
128'h1101495cbfcd050500b50023808200f6, /*  515 */
128'h3903cfa500958413e04ae426ec06e822, /*  516 */
128'h031348a5481586ca0200051347810185, /*  517 */
128'h146300a70e6327850006c703462d02e0, /*  518 */
128'h040500640023011795630e5007130107, /*  519 */
128'h00b94783fcc79ee30685040500e40023, /*  520 */
128'hc088f59ff0ef00f5842384ae01c90513, /*  521 */
128'h92238fd90087979b0189470301994783, /*  522 */
128'h8fd90087979b016947030179478300f4, /*  523 */
128'h690264a2644260e20004002300f49323, /*  524 */
128'h061302000593cf99873e611c80826105, /*  525 */
128'h869300c6986302d5fc630007468303a0, /*  526 */
128'hc683b7dd0705a00d577d00d706630017, /*  527 */
128'h66630ff6f593fd06869b577d46050007, /*  528 */
128'ha7178082853ae11c0006871b078900b6, /*  529 */
128'hc703cb85611cc915bfd586a747030000, /*  530 */
128'h02e69063008557030067d683c70d0007, /*  531 */
128'h00157793320060ef0017c503e4061141, /*  532 */
128'h808245258082014160a24525c3914501, /*  533 */
128'h8f5d0087979b468d01a5c70301b5c783, /*  534 */
128'h0145c6830155c78300d51d630007079b, /*  535 */
128'h853e27818fd90107979b8fd50087979b, /*  536 */
128'he84af4065904e44eec26f02271798082, /*  537 */
128'h8626468500154503842a03450993e052, /*  538 */
128'h02234c58505ce13125012ae060ef85ce, /*  539 */
128'h740270a2450100e7eb6340f487bb0004, /*  540 */
128'h00344903808261456a0269a2694264e2, /*  541 */
128'h9cbd4685001445034c5cff2a74e34a05, /*  542 */
128'hb7f94505b7e5397d26c060ef85ce8626, /*  543 */
128'h591c80824501f8dff06fc39900454783, /*  544 */
128'h02b787634401e04ae426ec06e8221101, /*  545 */
128'hc503ec190005041bfddff0ef892e84aa, /*  546 */
128'h25011f4060ef03448593864a46850014, /*  547 */
128'h644260e285220324a823597d4405c119, /*  548 */
128'he426ec06e822110180826105690264a2, /*  549 */
128'hfa3ff0ef842ad91c0005022357fde04a, /*  550 */
128'h979b45092324470323344783e52d2501, /*  551 */
128'h07134107d79b776d0107979b8fd90087, /*  552 */
128'h079bd59ff0ef06a4051302f71f63a557, /*  553 */
128'h049300544537fff50913010005370005, /*  554 */
128'h0864051300978c6345010127f7b31465, /*  555 */
128'h00a035338d05012575332501d33ff0ef, /*  556 */
128'hbfcd450d80826105690264a2644260e2, /*  557 */
128'hec56f052fc26e0a2e486f44ef84a715d, /*  558 */
128'hdd9ff0ef8932852e89aa00053023e85a, /*  559 */
128'h8793000097970035171302054e6347ad, /*  560 */
128'h0089b023c01547b184aa638097ba66e7, /*  561 */
128'h779313e060ef00144503cb8500044783, /*  562 */
128'h60a647a9c111891100090563e38d0015, /*  563 */
128'h853e6b426ae27a0279a2794274e26406, /*  564 */
128'h00a400a3000400230ff4f51380826161, /*  565 */
128'h00090463fb71478d00157713050060ef, /*  566 */
128'h1a634785ee1ff0ef85224581f5698911, /*  567 */
128'h478389a623a40a131fa40913848a04f5, /*  568 */
128'ha0232501c5bff0ef854ac7894501ffc9, /*  569 */
128'haa8301048913ff2a14e30991094100a9, /*  570 */
128'he9dff0ef852285d6000a876345090004, /*  571 */
128'h00e519634785470dfe9915e30491c10d, /*  572 */
128'h47b5c1194a81f6e504e34785470db7bd, /*  573 */
128'h8fd90087979b03f4470304044783bfb9, /*  574 */
128'hfef711e3200007134107d79b0107979b, /*  575 */
128'h00f9e9b30089999b04a4478304b44983, /*  576 */
128'h470501342e230444490329811a098663, /*  577 */
128'hfaf769e30ff7f793012401a3fff9079b, /*  578 */
128'hfffb079bfa0b03e30164012304144b03, /*  579 */
128'h1a1b0454478304644a03ffc900fb77b3, /*  580 */
128'hf3c100fa77930144142300fa6a33008a, /*  581 */
128'h0e638d450085151b0474448304844503, /*  582 */
128'h0087979b250104244703043447831405, /*  583 */
128'h9f3d004a571b2781033906bbdfb18fd9, /*  584 */
128'hd5bb40c504bbf4c564e3873200d7063b, /*  585 */
128'h00b93933664119556905dd8d84ae0364, /*  586 */
128'h248900ea873b490d00b6736309051655, /*  587 */
128'h470dd05c03542023cc04d458015787bb, /*  588 */
128'hb17ff0ef06040513f00a15e310e91263, /*  589 */
128'h24810094d49b1ff4849b0024949bd408, /*  590 */
128'h02a3f8000793c45cc81c57fdee99e7e3, /*  591 */
128'h064447030654478308f91963478d00f4, /*  592 */
128'h47054107d79b0107979b8fd90087979b, /*  593 */
128'h2501ce5ff0ef8522001a859b06f71b63, /*  594 */
128'h979b000402a32324470323344783e13d, /*  595 */
128'h07134107d79b776d0107979b8fd90087, /*  596 */
128'h57b7a99ff0ef0344051304f71263a557, /*  597 */
128'h2184051302f517632527879325014161, /*  598 */
128'h1c63272787932501614177b7a83ff0ef, /*  599 */
128'h22040513c808a6dff0ef21c4051300f5, /*  600 */
128'h27853f47d78300009797c448a63ff0ef, /*  601 */
128'h00f413233ef713230000971793c117c2, /*  602 */
128'h05840513b351478100042a2301240023, /*  603 */
128'hf0ef05440513b5b90005099ba33ff0ef, /*  604 */
128'h15634789d41c9fb5e00a05e3b545a25f, /*  605 */
128'h8885029787bb478db7010014949b00f9, /*  606 */
128'he426ec06e8221101bdc59cbd0017d79b, /*  607 */
128'h478d00044703ed692501bffff0ef842a, /*  608 */
128'h04930af71b634785005447030cf71063, /*  609 */
128'h0793a01ff0ef85264581200006130344, /*  610 */
128'h079322f409a3faa0079322f409230550, /*  611 */
128'h0b230610079302f40aa302f40a230520, /*  612 */
128'h02e40ba304100713481c20f40da302f4, /*  613 */
128'h0087571b0107571b0107971b20e40d23, /*  614 */
128'h0187d79b0107d71b20e40ea320f40e23, /*  615 */
128'h0107971b501020e40f23445c20f40fa3, /*  616 */
128'h07200693001445030087571b0107571b, /*  617 */
128'hd79b0107d71b260522e400a322f40023, /*  618 */
128'h01a322e4012320d40ca320d40c230187, /*  619 */
128'h000402a3599050ef85a64685d81022f4, /*  620 */
128'h3533250158d050ef4581460100144503, /*  621 */
128'h869b4d1c8082610564a2644260e200a0, /*  622 */
128'h85bb55480025458300f6f96337f9ffe5, /*  623 */
128'h0eb7f76347858082450180829d2d02d5, /*  624 */
128'h892ae44eec26f022f406e84a71794d18, /*  625 */
128'h06d70c63842e46890005470302e5f963, /*  626 */
128'h515c0015d49b00f71e6308d70e63468d, /*  627 */
128'hc9112501ac7ff0ef9dbd0094d59b9cad, /*  628 */
128'h6145853e69a2694264e2740270a257fd, /*  629 */
128'hf4930099d59b0014899b024927838082, /*  630 */
128'ha93ff0ef0344c483854a9dbd94ca1ff4, /*  631 */
128'h880503494783994e1ff9f993f5792501, /*  632 */
128'h157d6505bf658391c0198fc50087979b, /*  633 */
128'ha63ff0ef9dbd0085d59b515cbf458fe9, /*  634 */
128'h478399221fe474130014141bfd592501, /*  635 */
128'h515cb7598fc90087979b034945030359, /*  636 */
128'h151bf9352501a39ff0ef9dbd0075d59b, /*  637 */
128'h807ff0ef954a034505131fc575130024, /*  638 */
128'h8082853e4785b76517fd2501100007b7, /*  639 */
128'he852ec4ef426fc06f04a4540f8227139, /*  640 */
128'h450900f41c63892a478500b51523e456, /*  641 */
128'h61216aa26a4269e2790274a2744270e2, /*  642 */
128'hc683e02184aefee474e34f98611c8082, /*  643 */
128'h0087d703eb15579800e69463470d0007, /*  644 */
128'h0044d79bd171008928235788fce4f7e3, /*  645 */
128'h94be03478793049688bd000937839d3d, /*  646 */
128'hc9838722b75d450100993c2300a92a23, /*  647 */
128'h85a2000935034a8509925a7d843a0027, /*  648 */
128'he6fff0efbf752501e59ff0ef0134f663, /*  649 */
128'h00093783f68afbe301440c630005041b, /*  650 */
128'hb78d4505bfc1413484bbf6f476e34f9c, /*  651 */
128'hf0ef842aec06e426e822110100a55583, /*  652 */
128'h933ff0ef6008484ce4950005049bf33f, /*  653 */
128'hf0ef4581020006136c08ec990005049b, /*  654 */
128'h82234705601c00e7802357156c1cf3cf, /*  655 */
128'h71398082610564a28526644260e200e7, /*  656 */
128'h4a05e456ec4ef04af426f822fc06e852, /*  657 */
128'h47830af5f063498984aa4d1c16ba7563, /*  658 */
128'h8863470d0ae78f63842e893247090005, /*  659 */
128'h00ba0a3b515c0015da1b154794630ee7, /*  660 */
128'h96630005099b8b9ff0ef9dbd009a559b, /*  661 */
128'h1ffa7a130ff97793001a0a9b88050609, /*  662 */
128'hf71316c166850347c783014487b3cc19, /*  663 */
128'h9a260ff7f7938fd98ff50049179b00f7, /*  664 */
128'h009ad59b50dc00f48223478502fa0a23, /*  665 */
128'h00099f630005099b86bff0ef9dbd8526, /*  666 */
128'h9aa60ff979130049591bc40d1ffafa93, /*  667 */
128'h854e744270e200f482234785032a8a23, /*  668 */
128'h87b3808261216aa26a4269e2790274a2, /*  669 */
128'h9bc100f979130089591b0347c7830154, /*  670 */
128'hf0ef9dbd0085d59b515cb7e90127e933, /*  671 */
128'h74130014141bfc0992e30005099b811f, /*  672 */
128'h0109591b0109191b03240a2394261fe4, /*  673 */
128'h515cbf790144822303240aa30089591b, /*  674 */
128'h96e30005099bfd8ff0ef9dbd0075d59b, /*  675 */
128'h9aa603440a931fc474130024141bf809, /*  676 */
128'h69338d71f00006372501da0ff0ef8556, /*  677 */
128'h03240a230107d79b94260109179b0125, /*  678 */
128'h0189591b0109579b00fa80a30087d79b, /*  679 */
128'h7139bf3d4989b745012a81a300fa8123, /*  680 */
128'h84aae456e852f04af822fc06ec4ef426, /*  681 */
128'h77634d1c04090a6300c52903e19d89ae, /*  682 */
128'h04f4636324054c9c5afd4a05844a04f9, /*  683 */
128'h0005041bc43ff0efa8214401052a6063, /*  684 */
128'h8522547d00f41d6357fd0887f8634785, /*  685 */
128'h61216aa26a4269e2790274a2744270e2, /*  686 */
128'hbf554905b7d5faf47ee3894e4c9c8082, /*  687 */
128'h07e3c9012501c05ff0ef852685a24409, /*  688 */
128'h10000637b76dfb2411e305450863fd55, /*  689 */
128'h9063e9052501de9ff0ef852685a2167d, /*  690 */
128'hc89c37fdfae783e3577dc4c0489c0209, /*  691 */
128'h8622bf4900f482a30017e7930054c783, /*  692 */
128'h0fe34785dd612501dbbff0ef852685ce, /*  693 */
128'hfc0600a55903f04a7139bfad4405f6f5, /*  694 */
128'he456e852ec4ef426030917932905f822, /*  695 */
128'h69e2790274a2744270e24511eb9993c1, /*  696 */
128'h00f97993d7ed495c808261216aa26a42, /*  697 */
128'hc85c61082785480c00099d63842a8a2e, /*  698 */
128'h601cfcf775e30009071b00855783e18d, /*  699 */
128'h4501ec1c97ce03478793012415230996, /*  700 */
128'h0157fab337fd00495a9b00254783bf5d, /*  701 */
128'he46347850005049bb27ff0effc0a9fe3, /*  702 */
128'hb761450500f4946357fdbf4945090097, /*  703 */
128'hf0ef480cf60a0ee306f4e0634d1c6008, /*  704 */
128'hfcf48be34785d4bd451d0005049be81f, /*  705 */
128'hf5792501dd8ff0ef6008fcf48de357fd, /*  706 */
128'hbeeff0ef034505134581200006136008, /*  707 */
128'h02aa2823aa5ff0ef855285a600043a03, /*  708 */
128'h87bb591c00faed630025478360084a05, /*  709 */
128'hc848a83ff0ef85a6c8046008d91c4157, /*  710 */
128'h6018f1412501d1cff0ef01450223b7b9, /*  711 */
128'hf426f8227139b7e9db1c27855b1c2a85, /*  712 */
128'h0005c783e05ae456e852ec4ef04afc06, /*  713 */
128'h05c0071300e78663842e84aa02f00713, /*  714 */
128'h47fd000447030004a62304050ce79063, /*  715 */
128'h02e0099305c00a9302f00a130ae7fc63, /*  716 */
128'hb9030d5780630d478263000447834b21, /*  717 */
128'h4783b40ff0ef854a02000593462d0204, /*  718 */
128'h906300144783013900230d3792630004, /*  719 */
128'h8e630024478300f900a302e007930b37, /*  720 */
128'h05a302000793943a09479763470d1b37, /*  721 */
128'h100510632501adbff0ef8526458100f9, /*  722 */
128'h47836c98e96d2501cdaff0ef608848cc, /*  723 */
128'h8593709cef918ba100b74783c7e50007, /*  724 */
128'hc683fff74603078507050cb78d6300b7, /*  725 */
128'hbf75dfdff0ef85264581fed608e3fff7, /*  726 */
128'ha85ff0ef85264581b791c55c4bdc611c, /*  727 */
128'h69e2790274a2744270e20004bc232501, /*  728 */
128'h4709bf1d0405808261216b026aa26a42, /*  729 */
128'h943a12f6e06302000693f7578be3bf95, /*  730 */
128'h0313478145a147014681b7ad02400793, /*  731 */
128'h95130027e793a8dd0505a0d148650200, /*  732 */
128'h4711a06d268500e50023954a91010206, /*  733 */
128'h469500d515630e50069300094503c6ed, /*  734 */
128'h0ff7f7930027979b0165966300d90023, /*  735 */
128'h8bb10107671300b6946345850037f693, /*  736 */
128'h9432920116020087671300d794634691, /*  737 */
128'hc783709c4511bf654701bdfd00e905a3, /*  738 */
128'hf7930047f713f4e518e34711c50500b7, /*  739 */
128'he80703e30004bc230004a623cb890207, /*  740 */
128'h6c8cfbf58b91b73d4515fb0dbf154501, /*  741 */
128'hf0ef0007c503609cdbe58bc100b5c783, /*  742 */
128'hf7930027979b05659a63bdb9c4c8af2f, /*  743 */
128'h930117020017061b873245ad46a10ff7, /*  744 */
128'h04e3f94706e3f4e374e3000747039722, /*  745 */
128'h551b0187151b02b6f263fd370ae3f957, /*  746 */
128'h4883cfa505130000851700054c634185, /*  747 */
128'h051bbd6d4519f11710e3000886630005, /*  748 */
128'h7513f9f7051beea87ae30ff57513fbf7, /*  749 */
128'h0ff777130017e7933701eea866e30ff5, /*  750 */
128'hf406842ae44ee84aec26f0227179bdf9, /*  751 */
128'hc90de199484c49bd0e500913451184ae, /*  752 */
128'hc7036c1ce1292501afaff0ef6008a0b1, /*  753 */
128'h0327026303f7f79300b7c783c3210007, /*  754 */
128'h00979a630017b79317e18bfd03378063, /*  755 */
128'h8082614569a2694264e2740270a24501, /*  756 */
128'h00042a23d9452501c13ff0ef85224581, /*  757 */
128'he426ec06e82245811101bfe54511b7cd, /*  758 */
128'h484c0e500493e50d250188fff0ef842a, /*  759 */
128'h0007c7836c1ced092501a8cff0ef6008, /*  760 */
128'h2501bcdff0ef85224585cb9900978d63, /*  761 */
128'h64a2644260e2451d00f513634791dd79, /*  762 */
128'hf0ef842aec06e426e822110180826105, /*  763 */
128'ha42ff0ef6008484ce49d0005049bfa9f, /*  764 */
128'hf0ef4581020006136c08e0850005049b, /*  765 */
128'h4705601c82aff0ef462d6c08700c84cf, /*  766 */
128'h8082610564a28526644260e200e78223, /*  767 */
128'h740270a245098082450900b7ed634785, /*  768 */
128'h71794d1c808261456a0269a2694264e2, /*  769 */
128'h84ae842ae052e44ee84af406ec26f022, /*  770 */
128'h85a600f4fa634c1c59fd4a05fcf5fde3, /*  771 */
128'h4501000914630005091bec8ff0ef8522, /*  772 */
128'h852285a6460103390763fb490ce3bf75, /*  773 */
128'h278501378a63481cf15d25018afff0ef, /*  774 */
128'h049b00f402a30017e79300544783c81c, /*  775 */
128'hfc061028ec2a7139b7594505bf5d0009, /*  776 */
128'h97970405426383eff0eff42ee432e82e, /*  777 */
128'h6622631800a78733050e8da787930000, /*  778 */
128'h97aa00070023c319676200070023c319, /*  779 */
128'h080c460100f618634785cb114501e398, /*  780 */
128'h452d8082612170e22501a0eff0ef0828, /*  781 */
128'hf0d2f4cefca6e122e506f8ca7175bfe5, /*  782 */
128'h0005302314050d634925e42ee8daecd6, /*  783 */
128'h091b9d6ff0ef1028002c8a7984aa89b2, /*  784 */
128'hf0efe4be1028083c65a2140910630005, /*  785 */
128'h01c9f7934519e011e11964062501b6df, /*  786 */
128'h102800f516634791c54dc3e101f9fa13, /*  787 */
128'h77936406e949008a6a132501e75ff0ef, /*  788 */
128'h08a302100713046007937aa2cfcd008a, /*  789 */
128'h0823000407a30004072300f40ca300f4, /*  790 */
128'h05a300e40c2300040ba300040b2300e4, /*  791 */
128'h0fa300040f2300040ea300040e230004, /*  792 */
128'h0d234785fc9fe0ef85a2000ac5030004, /*  793 */
128'h099b00040aa300040a2300040da30004, /*  794 */
128'hab03855685ce04098b6300fa82230005, /*  795 */
128'h85da39fd7522e9112501e3fff0ef030a, /*  796 */
128'ha895892ac90d250183aff0ef01352623, /*  797 */
128'hf60981e30049f993e3d98bc500b44783, /*  798 */
128'he72d0107f71300b44783f565a0854921, /*  799 */
128'h008a7793e3ad8b85000984630029f993, /*  800 */
128'hf4800309a78385a279a2020a6a13c399, /*  801 */
128'he0ef0009c503000485a3d09c01448523, /*  802 */
128'h0069d783dbbfe0ef01c40513c8c8f33f, /*  803 */
128'h94230134b0230004ae230004a623c888, /*  804 */
128'h7a0679a6794674e6854a640a60aa00f4, /*  805 */
128'hb7d5491db7e54911808261496b466ae6, /*  806 */
128'hf0caf4a6fc86e4d6e8d2eccef8a27119, /*  807 */
128'h0006a023ec6ef06af466f862fc5ee0da, /*  808 */
128'h0005099be91fe0ef8ab6e4328a2e842a, /*  809 */
128'h0007899bc39d662200b4478300099863, /*  810 */
128'h6aa66a4669e6790674a6854e744670e6, /*  811 */
128'h808261096de27d027ca27c427be26b06, /*  812 */
128'h445c01042903160789638b8500a44783, /*  813 */
128'h0b930006091b00f67463893e40f907bb, /*  814 */
128'h77934458fa090ce35c7d03040b132000, /*  815 */
128'h0025478300975c9b6008120790631ff7, /*  816 */
128'heb11020c99630ffcfc930197fcb337fd, /*  817 */
128'h498900f405a3478900a7ec6347854848, /*  818 */
128'h01851763b7e52501bd6ff0ef4c0cb741, /*  819 */
128'h00043d83cc08b7a5498500f405a34785, /*  820 */
128'h000c861bd5792501b98ff0ef856e4c0c, /*  821 */
128'hc4b58d3a0007849b00a6073b0099579b, /*  822 */
128'hc503419684bb00f6f4639fb1002dc683, /*  823 */
128'hf94d25010a6050ef85d2863a86a6001d, /*  824 */
128'h41a507bb4c48c3850407f79300a44783, /*  825 */
128'h20000613910115020097951b0097fc63, /*  826 */
128'h020497930094949bc5ffe0ef955285da, /*  827 */
128'ha783c45c9fa54099093b445c9a3e9381, /*  828 */
128'h04e601634c50b70500faa0239fa5000a, /*  829 */
128'h4685001dc503c38d0407f79300a44783, /*  830 */
128'h00a44783f139250106c050efe43a85da, /*  831 */
128'h863a4685601c00f40523fbf7f7936722, /*  832 */
128'h2e23f1152501018050ef85da0017c503, /*  833 */
128'h40bb87bb1ff5f5930009049b444c01a4, /*  834 */
128'h95a28626030585930007849b0127f463, /*  835 */
128'hf0a27159b59d499dbf9dbd1fe0ef8552, /*  836 */
128'hf45ef85aeca6f486fc56e0d2e4cee8ca, /*  837 */
128'h8a2e842a0006a023e46ee86aec66f062, /*  838 */
128'h000997630005099bcb5fe0ef8ab68932, /*  839 */
128'h854e740670a60007899bc39d00b44783, /*  840 */
128'h7c027ba27b427ae26a0669a6694664e6, /*  841 */
128'h8b8900a44783808261656da26d426ce2, /*  842 */
128'h0b9304f76c630127873b445c18078f63, /*  843 */
128'h77930409046344585c7d03040b132000, /*  844 */
128'h0025478300975c9b6008140793631ff7, /*  845 */
128'hef01040c9a630ffcfc930197fcb337fd, /*  846 */
128'h05a3478902e798634705cb914581485c, /*  847 */
128'h0005079bd86ff0ef4c0cb759498900f4, /*  848 */
128'he79300a4478312f76a634818445cf3fd, /*  849 */
128'h05a3478501879763b79500f405230207, /*  850 */
128'h4783c85ce311cc1c4858bf99498500f4, /*  851 */
128'hc50346854c50601cc38d0407f79300a4, /*  852 */
128'h00a44783f969250170d040ef85da0017, /*  853 */
128'h856e4c0c00043d8300f40523fbf7f793, /*  854 */
128'h0099579b000c869bd159250197cff0ef, /*  855 */
128'h002dc703c4b58d320007849b00a6863b, /*  856 */
128'h86a6001dc503419704bb00f774639fb5, /*  857 */
128'h41a587bb4c4cf15125016bf040ef85d2, /*  858 */
128'h20000613918115820097959b0297f263, /*  859 */
128'hfbf7f79300a44783a4ffe0ef855a95d2, /*  860 */
128'h9a3e9381020497930094949b00f40523, /*  861 */
128'h9fa5000aa783c45c9fa54099093b445c, /*  862 */
128'h445c481800c78e634c5cbdd100faa023, /*  863 */
128'h623040ef85da4685001dc50300e7fa63, /*  864 */
128'h75130009049b444801a42e23fd092501, /*  865 */
128'h05130007849b0127f46340ab87bb1ff5, /*  866 */
128'h00a447839dbfe0ef952285d286260305, /*  867 */
128'h499db5f9c81cbf4100f405230407e793, /*  868 */
128'h2501acffe0ef842ae406e0221141bd2d, /*  869 */
128'h0407f793cf690207f71300a44783e175, /*  870 */
128'h030405930017c50346854c50601cc395, /*  871 */
128'hfbf7f79300a44783ed5525015e1040ef, /*  872 */
128'he15d2501b77fe0ef6008500c00f40523, /*  873 */
128'h481800e785a30207671300b7c703741c, /*  874 */
128'h00e78e230086d69b0106d69b0107169b, /*  875 */
128'h00d78f230187571b0107569b00d78ea3, /*  876 */
128'h8d2300078ba300078b23485800e78fa3, /*  877 */
128'h00e78a2327010107571b0107169b00e7, /*  878 */
128'h00e78aa30087571b0107571b0107171b, /*  879 */
128'h0086d69b00e78c23021007130106d69b, /*  880 */
128'h0007892300e78ca300d78da304600713, /*  881 */
128'h0523fdf7f793600800a44783000789a3, /*  882 */
128'he06f014160a2640200f50223478500f4, /*  883 */
128'he022114180820141640260a24505ebbf, /*  884 */
128'he0ef8522e9012501effff0ef842ae406, /*  885 */
128'h0141640260a200043023e11925019cbf, /*  886 */
128'h4a6395bfe0efec060028e42a11018082, /*  887 */
128'h610560e2450120a78323000087970005, /*  888 */
128'h1028002c4601e42a7159bfe5452d8082, /*  889 */
128'hec190005041bb3bfe0efeca6f486f0a2, /*  890 */
128'h0005041bcd2ff0efe4be1028083c65a2, /*  891 */
128'h70a68522cbd8575277a2e9916586e41d, /*  892 */
128'hcb998bc100b5c7838082616564e67406, /*  893 */
128'h4791b7c5c8c897bfe0ef0004c50374a2, /*  894 */
128'he506e42afca67175bfd94415fcf41ee3, /*  895 */
128'h460184ae00050023f0d2f4cef8cae122, /*  896 */
128'hecbe081ce5292501acdfe0ef1828002c, /*  897 */
128'h4a16c2be02f009934bdc597d842677e2, /*  898 */
128'h470300008717e50567a24501040a1263, /*  899 */
128'h80a303a0071300e780230307071b14e7, /*  900 */
128'h078d00e7812302f007130e94186300e7, /*  901 */
128'h7a0679a6794674e6640a60aa00078023, /*  902 */
128'hfd452501f89fe0ef1828458580826149, /*  903 */
128'h65c677e2f5552501e6eff0ef18284581, /*  904 */
128'he0ef18284581c2aa8cdfe0ef0007c503, /*  905 */
128'h2501e48ff0ef18284581f9492501f63f, /*  906 */
128'h25018a7fe0ef0007c50365c677e2e105, /*  907 */
128'hdd612501a9eff0ef1828458101450e63, /*  908 */
128'h1828100cb7594509f8e516e367a24711, /*  909 */
128'h973610949301020797134781f5cfe0ef, /*  910 */
128'h871b04e462630037871beb05fc974703, /*  911 */
128'h66a20206961300e586bb40f405bbfff7, /*  912 */
128'h01368023fff7c79301271a6396b29201, /*  913 */
128'h1088920102071613b7c12785b7319c3d, /*  914 */
128'h4545b7e900c68023377dfc964603962a, /*  915 */
128'h4703973692810204169367220789bddd, /*  916 */
128'hb709fe9465e3fee78fa3240507850007, /*  917 */
128'he456e852ec4efc06f04af426f8227139, /*  918 */
128'h000917630005091bfb4fe0ef84ae842a, /*  919 */
128'h854a744270e20007891bcf8900b44783, /*  920 */
128'h4818808261216aa26a4269e2790274a2, /*  921 */
128'h445884bae3918b8900a4478300977763, /*  922 */
128'hc81cfcf778e34818445ce4bd00042623, /*  923 */
128'h4481bf7d00f405230207e79300a44783, /*  924 */
128'h4783fc960ee34c50d3e51ff7f793445c, /*  925 */
128'h4685601cc3850407f7930304099300a4, /*  926 */
128'h4783ed51250126b040ef0017c50385ce, /*  927 */
128'h86264685601c00f40523fbf7f79300a4, /*  928 */
128'hcc44ed352501219040ef85ce0017c503, /*  929 */
128'h377dc7290097999b002547836008bf59, /*  930 */
128'h02c6ed630337563b0336d6bbfff4869b, /*  931 */
128'hd1c19c9dc45c27814c0c8ff9413007bb, /*  932 */
128'hf793c45c9fa5445c0499ea634a855a7d, /*  933 */
128'hd49bcd112501c87fe0ef6008d7b51ff4, /*  934 */
128'h059b814ff0efe595484cbfb19ca90094, /*  935 */
128'h490900f405a3478900f5976347850005, /*  936 */
128'h490500f405a3478500f5976357fdbded, /*  937 */
128'h8b89600800a44783b765cc0cc84cb5ed, /*  938 */
128'hbf6984cee5990005059bfddfe0efcb81, /*  939 */
128'hfabafee3fd4588e30005059bc4bfe0ef, /*  940 */
128'h413484bbcc0c445cfaf5fae34f9c601c, /*  941 */
128'he42ef822fc067139b7bdc45c013787bb, /*  942 */
128'h2501fe6fe0ef0828002c4601842ac52d, /*  943 */
128'hf0eff01c101ce01c852265a267e2e115, /*  944 */
128'h8bc100b5c783cd996c0ce529250197cf, /*  945 */
128'h0007c50367e2a02d000430234515e789, /*  946 */
128'h0067d7838522458167e2c448e30fe0ef, /*  947 */
128'hfcf50be347912501cbdfe0ef00f41423, /*  948 */
128'h4791bfdd452580826121744270e2f971, /*  949 */
128'he0ef842ae406e0221141b7c1fcf501e3, /*  950 */
128'h0141640260a200043023e1192501dbaf, /*  951 */
128'h892e842af406e84aec26f02271798082, /*  952 */
128'h458100091f63e8890005049bd98fe0ef, /*  953 */
128'h8526740270a20005049bc5ffe0ef8522, /*  954 */
128'h85224581022430238082614564e26942, /*  955 */
128'h00042a2302f5136347912501b32ff0ef, /*  956 */
128'hf8bfe0ef85224581c68fe0ef852285ca, /*  957 */
128'hd16dbf7d00042a2300f5166347912501, /*  958 */
128'h002c460184aee42aeca67159bf6584aa, /*  959 */
128'he00d0005041bedafe0eff486f0a21028, /*  960 */
128'h0005041b872ff0efe4be1028083c65a2, /*  961 */
128'hc10fe0ef102885a6c489cf816786e801, /*  962 */
128'hbfcd44198082616564e6740670a68522, /*  963 */
128'h002c46018b2ee42af85a8432f0a27159, /*  964 */
128'hf45efc56e4cee8caeca6f486e0d28522, /*  965 */
128'h000a1c6300050a1be7cfe0efec66f062, /*  966 */
128'h02f76263ffec871b481c01842c836000, /*  967 */
128'h69a6694664e68552740670a600fb2023, /*  968 */
128'h808261656ce27c027ba27b427ae26a06, /*  969 */
128'h59fd4481490902fb9f63478500044b83, /*  970 */
128'h093508632501a55fe0ef852285ca4a85, /*  971 */
128'hfef963e329054c1c2485e11109550863, /*  972 */
128'h202300f402a30017e793c80400544783, /*  973 */
128'h44814981490110000ab7504cb74d009b, /*  974 */
128'he0ef0015899b852200099e631afd4c09, /*  975 */
128'h200009930344091385cee9212501d10f, /*  976 */
128'h0087979b0009470300194783038b9163, /*  977 */
128'hfc0c94e33cfd39f909092485e3918fd9, /*  978 */
128'h015575332501abcfe0efe02e854ab745, /*  979 */
128'hb7494a05b7c539f109112485e1116582, /*  980 */
128'hec06e426e8221101bfad8a2abfbd4a09, /*  981 */
128'h4783e4910005049bbc4fe0ef842ae04a, /*  982 */
128'h69028526644260e20007849bcb9100b4, /*  983 */
128'hcf390027f71300a447838082610564a2, /*  984 */
128'h0523c8180207e793fed772e348144458, /*  985 */
128'h2a232501a58ff0ef484cef01600800f4, /*  986 */
128'he0ef4c0cbf7d84aa00a405a3c5390004, /*  987 */
128'hb7dd450502f9146357fd0005091b94df, /*  988 */
128'hf9792501b37fe0ef167d100006374c0c, /*  989 */
128'hb769449db7e12501a1cff0ef85ca6008, /*  990 */
128'hfcf96ae34d1c6008fcf900e345094785, /*  991 */
128'h46854c50601cdba50407f79300a44783, /*  992 */
128'hf55d2501648040ef030405930017c503, /*  993 */
128'h7175b7b100f40523fbf7f79300a44783, /*  994 */
128'hf8cafca6e122e5061008002c4605e42a, /*  995 */
128'he0be1008081c65a2e9052501ca0fe0ef, /*  996 */
128'h00b7c78345196786e1052501e3bfe0ef, /*  997 */
128'hf79300b5c483c59975e2eb890207f793, /*  998 */
128'h6149794674e6640a60aa451dcb810014, /*  999 */
128'h0005041bad8fe0ef0009450379028082, /* 1000 */
128'h0613fc878de301492783c89d88c1cc0d, /* 1001 */
128'hcaa200a8458996cfe0ef00a8100c0280, /* 1002 */
128'h836ff0ef00a84581f1612501951fe0ef, /* 1003 */
128'h9f5fe0ef1008faf518e34791d94d2501, /* 1004 */
128'hbf612501f20fe0ef7502e411f1552501, /* 1005 */
128'h7171b769d575250191cff0ef85a27502, /* 1006 */
128'he94aed26f506f1221028002c4605e42a, /* 1007 */
128'he8eaece6f0e2f4def8dafcd6e152e54e, /* 1008 */
128'h083c65a21c0414630005041bbd0fe0ef, /* 1009 */
128'h1c0409630005041bd67fe0efe4be1028, /* 1010 */
128'hf79300b7c783441967a61af417634791, /* 1011 */
128'h091bb45fe0ef4581752218079f630207, /* 1012 */
128'h57fd16f90f6344094785180902630005, /* 1013 */
128'h0005041ba98fe0ef752216f90b634405, /* 1014 */
128'he0ef85220109549b85ca742216041463, /* 1015 */
128'h00050c1b45812000061303440a13f6ef, /* 1016 */
128'he0ef855202000593462d898fe0ef8552, /* 1017 */
128'h949b0109199b0ff4fb1347c1248188cf, /* 1018 */
128'hd49b021007930109d99b02f40fa30104, /* 1019 */
128'h07930ff97a9304f4062302e00b930104, /* 1020 */
128'h061304f406a30084d49b0089d99b0460, /* 1021 */
128'h0723040405a30404052303740a230200, /* 1022 */
128'h85d2049404a305640423053407a30554, /* 1023 */
128'h468d05740aa3772280efe0ef05440513, /* 1024 */
128'h00f69363571400d6166357d200074603, /* 1025 */
128'h27810107d79b0107969b06f407234781, /* 1026 */
128'h0107d79b0106d69b0107979b06f40423, /* 1027 */
128'h06f404a306d407a30087d79b0086d69b, /* 1028 */
128'hf59fe0ef1028040b99634c8500274b83, /* 1029 */
128'h00e785a3752247416786e8350005041b, /* 1030 */
128'h00078b230460071300e78c2302100713, /* 1031 */
128'h01378da301578d2300e78ca300078ba3, /* 1032 */
128'he0ef00f50223478500978aa301678a23, /* 1033 */
128'h2823001c0d1b7522a82d0005041bd5af, /* 1034 */
128'hec090005041b8dcfe0ef019502230385, /* 1035 */
128'hfb93f61fd0ef3bfd8552458120000613, /* 1036 */
128'hf25fe0ef85ca7522441db7498c6a0ffb, /* 1037 */
128'h7ae66a0a69aa694a64ea740a70aa8522, /* 1038 */
128'h44218082614d6d466ce67c067ba67b46, /* 1039 */
128'h002c843284aee42aeca6f0a27159b7c5, /* 1040 */
128'h65a2e13125019cafe0eff48610284605, /* 1041 */
128'h67a6e9152501b65fe0efe4be1028083c, /* 1042 */
128'hc30d6706e39d0207f79300b7c7834519, /* 1043 */
128'h8c3d027474138c658cbd752200b74783, /* 1044 */
128'h2501c9efe0ef00f502234785008705a3, /* 1045 */
128'he02ee42a71718082616564e6740670a6, /* 1046 */
128'h964fe0efed26f122f5060088002c4605, /* 1047 */
128'hf4be008865a26786120796630005079b, /* 1048 */
128'h10079a630005079baf7fe0eff0be083c, /* 1049 */
128'h1007126302077713479900b7c7037786, /* 1050 */
128'hd0ef102805ad46550e058e63479165e6, /* 1051 */
128'h850ae49fd0ef10a8008c02800613e55f, /* 1052 */
128'he0ef10a865820c054d6347adf05fd0ef, /* 1053 */
128'h10a80ce793634711cbf90005079baadf, /* 1054 */
128'h0593464d648aefc50005079bdc5fe0ef, /* 1055 */
128'h640602814783e0dfd0ef00d4851302a1, /* 1056 */
128'hc78300f40223478500f485a30207e793, /* 1057 */
128'h450306f7086357d64736cbbd8bc100b4, /* 1058 */
128'he0ef85220005059bf2dfd0ef85a60004, /* 1059 */
128'hfc3fd0ef8522c5a547890005059bcaef, /* 1060 */
128'h0557468302e007936706efb10005079b, /* 1061 */
128'hd79b06f707230107969b57d602f69d63, /* 1062 */
128'h0107d79b0107979b06f7042327810107, /* 1063 */
128'h06f704a30086d69b0106d69b0087d79b, /* 1064 */
128'he24fe0ef008800f7022306d707a34785, /* 1065 */
128'h0005079bb50fe0ef6506e7910005079b, /* 1066 */
128'hbfcd47a18082614d853e64ea740a70aa, /* 1067 */
128'hec861028002c4605842ee42ae8a2711d, /* 1068 */
128'he4be1028083c65a2e9292501810fe0ef, /* 1069 */
128'h00b7c783451967a6e12925019abfe0ef, /* 1070 */
128'h752200645703cb856786eb950207f793, /* 1071 */
128'h0044570300e78ba30087571b00e78b23, /* 1072 */
128'h0223478500e78ca30087571b00e78c23, /* 1073 */
128'h80826125644660e62501ad6fe0ef00f5, /* 1074 */
128'h4601002c893284aee42ae0cae4a6711d, /* 1075 */
128'he0510005041bf9bfd0efec86e8a20828, /* 1076 */
128'he5592501ca8fe0efd20208284581c4b9, /* 1077 */
128'h462d75c2e93d2501b8ffe0ef08284585, /* 1078 */
128'h0200061346ad00b48713ca1fd0ef8526, /* 1079 */
128'h17820007869bfff6879bce8900070023, /* 1080 */
128'h0a63fec783e3177d0007c78397a69381, /* 1081 */
128'he0150005041be69fd0ef510c65620209, /* 1082 */
128'h00e684630005468304300793470d6562, /* 1083 */
128'h2023c29fd0ef953e0347879302700793, /* 1084 */
128'h80826125690664a6644660e6852200a9, /* 1085 */
128'hb7d5842abf550004802300f515634791, /* 1086 */
128'hd0efec86e8a21028002c4605e42a711d, /* 1087 */
128'h460100010c2366a2ec550005041bee3f, /* 1088 */
128'h0593eba10007c78397b6938102061793, /* 1089 */
128'h041bbd6fe0efda0210284581ea290200, /* 1090 */
128'he1792501abbfe0ef10284585e8410005, /* 1091 */
128'hbc7fd0ef082c462dc3dd650601814783, /* 1092 */
128'h8b230460071300e78c23021007136786, /* 1093 */
128'hb74d2605a06100e78ca300078ba30007, /* 1094 */
128'h9736930102079713fff6079bbf45863e, /* 1095 */
128'h43658e2e4781082cfeb706e300074703, /* 1096 */
128'hf9f7051b27850006c70348b107f00e93, /* 1097 */
128'h651793411742370100a36c6391411542, /* 1098 */
128'h00eef863a82100070f1b712505130000, /* 1099 */
128'hbfcdf36d80826125644660e685224419, /* 1100 */
128'hb7cdffe81be306080563000548030505, /* 1101 */
128'h00235795a885078500c6802300fe06b3, /* 1102 */
128'h041b8fefe0ef00f502234785752200f5, /* 1103 */
128'hdbd50181478302f51b634791b7c10005, /* 1104 */
128'h06136506f4450005041ba55fe0ef1028, /* 1105 */
128'hd0ef082c462d6506b07fd0ef45810200, /* 1106 */
128'hb751842abf1900e785a347216786ae5f, /* 1107 */
128'hf4c7e5e30585068500e58023f91780e3, /* 1108 */
128'h71e30007869b02000613472993811782, /* 1109 */
128'hbf89eaf71de30e50079301814703f8d7, /* 1110 */
128'h05c528830585230305452e0305052e83, /* 1111 */
128'h8646040502938f2ae44ae826ec221101, /* 1112 */
128'hc5b326af8f9300005f97887687f2869a, /* 1113 */
128'h000f2583000fa38300b647338dfd00c6, /* 1114 */
128'hff4fa3839db9007585bb0fc1008fa403, /* 1115 */
128'h0198581b0078159b0105883b004f2703, /* 1116 */
128'hc6339f3100f805bb0077073b0105e833, /* 1117 */
128'h00c6171b9e39008f23838e358e6d00f6, /* 1118 */
128'h83bb00c5873b008383bb8e590146561b, /* 1119 */
128'h86bb8ebd00cf24038ef900b7c6b300d3, /* 1120 */
128'h9fa100d3e6b30116969b00f6d39b0076, /* 1121 */
128'h77338f2d0007061b00d703bbffcfa403, /* 1122 */
128'h0167171b00a7579b9f3d8f2d9fa10077, /* 1123 */
128'h00e387bb0003869b0005881b0f418f5d, /* 1124 */
128'h00005f972ac5859300005597f45f17e3, /* 1125 */
128'h00d7cf332ac28293000052971e4f8f93, /* 1126 */
128'h0015c383000faf0301e6c73300cf7f33, /* 1127 */
128'h93aa038a0005c70300ef0f3b0025c403, /* 1128 */
128'ha70300ef0f3b942a040a4318972a070a, /* 1129 */
128'h01b8581b9e3900581f1b010f083b004f, /* 1130 */
128'hc6339f3100f80f3b010f68330003a703, /* 1131 */
128'h0096139b008fa7039e398e3d8e7501e7, /* 1132 */
128'h00cf03bb00c3e63340189eb90176561b, /* 1133 */
128'hc6b3fff5c4838efd007f46b305919f35, /* 1134 */
128'h941b94aa048affcfa7039eb90fc101e6, /* 1135 */
128'h00d3843b8ec140980126d69b9fb900e6, /* 1136 */
128'h9f3d0077473301e777330083c7339fb9, /* 1137 */
128'h861b000f081b8f5d0147171b00c7579b, /* 1138 */
128'h5f17f25599e300e407bb0004069b0003, /* 1139 */
128'h13838393000053978ffa1c2f0f130000, /* 1140 */
128'h942a040a00d7c2b30003a703010fc403, /* 1141 */
128'ha4039f21011fc4839f25400000c2c4b3, /* 1142 */
128'hc4830107083b40809e2194aa048a0043, /* 1143 */
128'h9e210107683301c8581b0048171b012f, /* 1144 */
128'h94aa00e2c2b3048a00f8073b0083a403, /* 1145 */
128'h013fc90300b6129b408000c2863b9ea1, /* 1146 */
128'h9c3500c702bb03c100c2e6330156561b, /* 1147 */
128'h9ea1090a0056c6b300e7c6b3ffc3a483, /* 1148 */
128'h000924830106d69b9fa50106941b992a, /* 1149 */
128'h9fa5005747330007081b00d2843b8ec1, /* 1150 */
128'h0f918f5d0177171b0097579b9f3d8f21, /* 1151 */
128'hf5f592e300e407bb0004069b0002861b, /* 1152 */
128'h45b38f5dfff647130b02829300005297, /* 1153 */
128'h9f2d022f4403021f43830002a70300d7, /* 1154 */
128'h040a418c95aa058a93aa038a020f4583, /* 1155 */
128'h0068171b0107083b0042a5839f2d942a, /* 1156 */
128'h073b0107683301a8581b0003a5839e2d, /* 1157 */
128'ha5839e2d8e3d8e59fff6c6139db100f8, /* 1158 */
128'he633400c9ead0166561b00a6139b0082, /* 1159 */
128'hfff7c593023f44839ead00c703bb00c3, /* 1160 */
128'h048a9db5ffc2a4038db902c10075e5b3, /* 1161 */
128'h40809fa18dd50115d59b94aa00f5969b, /* 1162 */
128'h9fa18f4dfff747130007081b00b385bb, /* 1163 */
128'h8f5d0157171b00b7579b9f3d00774733, /* 1164 */
128'h9de300e587bb0005869b0003861b0f11, /* 1165 */
128'h00d306bb00fe07bb010e883b6462f3ef, /* 1166 */
128'h64c2cd70cd34c97c0505282300c8863b, /* 1167 */
128'hf84afc26e0a2715d653c808261056922, /* 1168 */
128'h03f7f413ec56f052e486e45ee85af44e, /* 1169 */
128'h0b9304000b13e53c893289ae84aa97b2, /* 1170 */
128'h74639381178200078a1b408b07bb0400, /* 1171 */
128'h85ce020ada93020a1a9300090a1b00f9, /* 1172 */
128'h0933481020ef0144043b865600848533, /* 1173 */
128'h97824401852660bc0174176399d64159, /* 1174 */
128'h6ae27a0279a2794274e2640660a6b7c9, /* 1175 */
128'hf793f0227179653c808261616ba26b42, /* 1176 */
128'h00178513e84af406e44eec26842a03f7, /* 1177 */
128'h449d0400099300e7802397a2f8000713, /* 1178 */
128'h95224581920116020006091b40a9863b, /* 1179 */
128'h603cfc1c078e643c0124f5633c9020ef, /* 1180 */
128'h64e2740270a2fd24fde3450197828522, /* 1181 */
128'hd3078793000077978082614569a26942, /* 1182 */
128'hd287879300007797e93c04053423639c, /* 1183 */
128'h8082e13cb6c7879300000797ed3c639c, /* 1184 */
128'h3bf020efec06850a4641050505931101, /* 1185 */
128'h859300006597f6e68693000076974701, /* 1186 */
128'h070506890007c78300e107b345411a65, /* 1187 */
128'hc78397ae000646038bbd962e0047d613, /* 1188 */
128'h60e2fca71de3fef68fa3fec68f230007, /* 1189 */
128'he122717580826105f305051300007517, /* 1190 */
128'h85a26622f71ff0efe42ee5060808842a, /* 1191 */
128'hf0ef0808f01ff0ef0808e85ff0ef0808, /* 1192 */
128'h711c46a1595880826149640a60aaf83f, /* 1193 */
128'hcf980200071300d71763469100d70d63, /* 1194 */
128'h11018082556dbfe50007ac2380824501, /* 1195 */
128'h026384ae842a200007b7ec06e426e822, /* 1196 */
128'h659708800613e5e686930000569702f5, /* 1197 */
128'h30ef11a505130000651710a585930000, /* 1198 */
128'h11018082610564a2644260e2fc240f70, /* 1199 */
128'h026384ae200007b7ec06e4266100e822, /* 1200 */
128'h659702f00613e36686930000569702f4, /* 1201 */
128'h30ef0da50513000065170ca585930000, /* 1202 */
128'h11018082610564a2644260e2e0040b70, /* 1203 */
128'h026384ae200007b7ec06e4266100e822, /* 1204 */
128'h659703600613e06686930000569702f4, /* 1205 */
128'h30ef09a505130000651708a585930000, /* 1206 */
128'h11018082610564a2644260e2e4040770, /* 1207 */
128'h8263842e200007b7ec06e8226104e426, /* 1208 */
128'h659703e00613cae686930000769702f4, /* 1209 */
128'h30ef05a505130000651704a585930000, /* 1210 */
128'h610564a2644260e2e880900114020370, /* 1211 */
128'h200007b7ec06e8226104e42611018082, /* 1212 */
128'h0613c62686930000769702f48263842e, /* 1213 */
128'h05130000651700658593000065970450, /* 1214 */
128'h644260e2ec80900114027f2030ef0165, /* 1215 */
128'hec06e4266100e82211018082610564a2, /* 1216 */
128'h86930000569702f4026384ae200007b7, /* 1217 */
128'h6517fc2585930000659704c00613d4e6, /* 1218 */
128'h644260e2f0047ae030effd2505130000, /* 1219 */
128'hec06e4266100e82211018082610564a2, /* 1220 */
128'h86930000569702f4026384ae200007b7, /* 1221 */
128'h6517f82585930000659705300613d1e6, /* 1222 */
128'h644260e2f40476e030eff92505130000, /* 1223 */
128'hf82200053983ec4e71398082610564a2, /* 1224 */
128'h8436893284ae200007b7fc06f04af426, /* 1225 */
128'h05a00613ce4686930000569702f98463, /* 1226 */
128'hf485051300006517f385859300006597, /* 1227 */
128'h8b0589890014159b6722722030efe43a, /* 1228 */
128'he5b30034949b8dd9004979130029191b, /* 1229 */
128'h74a202b9b8238dc5744270e288a10125, /* 1230 */
128'h47057100e02211418082612169e27902, /* 1231 */
128'h8522f7dff0efe4064581852246054681, /* 1232 */
128'h45814605468547058522f35ff0ef4581, /* 1233 */
128'h640260a2d97ff0ef45816008f67ff0ef, /* 1234 */
128'h46814705e022e4061141808201414501, /* 1235 */
128'hf0ef842a45810405302302053c234605, /* 1236 */
128'h470545818522ef1ff0ef45818522f39f, /* 1237 */
128'h458160a264026008f23ff0ef46054685, /* 1238 */
128'hec06e8226104e4261101d4dff06f0141, /* 1239 */
128'h86930000569702f48263842e200007b7, /* 1240 */
128'h6517e52585930000659706100613c0e6, /* 1241 */
128'hfc809041144263e030efe62505130000, /* 1242 */
128'h6104e42611018082610564a2644260e2, /* 1243 */
128'h569702f48263842e200007b7ec06e822, /* 1244 */
128'h85930000659706800613bda686930000, /* 1245 */
128'h67855fa030efe1e5051300006517e0e5, /* 1246 */
128'h8082610564a2644260e2e0a08c7d17fd, /* 1247 */
128'h84ae200007b7ec06e4266100e8221101, /* 1248 */
128'h06f00613ba4686930000569702f40263, /* 1249 */
128'hdd85051300006517dc85859300006597, /* 1250 */
128'h8082610564a2644260e2e4245b4030ef, /* 1251 */
128'h07b7ec06e426e82200053903e04a1101, /* 1252 */
128'h86930000569702f9026384ae842a2000, /* 1253 */
128'h6517d82585930000659707600613b6e6, /* 1254 */
128'hc84404993c2356e030efd92505130000, /* 1255 */
128'hf0a2715980826105690264a2644260e2, /* 1256 */
128'hf85afc56e0d2e4cef486e8caeca67100, /* 1257 */
128'h892e0005d783020408a3ec66f062f45e, /* 1258 */
128'h20ef00c9051345814611d01ce03084b2, /* 1259 */
128'h3983bf5ff0ef458560080e049c636ca0, /* 1260 */
128'h278316f99a6304043a03200007b70004, /* 1261 */
128'he391448d8b89c7090017f71344810049, /* 1262 */
128'h2783000a09638cdd03243c234c1c4485, /* 1263 */
128'h468147050144e493160786638b85008a, /* 1264 */
128'hf0ef85224581d71ff0ef852245814605, /* 1265 */
128'hae8c0c1300005c17852200892583be1f, /* 1266 */
128'h0a1300006a17852200095583c4fff0ef, /* 1267 */
128'h4581cbdff0ef852285a6c81ff0efcaea, /* 1268 */
128'h85224581460546854705cf5ff0ef8522, /* 1269 */
128'hf0ef852224058593000f45b7d27ff0ef, /* 1270 */
128'h85220d89b583cd1ff0ef85224585e93f, /* 1271 */
128'h8993eb7ff0ef25810015e593009899b7, /* 1272 */
128'h70a6efe9485cc6ea8a9300006a976819, /* 1273 */
128'h7ba27b427ae26a0669a6694664e67406, /* 1274 */
128'he024852244cc8082616545016ce27c02, /* 1275 */
128'h8b85449cdf3ff0ef8522488cdb7ff0ef, /* 1276 */
128'h0107e683654100043883603cee079be3, /* 1277 */
128'h051300ff0e3743114701478145816390, /* 1278 */
128'h00371f1b00064803ec0689e36e89f005, /* 1279 */
128'h16fd060527810107e7b301e8183b0705, /* 1280 */
128'h67330187971b0187d81bf2e500670363, /* 1281 */
128'h67330087d79b01c878330087981b0107, /* 1282 */
128'h83751782170200be873b8fd98fe90107, /* 1283 */
128'h5697b765470147812585e31c97469381, /* 1284 */
128'h8593000065971490061398a686930000, /* 1285 */
128'hbd8537a030efb9e5051300006517b8e5, /* 1286 */
128'h1d633b7d20000bb78b4ebd6100c4e493, /* 1287 */
128'h05130000651796e5859300005597000b, /* 1288 */
128'h0179096300043903b7116f6000efb8e5, /* 1289 */
128'h348333a030ef855685d20f20061386e2, /* 1290 */
128'h370312048e6324818cfd4c81485c0709, /* 1291 */
128'h0793c7817c1c00f76f630c8937830209, /* 1292 */
128'h85224581b6fff0ef85224581cc5cf920, /* 1293 */
128'h852201442903c3950044f793b27ff0ef, /* 1294 */
128'h85cad47ff0ef85ca00896913ff397913, /* 1295 */
128'h0084f793680000efb305051300006517, /* 1296 */
128'h00496913ff397913852201442903c395, /* 1297 */
128'hb30505130000651785cad1fff0ef85ca, /* 1298 */
128'h390300043c83cfb50014f793658000ef, /* 1299 */
128'h06138da6869300005697017c8c630384, /* 1300 */
128'h2783cba97c1c28e030ef855685d209c0, /* 1301 */
128'h08e69f630037f693470d02043c230049, /* 1302 */
128'h63104591480d468100c90793018c8713, /* 1303 */
128'h370301068763c3900086161bff870513, /* 1304 */
128'h90e30791872a2685c3988f518361ff87, /* 1305 */
128'h485cc85c0027e793485ccbb5603cfeb6, /* 1306 */
128'h040439036004cc9d4c858889c85c9bf9, /* 1307 */
128'h0ca00613874686930000569701748c63, /* 1308 */
128'h0009096304043023210030ef855685d2, /* 1309 */
128'h485cb4dff0ef8522ef8d8b8500892783, /* 1310 */
128'h8ee3c47ff0ef8522484cc85c9bf54c85, /* 1311 */
128'hb783dbd98b85bd9560f020ef4505d80c, /* 1312 */
128'hbf41b1dff0ef8522b77100f92623000c, /* 1313 */
128'h8de394be00093c830109648397a667a1, /* 1314 */
128'he43e002c46218566639c00878913fa97, /* 1315 */
128'h08b041635535b7dd87ca0ca139a020ef, /* 1316 */
128'he44ef406e84aec26f022048005137179, /* 1317 */
128'h85a2cc1d5551842a100030ef892e84b2, /* 1318 */
128'h85aa89aa785010ef7e05051300004517, /* 1319 */
128'h8b634fe000ef9fe50513000065178622, /* 1320 */
128'hf793f40401242423e01c200007b70209, /* 1321 */
128'h64e2740270a24501c45c4789cb990024, /* 1322 */
128'h4785d4fd450188858082614569a26942, /* 1323 */
128'h8082bff9557d0e8030ef8522b7e5c45c, /* 1324 */
128'h200007b7f73ff06f2000053745814609, /* 1325 */
128'he0221141711c808225016108953e050e, /* 1326 */
128'h0000469702f40263200007b7e4066380, /* 1327 */
128'h8e0585930000659734c0061377c68693, /* 1328 */
128'h4505703c0cc030ef8f05051300006517, /* 1329 */
128'he822110180820141640260a2557de391, /* 1330 */
128'h644285a24d3010efe42eec064501842a, /* 1331 */
128'h051371797940006f6105468560e26622, /* 1332 */
128'h30efe052e44ee84aec26f022f4062000, /* 1333 */
128'h10e030ef954505130000651784aa0060, /* 1334 */
128'h842a491010ef450144b010ef0001b503, /* 1335 */
128'h638c93a5051300006517681c206010ef, /* 1336 */
128'h938505130000651706f445833f8000ef, /* 1337 */
128'hd59b9425051300006517546c3e8000ef, /* 1338 */
128'h06c44583583c3d2000ef91c115c20085, /* 1339 */
128'h0107d69b0087d71b9385051300006517, /* 1340 */
128'h0ff6f6930ff7f7930ff777130187d61b, /* 1341 */
128'h92850513000065175c0c3a6000ef2601, /* 1342 */
128'hc7898b25859300006597545c398000ef, /* 1343 */
128'h91850513000065178a05859300006597, /* 1344 */
128'h05e030ef9245051300006517378000ef, /* 1345 */
128'h2783db5fb0efe9658593000065977448, /* 1346 */
128'h6617e78987c6061300006617584c19c4, /* 1347 */
128'h00ef9025051300006517bda606130000, /* 1348 */
128'h6a174481ed5ff0ef84264581852633a0, /* 1349 */
128'h09139029899300006997902a0a130000, /* 1350 */
128'h30c000ef855285a6e78901f4f7932000, /* 1351 */
128'h00ef819100f5f6132485854e00044583, /* 1352 */
128'he205051300006517fd249fe304052fa0, /* 1353 */
128'h6a0269a2694264e2740270a22e8000ef, /* 1354 */
128'hb6830083b7830103b703808261454501, /* 1355 */
128'h00d7fe6393811782278540f707b30003, /* 1356 */
128'h0103b78300a7002300f3b82300170793, /* 1357 */
128'h0083b703808245018082000780234505, /* 1358 */
128'h0003b7038f999201020596130103b783, /* 1359 */
128'h9d9dfff7059b00c6f5638e9dfff70693, /* 1360 */
128'h002300b6e6630103b70340a786bb87aa, /* 1361 */
128'hc68300d3b823001706938082852e0007, /* 1362 */
128'h000556634881bfe900d7002307850007, /* 1363 */
128'h0693c21906100693488540a0053be681, /* 1364 */
128'h0005061b385986ba4e250ff6f8130410, /* 1365 */
128'h0305051b046e67630ff3751302b6733b, /* 1366 */
128'h8532fea68fa306850ff5751302b6563b, /* 1367 */
128'h876302f5e9630300051340e685bbfe71, /* 1368 */
128'h40e6853b068500f6802302d007930008, /* 1369 */
128'hfff5081b86ba2581000680230015559b, /* 1370 */
128'h8fa30685bf5d00a8053b808200b61b63, /* 1371 */
128'h97ba9381178240c807bbb7d92585fea6, /* 1372 */
128'h80230066802326050006c8830007c303, /* 1373 */
128'hf8a2597d011cf0ca7119b7f106850117, /* 1374 */
128'h843684b2e0dafc86e4d6e8d2eccef4a6, /* 1375 */
128'h06c00a1302500993f82af02ef42afc3e, /* 1376 */
128'h0004c50377a277420209591303000a93, /* 1377 */
128'hff639381178276820017079bc52d8f1d, /* 1378 */
128'he7bff0ef0201039304850135086304d7, /* 1379 */
128'h10634781048905450f630014c503bfe1, /* 1380 */
128'h0ff7f793fd07879bcb9d0004c7830355, /* 1381 */
128'h069304890014c503478100f6f36346a5, /* 1382 */
128'h0f630580069302a6eb6306d50f630640, /* 1383 */
128'h744670e6f55d08f509630630079304d5, /* 1384 */
128'h0007051b6b066aa66a4669e6790674a6, /* 1385 */
128'h07300713b74d048d0024c50380826109, /* 1386 */
128'hf6e51ee30700071300a76c6306e50e63, /* 1387 */
128'h07500713a00d46014685003800840b13, /* 1388 */
128'hfa850613f6e510e30780071302e50063, /* 1389 */
128'ha81145c1001636134685003800840b13, /* 1390 */
128'h46010016b693003800840b13f8b50693, /* 1391 */
128'h020103930005059be37ff0ef400845a9, /* 1392 */
128'h0201039300044503a809ddbff0ef0028, /* 1393 */
128'h00840b13b5fd845ad93ff0ef00840b13, /* 1394 */
128'h0005059b4db010ef8522012474336000, /* 1395 */
128'hec061034f436715db7f1852202010393, /* 1396 */
128'h60e2e8dff0efe436e4c6e0c2fc3ef83a, /* 1397 */
128'h05931014862ef436f032715d80826161, /* 1398 */
128'hf0efe436e4c6e0c2fc3ef83aec061000, /* 1399 */
128'hfe36fa32f62e710d8082616160e2e69f, /* 1400 */
128'he2baea22ee060808100005931234862a, /* 1401 */
128'h0808842ae3fff0efe436eec6eac2e6be, /* 1402 */
128'h691c80826135645260f285220f7020ef, /* 1403 */
128'h808245018302000303630087b303679c, /* 1404 */
128'h0713000047170205979304b7ee63479d, /* 1405 */
128'he426e822ec061101439c97ba83f92d67, /* 1406 */
128'h10ef7540f55c08c52483795c878297ba, /* 1407 */
128'h644260e202f457b39381020497930c50, /* 1408 */
128'h617cbfe97d5c808261054501e91c64a2, /* 1409 */
128'h557db7e9659c95aa058e05e135f1bfd9, /* 1410 */
128'hf0ef842ae406e02211418082557d8082, /* 1411 */
128'h07630207b303679c681c00055e63ff5f, /* 1412 */
128'h60a245018302014160a2640285220003, /* 1413 */
128'h00a7eb6347ad8082557d808201416402, /* 1414 */
128'h6108953e817525e78793000047971502, /* 1415 */
128'h679c691c80824fe50513000055178082, /* 1416 */
128'h47d502f1102347a1715d83020007b303, /* 1417 */
128'h07930030e83ee42e078517824785d23e, /* 1418 */
128'h60a6fd3ff0efcc3ed402e486100c2000, /* 1419 */
128'h450100e6fe63400407374d1480826161, /* 1420 */
128'h22813483230134032381308345018082, /* 1421 */
128'h041322813823dc010113808224010113, /* 1422 */
128'h348322113c232291342385a2980101f1, /* 1423 */
128'h0a0447830a04c703f579f95ff0ef1a05, /* 1424 */
128'h02f716630dd447830dd4c70302f71c63, /* 1425 */
128'h0e04c70302f710630c0447830c04c703, /* 1426 */
128'h85130d440593461100f71a630e044783, /* 1427 */
128'h7179b761fb600513d55156f010ef0d44, /* 1428 */
128'h85226b8020eff4063e800513842af022, /* 1429 */
128'hf21ff0efc202c40200011023858a4601, /* 1430 */
128'h70a2852269a020ef7d000513e509842a, /* 1431 */
128'h478500f1102347857179808261457402, /* 1432 */
128'h45386914c195842ac402c23ef406f022, /* 1433 */
128'h06b78ff58ff9f80787934ad4008007b7, /* 1434 */
128'h4601c43e8fd98f55400006b78f756000, /* 1435 */
128'h70a2c43c47b2e119ec9ff0ef8522858a, /* 1436 */
128'h47d500f1102347b5711d808261457402, /* 1437 */
128'h0107979bf852fc4ee0ca07c55783c23e, /* 1438 */
128'hec86f456e4a6e8a26a056989fdf94937, /* 1439 */
128'he0098993080909134495c43e842e8aaa, /* 1440 */
128'hed0de73ff0ef8556858a4601e00a0a13, /* 1441 */
128'h054793630135f7b3c7891005f79345b2, /* 1442 */
128'hf0ef35a5051300005517c78d0125f7b3, /* 1443 */
128'h79e2690664a6644660e6fba00513d4bf, /* 1444 */
128'h347dfe04c6e334fd808261257aa27a42, /* 1445 */
128'h5a6020ef3e80051300f057630014079b, /* 1446 */
128'h3305051300005517fc8049e34501b755, /* 1447 */
128'he7a919c52783bf7df9200513d09ff0ef, /* 1448 */
128'h858a460147d5c42e00f1102347c17139, /* 1449 */
128'hc11dde3ff0efc23e842af426fc06f822, /* 1450 */
128'h8522858a46014495cb918b891b842783, /* 1451 */
128'h74a2744270e2f8ed34fdc901dcdff0ef, /* 1452 */
128'he4a6711d80824501bfd5450180826121, /* 1453 */
128'h06d7f66384b6892a4785e8a2ec86e0ca, /* 1454 */
128'h08c92783260102f1102302c9270347c9, /* 1455 */
128'h100c47850030cc3ee42e4755d432cf31, /* 1456 */
128'he529842ad75ff0efc83eca26d23a854a, /* 1457 */
128'h47f5460102f1102347b10497f0634785, /* 1458 */
128'h5517c11dd55ff0efd23ed402854a100c, /* 1459 */
128'h644660e68522c43ff0ef28a505130000, /* 1460 */
128'h02f6063bbf6147c580826125690664a6, /* 1461 */
128'hfc067139b7c54401b7d50004841bb74d, /* 1462 */
128'h842ace05e456e852ec4ef04af426f822, /* 1463 */
128'hc11d892a482010ef8ab684b28a2e4148, /* 1464 */
128'h681000054d638dffa0ef852200b44583, /* 1465 */
128'h240505130000551700b67a63014485b3, /* 1466 */
128'hf0ef854a08c92583a0894481bd9ff0ef, /* 1467 */
128'hf3630207e4030109378389a6f96decdf, /* 1468 */
128'hf01ff0ef854a85d6865286a2844e0089, /* 1469 */
128'h84339a22408989b308c96783fc851ae3, /* 1470 */
128'h79028526744270e2fc0999e39aa20287, /* 1471 */
128'h47997139808261216aa26a4269e274a2, /* 1472 */
128'h030007b70086969bc23e47f500f11023, /* 1473 */
128'h84aafc06f426f8228ed10106161b8edd, /* 1474 */
128'he919c53ff0ef8526858a4601440dc436, /* 1475 */
128'h74a2744270e2d91ff0ef85263e800593, /* 1476 */
128'hdb0101134d18bfcdfc79347d80826121, /* 1477 */
128'h3023241134239fb923213823bffc07b7, /* 1478 */
128'h49013ffc07372331342322913c232481, /* 1479 */
128'hf0ef84aa85a2980101f104131ce7f563, /* 1480 */
128'h0513e7991a04b7831e051863892ac09f, /* 1481 */
128'h03631a04b5031aa4b0236c2020ef2000, /* 1482 */
128'h0c044783123010ef85a2200006131e05, /* 1483 */
128'h078ae0a70713000047171cf76b634721, /* 1484 */
128'hfd63cc981ff78793400407b753b897ba, /* 1485 */
128'hd69307a68007071367050d44278300e7, /* 1486 */
128'h09b449830a044783f8dc00d773630147, /* 1487 */
128'h0e244783e7810019f9938b8506f48f23, /* 1488 */
128'h478300098a6308f480a30b344783c789, /* 1489 */
128'h478306f48fa309c44783c7898b890a04, /* 1490 */
128'h4783fcdc07c60c848613091407130e24, /* 1491 */
128'hfff74783e0fc07c6468109d405130a84, /* 1492 */
128'h45839fad0105959b0087979b00074583, /* 1493 */
128'h0e04458300098c634685c39197aeffe7, /* 1494 */
128'he21c07ce02b787b30dd4478302f585b3, /* 1495 */
128'h08e4478304098f63fca714e30621070d, /* 1496 */
128'h9fb90087171b0107979b468508d44703, /* 1497 */
128'h478302f707330e04470397ba08c44703, /* 1498 */
128'h470308b44783f8fc07ce02e787b30dd4, /* 1499 */
128'h089447039fb90107171b0187979b08a4, /* 1500 */
128'hf4fc54d89fb9088447039fb90087171b, /* 1501 */
128'h4783c7898b850a044783f4fc07a6c319, /* 1502 */
128'h45850af006134685ce81e3918bfd09c4, /* 1503 */
128'h47830af407a34785ed35e0bff0ef8526, /* 1504 */
128'haa2300a6979bc7b98b850e0446830af4, /* 1505 */
128'h07a60d44278300098663c79954dc08f4, /* 1506 */
128'hac2302f686bb00a6969b0dd44783f8dc, /* 1507 */
128'h34032481308308f480230a74478308d4, /* 1508 */
128'h228139832301390323813483854a2401, /* 1509 */
128'h0057d79b00a7d71b50fc808225010113, /* 1510 */
128'h08f4aa2302f707bb278527058bfd8b7d, /* 1511 */
128'hb023524020efd1691a04b503892abf4d, /* 1512 */
128'hdc010113bf455929bf555951bf651a04, /* 1513 */
128'h23213023229134232281382322113c23, /* 1514 */
128'h54a9c585468102b7e16302f588634789, /* 1515 */
128'h34832201390385262301340323813083, /* 1516 */
128'h60e34705ffc5879b8082240101132281, /* 1517 */
128'hf0ef892a45850b900613842e4685fef7, /* 1518 */
128'hf1e9258199f5ffe4059bf57184aad1ff, /* 1519 */
128'he51998dff0ef854a85a2980101f10413, /* 1520 */
128'hb74d84aab75ddf400493f7d50b944783, /* 1521 */
128'h08154783f022f406e44ee84aec267179, /* 1522 */
128'h06138edd892e9be10079f6930ff5f993, /* 1523 */
128'h842a57b5c519cc7ff0ef84aa45850b30, /* 1524 */
128'h875ff0ef852685ca00091c6300f51e63, /* 1525 */
128'h70a28522013505a315e010ef8526842a, /* 1526 */
128'hd60101138082614569a2694264e27402, /* 1527 */
128'h29213023289134232881382328113c23, /* 1528 */
128'h27613023275134232741382327313c23, /* 1529 */
128'h25a13023259134232581382325713c23, /* 1530 */
128'hbffc07b74d180ac7e963478923b13c23, /* 1531 */
128'h892abfe787933ffc07b79f3dbff7879b, /* 1532 */
128'h00e7eb63e44505130000551784ae8b32, /* 1533 */
128'h051300005517e7b90016779307e94603, /* 1534 */
128'h298130838522f8400413f96ff0efe665, /* 1535 */
128'h27813983280139032881348329013403, /* 1536 */
128'h25813b8326013b0326813a8327013a03, /* 1537 */
128'h23813d8324013d0324813c8325013c03, /* 1538 */
128'h0513000055170989270380822a010113, /* 1539 */
128'h02eaf7bb060a81630045aa83db45e3e5, /* 1540 */
128'h00005517cb8902ecf7bb0005ac83e791, /* 1541 */
128'h02c92783bf415429f24ff0efe4450513, /* 1542 */
128'h88138c0a009c9c9be3994b8502eadabb, /* 1543 */
128'h000828834e114e85478189d6856200c4, /* 1544 */
128'h0000551700030d6302e8f33b0017859b, /* 1545 */
128'h4b814a814c81b7c1ee4ff0efe3c50513, /* 1546 */
128'h078e020880630065202302e8d33bb7f1, /* 1547 */
128'hebb300be96bbcb898b850107c78397a6, /* 1548 */
128'h87ae05110821013309bb0ffbfb9300db, /* 1549 */
128'h0513000055178a09000b8963fbc596e3, /* 1550 */
128'h85d2fe0a7a1302f10a13f00600e3e1e5, /* 1551 */
128'h09fa4603ee0519e3842af94ff0ef854a, /* 1552 */
128'h47839e3d0087979b0106161b09ea4783, /* 1553 */
128'h05130000551785ce01367a63963e09da, /* 1554 */
128'h0a7a46830084c783b5c1e56ff0efe0e5, /* 1555 */
128'hc3990fe6f9938b89c71989b60017f713, /* 1556 */
128'h070e0017059b4611450547010016e993, /* 1557 */
128'h02080463001878130017581b4b189726, /* 1558 */
128'h0189999b0187979b0027571b00b517bb, /* 1559 */
128'h00f9e9b3c70d4189d99b4187d79b8b05, /* 1560 */
128'h478302d98263fcc592e3872e0ff9f993, /* 1561 */
128'h20efdc25051300005517ef898b850a6a, /* 1562 */
128'h4783bfd100f9f9b3fff7c793b5912cc0, /* 1563 */
128'hf0efdf25051300005517cb898b8509ba, /* 1564 */
128'h8b850afa4783e20b02e3b51d547ddbaf, /* 1565 */
128'ha21ff0ef854a45850af006134685e395, /* 1566 */
128'h00a7979b0e0a47830afa07a34785e569, /* 1567 */
128'hd6bb08c00d934d010880049308f92a23, /* 1568 */
128'h9f1ff0ef854a458586260ff6f69301ac, /* 1569 */
128'h4c81ffb492e32d210ff4f4932485ed49, /* 1570 */
128'h458586260ff6f693019ad6bb08f00d13, /* 1571 */
128'h2ca10ff4f4932485e9359cbff0ef854a, /* 1572 */
128'h26834c818aa609b00d934d61ffa492e3, /* 1573 */
128'h854a0ff6f6930196d6bb45858656000c, /* 1574 */
128'h90e30ffafa932ca12a85e13999dff0ef, /* 1575 */
128'h86defdb498e30c110ff4f493248dffac, /* 1576 */
128'h4785ed19975ff0ef854a458509c00613, /* 1577 */
128'h0613468501379b630a7a4783d4fb0de3, /* 1578 */
128'h86cebb3d842a957ff0ef854a458509b0, /* 1579 */
128'hdd79842a945ff0ef854a45850a700613, /* 1580 */
128'h5e63810ff0ef842ae406e0221141b32d, /* 1581 */
128'h8522000307630187b303679c681c0005, /* 1582 */
128'h0141640260a245058302014160a26402, /* 1583 */
128'h84aa4791f04af822fc06f42671398082, /* 1584 */
128'h0370079304f592635529478500f58663, /* 1585 */
128'h0107979b4955842e07c4d78300f11023, /* 1586 */
128'hed19d52ff0efc43ec24a8526858a4601, /* 1587 */
128'h478900f41f634791c24a00f110234799, /* 1588 */
128'h744270e2d34ff0ef8526858a4601c43e, /* 1589 */
128'hc402fef414e3478580826121790274a2, /* 1590 */
128'h4f1887ae00f5f3634f5c6918ee09b7cd, /* 1591 */
128'h0823dd0c0007059b00e7f46385be2781, /* 1592 */
128'h10000737691c80828082c2cff06f02c5, /* 1593 */
128'heccef0caf4a6fc86f8a2070d4b9c7119, /* 1594 */
128'hc17c8fd9f466f862fc5ee0dae4d6e8d2, /* 1595 */
128'heb8d6b9c679c681cc509f11ff0ef842a, /* 1596 */
128'hbacff0efc04505130000551702042423, /* 1597 */
128'h69e674a679068526744670e6f8500493, /* 1598 */
128'h808261097ca27c427be26b066aa66a46, /* 1599 */
128'h1af42c23478df93ff0eff3e54481541c, /* 1600 */
128'hba2ff0ef852202042c2302f408234785, /* 1601 */
128'h6b9c679c8522681c3ef010ef7d000513, /* 1602 */
128'h282318042e2308842783f94584aa9782, /* 1603 */
128'hb72ff0ef8522d85c478508f422231a04, /* 1604 */
128'hcf2ff0ef8522f1dff0ef852245814601, /* 1605 */
128'h47a1000505a345d000ef8522f14984aa, /* 1606 */
128'h07138ff94bdc00ff8737681c00f11023, /* 1607 */
128'h8522858a460147d50aa00713e3991aa0, /* 1608 */
128'h079300c14703e911bf8ff0efc23ec43a, /* 1609 */
128'h3e900913cc1c800207b700f715630aa0, /* 1610 */
128'h00ff8bb74b0502900a934a5503700993, /* 1611 */
128'h10238522858a460140000cb780020c37, /* 1612 */
128'h4c18681ce13dbb6ff0efc402c2520131, /* 1613 */
128'h1563c43e0177f7b3c25a4bdc01511023, /* 1614 */
128'hf0ef8522858a4601c43e0197e7b30187, /* 1615 */
128'h06090863397d0007ca6347b2ed1db8ef, /* 1616 */
128'h800207374c14bf452ff010ef3e800513, /* 1617 */
128'h41e7d79bc43ccc188001073700e68563, /* 1618 */
128'hb55d18f40ca3478506041e23d45c8b85, /* 1619 */
128'h4581c04ff0ef852202f51f63f9200793, /* 1620 */
128'h47850007d663443ced09c34ff0ef8522, /* 1621 */
128'hd965c1cff0ef85224585bfd118f40c23, /* 1622 */
128'hfa100493a10ff0efa805051300005517, /* 1623 */
128'hef26f706f3227161551cb58584aab595, /* 1624 */
128'heee6f2e2f6defadafed6e352e74eeb4a, /* 1625 */
128'h1cd010ef45018baae3b54401e6eeeaea, /* 1626 */
128'he7b5180b8ca3198bc783c7b1199bc783, /* 1627 */
128'hc2be855e008c479d460104f110234789, /* 1628 */
128'h1b8ba783120500e3842aabaff0efc482, /* 1629 */
128'haa0ff0ef855e008c46014495cf818b85, /* 1630 */
128'ha031020ba423f4fd34fd100503e3842a, /* 1631 */
128'h741a70ba8522d55d842ad99ff0ef855e, /* 1632 */
128'h7c167bb67b567af66a1a69ba695a64fa, /* 1633 */
128'h8c23048ba7838082615d6db66d566cf6, /* 1634 */
128'h10ef4501b16ff0ef855e0407c163180b, /* 1635 */
128'h855e45853e80091390810205149313b0, /* 1636 */
128'h0007cc63048ba783f155842ab36ff0ef, /* 1637 */
128'h10ef0640051312a96ee3117010ef8526, /* 1638 */
128'h048ba78300fbac23400007b7bfe91a50, /* 1639 */
128'h06fb9e23478502fba6238b8541e7d79b, /* 1640 */
128'h06370ea61ee345111aa60f63450dbf05, /* 1641 */
128'h00cbac234006061b40010637a0294004, /* 1642 */
128'h8a3d41a98993000039978a9d0036d61b, /* 1643 */
128'h45051086a6830f86460396ce964e068a, /* 1644 */
128'ha8238a0500c7d61b02d606bb018ba883, /* 1645 */
128'ha22308dba42304cba823180bae231a0b, /* 1646 */
128'h090ba62300d5183b8abd0107d69b08db, /* 1647 */
128'h14068e6302cba683090ba8231408dc63, /* 1648 */
128'h8fd98ff50107571b003f06b70107979b, /* 1649 */
128'h87b300e797b307090785472193811782, /* 1650 */
128'hb8230c0bb4230c0bb0230a0bbc230307, /* 1651 */
128'h07930afbb8230e0bb0230c0bbc230c0b, /* 1652 */
128'h0793090ba70308fba6230107d4632000, /* 1653 */
128'h04cba783c21508fba82300e7f4632000, /* 1654 */
128'h008c46010107979b471100e78e63577d, /* 1655 */
128'h479d902ff0efc282c4be04e11023855e, /* 1656 */
128'h0107979b4601495507cbd78304f11023, /* 1657 */
128'h16e3842a8e4ff0efc4bec2ca855e008c, /* 1658 */
128'h855e08fb80a357fd08fbaa234785e405, /* 1659 */
128'h0f7000ef855ee2051ae3842ac9aff0ef, /* 1660 */
128'he0051fe3842affbfe0ef855e00b54583, /* 1661 */
128'ha0232789100007b754075a63018ba703, /* 1662 */
128'h460107cbd78306f110230370079304fb, /* 1663 */
128'h880ff0efd4bed2ca855e0107979b108c, /* 1664 */
128'h1a93033007930bf104934905d2caed05, /* 1665 */
128'h4b210a854a11d48206f1102398810209, /* 1666 */
128'h850ff0efd05aec56e826855e108c0810, /* 1667 */
128'h40020637bb45842afe0a16e33a7dc131, /* 1668 */
128'h15bb89bd0165d59bbd9940030637a7a9, /* 1669 */
128'h0027979b16f16685b54d08bba82300b5, /* 1670 */
128'h938100f7571b17828fd501e7569b8ff5, /* 1671 */
128'h179b0187569b00ff05374098b5558b1d, /* 1672 */
128'h67410087569b8e698fd50087161b0187, /* 1673 */
128'h04fbaa2327818fd58ef1f00706138fd1, /* 1674 */
128'h0087159b8ecd0187169b0187559b40d8, /* 1675 */
128'h04ebac238f558f718ecd0087571b8de9, /* 1676 */
128'h20d702634689212700638b3d0187d71b, /* 1677 */
128'h0007596302d7971300ebac2380010737, /* 1678 */
128'ha70304fba0238fd920000737040ba783, /* 1679 */
128'h8793000057971ef71863800107b7018b, /* 1680 */
128'h044ba783f0be4d05040ba903639ce1e7, /* 1681 */
128'h00f979332344849300003497020d1a13, /* 1682 */
128'h40980a05fe07fc1383f979130ff10793, /* 1683 */
128'h16078563278100f977b300e797bb4785, /* 1684 */
128'hac8397d6109c840b0b1b4a81017d8b37, /* 1685 */
128'h140781630197f7b300f977b340dc0007, /* 1686 */
128'h4591200007b700fc8d6345a1400007b7, /* 1687 */
128'h0015b59340bc85b3100005b700fc8863, /* 1688 */
128'h400007370e051c638daa971ff0ef855e, /* 1689 */
128'h00ec886347912000073700ec8d6347a1, /* 1690 */
128'h02fbaa23001cb79340fc8cb3100007b7, /* 1691 */
128'h9163470d01a78663409cdfdfe0ef855e, /* 1692 */
128'h07b7d33e47d50af1102347994d850ce7, /* 1693 */
128'h07930110d53e00fde7b317c12d818100, /* 1694 */
128'he91fe0efc93ee552e162855e110c0400, /* 1695 */
128'ha823409c09b794638bbd010c4783e941, /* 1696 */
128'h0017b79317ed088ba58314079a631afb, /* 1697 */
128'h947ff0ef855e460118fbae2308bba223, /* 1698 */
128'h0af1102303700793fe07fd930ff10793, /* 1699 */
128'h855e110c0107979b4601475507cbd783, /* 1700 */
128'h6702e915e35fe0efd53ee03ad33a8cee, /* 1701 */
128'h040007134791d502d33a0af1102347b5, /* 1702 */
128'he03ac93ae552e16ee43e855e110c0110, /* 1703 */
128'hf3ed37fd670267a20e050c63e0dfe0ef, /* 1704 */
128'hae23096ba2231afba823017d85b74785, /* 1705 */
128'h0a918c9ff0ef855e840585934601180b, /* 1706 */
128'h0b0787930000379704a1eafa94e347a1, /* 1707 */
128'hcbdfe0ef55c5051300004517e6f49fe3, /* 1708 */
128'hb519a007071b80011737b61ddf400413, /* 1709 */
128'hde075ee30307971300ebac2380020737, /* 1710 */
128'h01000ab70ff104934905bbc580030737, /* 1711 */
128'h020a08633a7d09053ac54a1598811902, /* 1712 */
128'h040007931030c33e47d508f110234799, /* 1713 */
128'hd61fe0efdc3ef84af426c556855e010c, /* 1714 */
128'h66c144dcfbe18b8583a54cdcd0051ce3, /* 1715 */
128'h8fd18ff50087d79b0087961bf0068693, /* 1716 */
128'h00876793da06d9e3040ba70302e79693, /* 1717 */
128'h9713eaf768e34581472db35d04fba023, /* 1718 */
128'h859366c1b54511872583974e83790207, /* 1719 */
128'h0d91000da783f006869300ff0537040d, /* 1720 */
128'h8e690087961b8f510187971b0187d61b, /* 1721 */
128'h9ee3fefdae238fd98ff58f510087d79b, /* 1722 */
128'hf8638bbd00c7579b46a5008ca703fdb5, /* 1723 */
128'h369704d61c63800306b7018ba60300f6, /* 1724 */
128'h171b1487a78397b6078af02686930000, /* 1725 */
128'h8ff917fd67c100cca68308fbae230087, /* 1726 */
128'h03f7771327810126d71b8fd10186d61b, /* 1727 */
128'h0106d69b02e6073b3e800613c305c38d, /* 1728 */
128'ha2230afba02302d606bb02f757bb8a8d, /* 1729 */
128'hc79919cba7831afbaa231b0ba7830adb, /* 1730 */
128'h00ef855e08fba82308fba62320000793, /* 1731 */
128'hb7b708cba70300050623000515234840, /* 1732 */
128'h8ff9ccc68693aaa78793ccccd6b7aaaa, /* 1733 */
128'h9fb500f037b3068600d036b327818ef9, /* 1734 */
128'h068a00d036b38ef90f068693f0f0f6b7, /* 1735 */
128'h00d036b38ef9f0068693ff0106b79fb5, /* 1736 */
128'h00e037338f750207161376c19fb5068e, /* 1737 */
128'hd7b3ed1092010a8bb783d11c9fb90712, /* 1738 */
128'h84aa06fbc603074bd68307abd70302c7, /* 1739 */
128'hfef53623024505133985859300004597, /* 1740 */
128'h06cbc603077bc883070ba803a95fe0ef, /* 1741 */
128'h0ff7f7930188569b0108571b0088579b, /* 1742 */
128'h85930000459726810ff777130ff87813, /* 1743 */
128'h4597074ba603a5ffe0ef04d485133765, /* 1744 */
128'h561b0106569b06248513372585930000, /* 1745 */
128'h740010ef8526a3ffe0ef8a3d8abd0146, /* 1746 */
128'ha0232785100007b7b8d102fba4234785, /* 1747 */
128'he691ecf76ce31a0bb683400407b704fb, /* 1748 */
128'h079b70000737bb952f05051300004517, /* 1749 */
128'ha42303f7f6930c46c78304fba0230017, /* 1750 */
128'h071bc68900c7f693ce910027f6931adb, /* 1751 */
128'ha02301076713040ba70304eba0230217, /* 1752 */
128'ha02300c7e793040ba783c7998b8504eb, /* 1753 */
128'h4601088ba583044ba783040baa0304fb, /* 1754 */
128'hf0efdb2484930000349700fa7a33855e, /* 1755 */
128'h3c974c2ddc4b0b1300003b174a85db4f, /* 1756 */
128'h00fa77b300fa97bb409cdf6c8c930000, /* 1757 */
128'h20000d37da49091300003917cbb52781, /* 1758 */
128'h0017b79317ed00494703409c10000db7, /* 1759 */
128'h8ff900fa77b30009270340dc04f71863, /* 1760 */
128'h0fb6f69345850b70061300894683c3a1, /* 1761 */
128'h45850b7006134681c131debfe0ef855e, /* 1762 */
128'hae231a0ba823088ba783ddbfe0ef855e, /* 1763 */
128'h973fe0ef855e035baa2308fba223180b, /* 1764 */
128'h00004517f7649fe304a1fb9911e30931, /* 1765 */
128'h06b700092783bb6d925fe0ef1c450513, /* 1766 */
128'h87b301a78663471100d7896347214000, /* 1767 */
128'h933fe0ef855e02ebaa230017b71341b7, /* 1768 */
128'hf79300892683f941808ff0ef855e408c, /* 1769 */
128'h088ba583ef8d1afba823409ce79d0046, /* 1770 */
128'h460118fbae2308bba2230017b79317ed, /* 1771 */
128'hbb91fd319fdfe0ef855ecb0ff0ef855e, /* 1772 */
128'hd31fe0ef855e45850b7006130ff6f693, /* 1773 */
128'h837902079713fcfc65e34581b7c9f521, /* 1774 */
128'h06cb851300ec4641bf6d11872583974e, /* 1775 */
128'h460107cbd78304f11023478d6da000ef, /* 1776 */
128'he0efc2be47d5855ec4be0107979b008c, /* 1777 */
128'h0007d663018ba783ec051b63842a96ff, /* 1778 */
128'h479d04f1102347a506fb9e2304e15783, /* 1779 */
128'h855e0107979b008c460107cbd783c2be, /* 1780 */
128'h47c646b6ea051163842a93bfe0efc4be, /* 1781 */
128'h06fba02304dbae23018ba50345e64756, /* 1782 */
128'hf2c51a634000063706bba42306eba223, /* 1783 */
128'hf0c543638ca602e345098a3d01a6d61b, /* 1784 */
128'hf06f2006061b40010637f0a609634505, /* 1785 */
128'h80824501c56ce54ff06ffa100413f0ef, /* 1786 */
128'h5797808218b50d238082557d8082557d, /* 1787 */
128'he02247851141ef9d439c9f6787930000, /* 1788 */
128'h12a000ef9ef7202300005717842ae406, /* 1789 */
128'hfc5ff0ef852200055563aeefe0ef8522, /* 1790 */
128'h640260a20dc000ef13e000ef02c00513, /* 1791 */
128'h07130000571780824501808201414501, /* 1792 */
128'h451785aa114102e790636394631c9ae7, /* 1793 */
128'h478160a2f60fe0efe406172505130000, /* 1794 */
128'h87b600a604630fc7a60380820141853e, /* 1795 */
128'hf0efe42eec06110141488082853ebfd1, /* 1796 */
128'h470302b7006365a210354703c105fbdf, /* 1797 */
128'he06f610560e200f70c630ff007930815, /* 1798 */
128'h0513bfe545018082610560e25535eb3f, /* 1799 */
128'hf0ef84aee822ec06e4261101bfcdf840, /* 1800 */
128'h0f840413e501cf0ff0ef842acd09f7df, /* 1801 */
128'hbfd555358082610564a2644260e2e080, /* 1802 */
128'hc3980015071b43887987879300004797, /* 1803 */
128'h780787930000479780820f8505138082, /* 1804 */
128'he8228e27879300005797110180824388, /* 1805 */
128'h644260e20094176384beec06e4266380, /* 1806 */
128'hf0ef8522c78119a447838082610564a2, /* 1807 */
128'he39c8b27879300005797b7d56000a9cf, /* 1808 */
128'h5797e50880827207ab2300004797e79c, /* 1809 */
128'he308e518e11ce788679889a787930000, /* 1810 */
128'he8a28824849300005497e4a6711d8082, /* 1811 */
128'he466e862ec5ef05af456f852fc4e6080, /* 1812 */
128'h060a0a1300004a1789aae0caec86e06a, /* 1813 */
128'h058b0b1300004b17050a8a9300004a97, /* 1814 */
128'h00003c9700050c1b058b8b9300004b97, /* 1815 */
128'h64a660e66446029415634d295ecc8c93, /* 1816 */
128'h6ca26c426be27b027aa27a4279e26906, /* 1817 */
128'hddcfe06f612511650513000045176d02, /* 1818 */
128'h89560007c36389524c1cc7914901541c, /* 1819 */
128'h0663dbefe0ef638c855a0fc42603681c, /* 1820 */
128'h00978e63601cdb2fe0ef855e85ca0009, /* 1821 */
128'h0000351701a98863da4fe0ef856685e2, /* 1822 */
128'he8221101b7716000286010ef57450513, /* 1823 */
128'hcfad44014d1cc1414401e04ae426ec06, /* 1824 */
128'hc7ad639cc7bd651ccbad511ccbbd4d5c, /* 1825 */
128'h842a15c010ef45051c00059384aa892e, /* 1826 */
128'h02a347850ef52c234799c57c57fdcd21, /* 1827 */
128'he65ff0ef0405282303253023e90410f5, /* 1828 */
128'h0000179716f43c2391c78793fffff797, /* 1829 */
128'h20a787930000179718f4302321a78793, /* 1830 */
128'h0247c78385220ea42e23681c18f43423, /* 1831 */
128'h64a2644260e28522e99ff0ef10f40023, /* 1832 */
128'h8693000046971180106f808261056902, /* 1833 */
128'h0017671302d786b365186294611c4966, /* 1834 */
128'h553b93ed836d8f3d0127d713e1189736, /* 1835 */
128'h808225018d5d00f717bb40f007b300f7, /* 1836 */
128'he4061141fc3ff06f6f85051300004517, /* 1837 */
128'h0105151bfe9ff0ef842afefff0efe022, /* 1838 */
128'he4061141808201412501640260a28d41, /* 1839 */
128'hfd1ff0ef14020005041bfdbff0efe022, /* 1840 */
128'h87aa80820141640260a28d4115029001, /* 1841 */
128'h8082fb75fee78fa30785fff5c7030585, /* 1842 */
128'h0785fff5c703058500c7896387aa962a, /* 1843 */
128'h86930007c70387aa8082fb65fee78fa3, /* 1844 */
128'hfee78fa30785fff5c7030585eb090017, /* 1845 */
128'h87b68082e21987aab7d587b68082fb75, /* 1846 */
128'hc6830585963efb7d001786930007c703, /* 1847 */
128'h15638082e291fed70fa300178713fff5, /* 1848 */
128'h47030585b7cd87ba8082000780a300c7, /* 1849 */
128'hd79b0187979b40f707bbfff5c7830005, /* 1850 */
128'h9463962e8082853ef37d0505e3994187, /* 1851 */
128'hfff5c783000547030585a839478100c5, /* 1852 */
128'h0505e3994187d79b0187979b40f707bb, /* 1853 */
128'h9363000547830ff5f5938082853eff79, /* 1854 */
128'hf59380824501bfcd0505c399808200b7, /* 1855 */
128'h0505dffd808200b79363000547830ff5, /* 1856 */
128'h808240a78533e7010007c70387aabfcd, /* 1857 */
128'hf0efec06842ae42ee8221101bfcd0785, /* 1858 */
128'h8663000547830ff5f593952265a2fe5f, /* 1859 */
128'h6105644260e24501fe857be3157d00b7, /* 1860 */
128'he7010007c70300b7856387aa95aa8082, /* 1861 */
128'hc68387aa862ab7fd0785808240a78533, /* 1862 */
128'h0705fed80fe38082ea9940c785330007, /* 1863 */
128'hbfcd872eb7d50785fe081be300074803, /* 1864 */
128'h8082ea1140d785330007c60387aa86aa, /* 1865 */
128'h8082fe081be300074803070500c80a63, /* 1866 */
128'h4501eb1900054703bff90785bfd5872e, /* 1867 */
128'h0505fafd0007c6830785fee68fe38082, /* 1868 */
128'h84aeec06e426e8221101bfd587aeb7e5, /* 1869 */
128'hcc1163804f47879300004797e519842a, /* 1870 */
128'hef8100044783942af9dff0ef85a68522, /* 1871 */
128'h644260e2852244014c07bc2300004797, /* 1872 */
128'hc519f9fff0ef852285a68082610564a2, /* 1873 */
128'h00004797050500050023c78100054783, /* 1874 */
128'he822ec066104e4261101bfd94aa7b623, /* 1875 */
128'h00050023c501f73ff0ef8526842ac891, /* 1876 */
128'h8082610564a28526644260e2e0080505, /* 1877 */
128'hce810007c68387aacf9900054783c11d, /* 1878 */
128'h00d780a300e780238082e3110017c703, /* 1879 */
128'h87aacb9d0075779380824501b7e50789, /* 1880 */
128'hff6d377d8fd507a2808204c79063963e, /* 1881 */
128'h0106ef6340e88833469d00c508b3872a, /* 1882 */
128'h963a97aa078e02e78733576100365793, /* 1883 */
128'hfef73c230721bfd10ff5f6934725bfc1, /* 1884 */
128'he7b300b50a63bf6dfeb78fa30785bfe1, /* 1885 */
128'h808202c79e63963e87aacb9d8b9d00a5, /* 1886 */
128'h40f88833ff07bc2307a1ff8738030721, /* 1887 */
128'h070e02f707b357e100365713ff06e8e3, /* 1888 */
128'h08b387aa872ebfc100e507b3963e95ba, /* 1889 */
128'h8fa30785fff5c7030585bfe1469d00c5, /* 1890 */
128'he432ec26852e842af0227179bf65fee7, /* 1891 */
128'hce1184aa6622dcdff0efe02ee84af406, /* 1892 */
128'h864a8522fff6091300c564636582892a, /* 1893 */
128'h8526740270a200040023f79ff0ef944a, /* 1894 */
128'h842ae406e02211418082614564e26942, /* 1895 */
128'h0141640260a28522f57ff0ef00a5e963, /* 1896 */
128'h00e587b340b6073300c506b395b28082, /* 1897 */
128'hb7fd00f6802316fd0005c78315fdd7e5, /* 1898 */
128'h000547838082853e478100c51563962a, /* 1899 */
128'h962ab7dd05850505fbed9f990005c703, /* 1900 */
128'h0505feb78de300054783808200c51363, /* 1901 */
128'hf406e44eec26852e842af0227179bfc5, /* 1902 */
128'h8522c8890005049bd1fff0ef89aee84a, /* 1903 */
128'h8522440100995b630005091bd13ff0ef, /* 1904 */
128'h86268082614569a2694264e2740270a2, /* 1905 */
128'hbfe90405d175f8bff0ef397d852285ce, /* 1906 */
128'h47038082450100c514630ff5f593962a, /* 1907 */
128'h47c1b7ed853efeb70be3001507930005, /* 1908 */
128'h4781e60187aa260100c7ef630ff5f593, /* 1909 */
128'h367d0785feb71ce30007c7038082853e, /* 1910 */
128'h069b40e7873b47a1c31d00757713b7f5, /* 1911 */
128'h078536fdfcb81ce30007c80387aa0007, /* 1912 */
128'h008597938e1d953e938102071793faf5, /* 1913 */
128'h5713020796938fd90107179300b7e733, /* 1914 */
128'hc703d24d8a1deb1187aa27018edd0036, /* 1915 */
128'h0007b803bfcd367d0785f8b71fe30007, /* 1916 */
128'hf8b712e30007c70300d80a6300878513, /* 1917 */
128'h419cb7f1377d87aabfa5fef51be30785, /* 1918 */
128'h470308f711630300079300054703e7a9, /* 1919 */
128'hc68300e786b3efe78793000027970015, /* 1920 */
128'h06930ff777130207071bc6898a850006, /* 1921 */
128'h0007c78397ba0025470304d71b630780, /* 1922 */
128'h1c6347c14198c19c47c1c3b10447f793, /* 1923 */
128'h478302f71663030007930005470302f7, /* 1924 */
128'h00074703973eeae70713000027170015, /* 1925 */
128'h078007130ff7f7930207879bc7098b05, /* 1926 */
128'hbf6d47a9bf7d47a18082050900e79363, /* 1927 */
128'hf63ff0efc632ec06006c842ee8221101, /* 1928 */
128'h4703e6a8081300002817468100c16583, /* 1929 */
128'h78930006460300f806330007079b0005, /* 1930 */
128'h61058536644260e2ec05000898630446, /* 1931 */
128'hf4e3fd07879b00088b63004678938082, /* 1932 */
128'hc6098a09b7d196be050502d586b3feb7, /* 1933 */
128'he008b7cdfc97879b0ff7f793fe07079b, /* 1934 */
128'h00063023f04afc06f426f8227139b7e1, /* 1935 */
128'h5529e90165a2b0dff0ef84b2842ae42e, /* 1936 */
128'h892a862e80826121790274a2744270e2, /* 1937 */
128'hc703fe8782e367e2f5dff0ef8522082c, /* 1938 */
128'h18e347a9fd279be307858f81cb010007, /* 1939 */
128'h02d0071300054683b7e94501e088fcf7, /* 1940 */
128'hf0efe40605051141f2dff06f00e68463, /* 1941 */
128'he02211418082014140a0053360a2f23f, /* 1942 */
128'hc70304b00693601cf0dff0ef842ee406, /* 1943 */
128'h0e630470069300e6ea6302d704630007, /* 1944 */
128'h076304d0069380820141640260a202d7, /* 1945 */
128'h07130017c683fed716e306b0069302d7, /* 1946 */
128'h042007130027c683fce69fe3052a0690, /* 1947 */
128'hbff1052a052ab7e9e01c078d00e69863, /* 1948 */
128'hc632ec06006c842ee8221101bfd50789, /* 1949 */
128'h081300002817468100c16583e0fff0ef, /* 1950 */
128'h460300f806330007079b00054703d168, /* 1951 */
128'h644260e2ec0500089863044678930006, /* 1952 */
128'h879b00088b6300467893808261058536, /* 1953 */
128'hb7d196be050502d586b3feb7f4e3fd07, /* 1954 */
128'hfc97879b0ff7f793fe07079bc6098a09, /* 1955 */
128'hf0ef842ee406e0221141b7e1e008b7cd, /* 1956 */
128'h02d704630007c70304b00693601cf87f, /* 1957 */
128'h640260a202d70e630470069300e6ea63, /* 1958 */
128'h06b0069302d7076304d0069380820141, /* 1959 */
128'h9fe3052a069007130017c683fed716e3, /* 1960 */
128'h078d00e69863042007130027c683fce6, /* 1961 */
128'h1141bfd50789bff1052a052ab7e9e01c, /* 1962 */
128'h00a405b395bff0efe589842ae406e022, /* 1963 */
128'hfff58513c3c7879300002797fff5c703, /* 1964 */
128'h557d640260a2e7198b1100074703973e, /* 1965 */
128'h973e00054703fea47ae3157d80820141, /* 1966 */
128'h4581462960a26402f77d8b1100074703, /* 1967 */
128'h1141fa5ff06f4581d7dff06f01410505, /* 1968 */
128'h014100e1550300a10723812100a107a3, /* 1969 */
128'h853ee3190005470345a9462547818082, /* 1970 */
128'h87bb00d667630ff6f693fd07069b8082, /* 1971 */
128'he0221141bff90505fd07879b9fb902f5, /* 1972 */
128'h45a900b7f86347a500a04563842ee406, /* 1973 */
128'h02a4753b4529fe7ff0ef357d02b455bb, /* 1974 */
128'h47854e60006f03050513014160a26402, /* 1975 */
128'h37230000471706f737230000471707fe, /* 1976 */
128'h0604041300004417e8221101808206f7, /* 1977 */
128'ha2fff0efec06600885aa84ae862ee426, /* 1978 */
128'h8082610564a26442e00c95a660e2600c, /* 1979 */
128'h000044970347879300004797e4261101, /* 1980 */
128'h35170004b9036380e04ae82202448493, /* 1981 */
128'hd0ef85a24124043bec065fa505130000, /* 1982 */
128'h862286aa608ce77fc0ef85a26088b9bf, /* 1983 */
128'h0000100fb81fd0ef5f05051300003517, /* 1984 */
128'h834a64a260e26442f14025730ff0000f, /* 1985 */
128'h83026105250106e58593000025976902, /* 1986 */
128'h008503638c0fa0ef8432e406e0221141, /* 1987 */
128'h71698082450180820141640260a2557d, /* 1988 */
128'hee26f606852289aae64e01258413f222, /* 1989 */
128'h852600a404b30505faeff0ef892eea4a, /* 1990 */
128'hfff5071beabff0ef95260505fa2ff0ef, /* 1991 */
128'hf6a7a0230000479704e7ee631ff00793, /* 1992 */
128'h380505130000351784aaf80ff0ef8522, /* 1993 */
128'h852204a7f2630ff007939526f72ff0ef, /* 1994 */
128'hf0ef3625051300003517842af62ff0ef, /* 1995 */
128'hd0ef542505130000351700a405b3f54f, /* 1996 */
128'h8082615569b2695264f2741270b2abbf, /* 1997 */
128'h0613b755f0f722230000471720000793, /* 1998 */
128'h859300003597893ff0ef850a45811000, /* 1999 */
128'h02f0079301294703e1aff0ef850a31e5, /* 2000 */
128'hf0ef850a514585930000359700f70963, /* 2001 */
128'h879300004797e22ff0ef850a85a2e2af, /* 2002 */
128'hd0ef4fa5051300003517858a4390ebe7, /* 2003 */
128'h332300004717451101f417934405a4bf, /* 2004 */
128'h4797db5ff0efeaf7332300004717eaf7, /* 2005 */
128'h00004797da7ff0ef4501c8a791230000, /* 2006 */
128'h854ec6a58593000045974611c6a79b23, /* 2007 */
128'h1101b799e687942300004797eb1ff0ef, /* 2008 */
128'h08c7df638432478de04ae426ec06e822, /* 2009 */
128'h25010004d783d69ff0ef84ae450d892a, /* 2010 */
128'hd53ff0efe38555030000451708a79563, /* 2011 */
128'h8513ffc4059b06a79a6325010024d783, /* 2012 */
128'h00004797d37ff0ef4511dc3ff0ef0044, /* 2013 */
128'hd23ff0efe085550300004517c0a79223, /* 2014 */
128'h859300004597bea79823000047974611, /* 2015 */
128'h4597256000ef4535e2dff0ef854abe65, /* 2016 */
128'h02000513d35ff0ef4515dde5d5830000, /* 2017 */
128'h0007d783dc87879300004797240000ef, /* 2018 */
128'h879300004797daf71d23000047172785, /* 2019 */
128'h0513000035170087cf63278d439cdae7, /* 2020 */
128'h6105690264a260e26442937fd0ef4065, /* 2021 */
128'h80826105690264a2644260e2d61ff06f, /* 2022 */
128'h00f10fa347090105c783f022f4067179, /* 2023 */
128'h00e78e6301e1578300f10f230115c783, /* 2024 */
128'h05130000351770a2740202e78a63470d, /* 2025 */
128'h051300003517842a8e5fd06f61453e65, /* 2026 */
128'h70a265a2740285228d5fd0efe42e3be5, /* 2027 */
128'h614505c170a241907402d8dff06f6145, /* 2028 */
128'h2291342322813823dc010113ebfff06f, /* 2029 */
128'h218006134581893284ae842a23213023, /* 2030 */
128'h2040061385a6e92ff0ef22113c230028, /* 2031 */
128'hf0ef8522002ced4ff0efe802c44a0828, /* 2032 */
128'h3903228134832301340323813083f63f, /* 2033 */
128'hcc47d783000047978082240101132201, /* 2034 */
128'hcf5ff06faac58593000045974611cb81, /* 2035 */
128'h878e1041e703492000efe40611418082, /* 2036 */
128'ha22310e1a02327051001a70300e57763, /* 2037 */
128'h8d5d91011782150260a21007e78310a7, /* 2038 */
128'he426e822ec0611018082450180820141, /* 2039 */
128'h3e8007933ce000ef842afc1ff0ef84aa, /* 2040 */
128'h02a7d533644260e29101150202f407b3, /* 2041 */
128'hf0efe022e40611418082610564a28d05, /* 2042 */
128'h24078793000f47b73a2000ef842af95f, /* 2043 */
128'hd533014191011502640260a202f407b3, /* 2044 */
128'h84aae04ae426e822ec061101808202a7, /* 2045 */
128'h443702a48533370000ef892af63ff0ef, /* 2046 */
128'hf0ef0405944a0285543324040413000f, /* 2047 */
128'h6105690264a2644260e2fe856ee3f45f, /* 2048 */
128'he04aec06e822009894b7e42611018082, /* 2049 */
128'h854a89260084f363892268048493842a, /* 2050 */
128'h64a2644260e2f47dfa1ff0ef41240433, /* 2051 */
128'h00054503808200b50023808261056902, /* 2052 */
128'h8082020575130147c503100007b78082, /* 2053 */
128'h0023dfe50207f7930147478310000737, /* 2054 */
128'hf800071300078223100007b7808200a7, /* 2055 */
128'h470d0007822300e78023476d00e78623, /* 2056 */
128'h0200071300e78423fc70071300e78623, /* 2057 */
128'h4503842ae406e0221141808200e78823, /* 2058 */
128'hfa5ff0ef80820141640260a2e5090004, /* 2059 */
128'h00f57713b947879300002797b7f50405, /* 2060 */
128'h80a30007c7830007470397aa973e8111, /* 2061 */
128'h842a002ce8221101808200f5802300e5, /* 2062 */
128'hf65ff0ef00814503fd1ff0efec068121, /* 2063 */
128'hf0ef0ff47513002cf5dff0ef00914503, /* 2064 */
128'hf0ef00914503f4bff0ef00814503fb7f, /* 2065 */
128'hec26f022717980826105644260e2f43f, /* 2066 */
128'h002c0089553b54e14461892af406e84a, /* 2067 */
128'hf0ef346100814503f81ff0ef0ff57513, /* 2068 */
128'h70a2fe9410e3f0bff0ef00914503f13f, /* 2069 */
128'hec26f022717980826145694264e27402, /* 2070 */
128'h0089553354e103800413892af406e84a, /* 2071 */
128'h346100814503f3fff0ef0ff57513002c, /* 2072 */
128'hfe9410e3ec9ff0ef00914503ed1ff0ef, /* 2073 */
128'h002c110180826145694264e2740270a2, /* 2074 */
128'h4503ea7ff0ef00814503f13ff0efec06, /* 2075 */
128'h0000100f8082610560e2e9fff0ef0091, /* 2076 */
128'h8593000025974305f14025730ff0000f, /* 2077 */
128'h000035974605d90101138302037eab65, /* 2078 */
128'h26113423a145051300004517e2c58593, /* 2079 */
128'h253134232521382324913c2326813023, /* 2080 */
128'h00003517c5152501e75fa0ef25413023, /* 2081 */
128'h2601340326813083d64fd0ef08450513, /* 2082 */
128'h24013a03248139832501390325813483, /* 2083 */
128'hd0ef07a5051300003517808227010113, /* 2084 */
128'ha0ef080808c58593000035974605d3af, /* 2085 */
128'h3a1709620bf00913e12d44812501e85f, /* 2086 */
128'h6605007491810204959314aa0a130000, /* 2087 */
128'h00c4d41be5052501fedfa0ef080895ca, /* 2088 */
128'h45039452dc9ff0ef880d45210004099b, /* 2089 */
128'h9cbd47b2286010ef854edbfff0ef0004, /* 2090 */
128'h3517c9192501c96fb0ef54020808f3f9, /* 2091 */
128'h0285051300003517bfb904a505130000, /* 2092 */
128'ha0ef4501d4458593000035974605bf91, /* 2093 */
128'hbf1d03a5051300003517c5112501dabf, /* 2094 */
128'h0000351785a20184961386a20bf00493, /* 2095 */
128'h0785051300003517c84fd0ef03c50513, /* 2096 */
128'h059b962f90ef0184951385a2c78fd0ef, /* 2097 */
128'hd0ef0725051300003517c981c62e0005, /* 2098 */
128'hc4cfd0ef8445051300003517bdddc5af, /* 2099 */
128'he40625011141900200000023e8dff0ef, /* 2100 */
128'h808224050513000f4537a001ddbff0ef, /* 2101 */
128'h157d631c89c707130000471780824501, /* 2102 */
128'h10d00513e30895360017869300756513, /* 2103 */
128'hec06e822110102b506338082953e055e, /* 2104 */
128'h45816622c509842afd1ff0efe4328532, /* 2105 */
128'h808280826105644260e285229e8ff0ef, /* 2106 */
128'hbccfd0efe40600e50513000035171141, /* 2107 */
128'h80820141450160a2f89fc0ef20000537, /* 2108 */
128'h553347a9b00025738082450180824501, /* 2109 */
128'h351785aa862e86b287361141808202f5, /* 2110 */
128'hf0ef4505b90fd0efe406ffa505130000, /* 2111 */
128'hf0efe406952e842ae0221141a001d2df, /* 2112 */
128'h01418d7d640260a29522408007b3f57f, /* 2113 */
128'h71798082450580824505808245058082, /* 2114 */
128'h0096186300c684bb842ef406ec26f022, /* 2115 */
128'h852285b280826145450164e2740270a2, /* 2116 */
128'hbff92605200404136622edbfc0efe432, /* 2117 */
128'h80828082808245098082450980824509, /* 2118 */
128'h1101c2dff06f80824501808245018082, /* 2119 */
128'h00d584b3003796934781e426e822ec06, /* 2120 */
128'h450164a2644260e200c7986300d50433, /* 2121 */
128'h600c02e8036360980004380380826105, /* 2122 */
128'h8626acefd0eff6e50513000035176090, /* 2123 */
128'ha001abefd0eff86505130000351785a2, /* 2124 */
128'h051300003517892ae0ca711dbf5d0785, /* 2125 */
128'he862ec5ef05af456f852fc4ee8a2f865, /* 2126 */
128'h3a17a8efd0ef44018b2ee466e4a6ec86, /* 2127 */
128'h4993f7ab8b9300003b97f72a0a130000, /* 2128 */
128'hd0ef85524ac1f7ec0c1300003c17fff9, /* 2129 */
128'h87caa5efd0ef855e85e600040c9ba6af, /* 2130 */
128'h856285e6a50fd0ef8552036498634481, /* 2131 */
128'h17e3040502b49b63458187caa48fd0ef, /* 2132 */
128'h4501a2efd0effa65051300003517fd54, /* 2133 */
128'h00349713c689873e8a85008486b3a889, /* 2134 */
128'h86b3bf5d07a104856398e39840e98733, /* 2135 */
128'h873300359713c689873e8a8563900085, /* 2136 */
128'hf085051300003517058e02e60d6340e9, /* 2137 */
128'h9dcfd0eff3450513000035179e8fd0ef, /* 2138 */
128'h7aa27a4279e2690664a6644660e6557d, /* 2139 */
128'h07a10585808261256ca26c426be27b02, /* 2140 */
128'h020005138aaa6a05fc56e0d27159bfa5, /* 2141 */
128'he8caf0a2f486f062f45ef85ae4ceeca6, /* 2142 */
128'hbb1ff0ef44818bb28b2ee46ee86aec66, /* 2143 */
128'h9793252c0c1300003c179c4a0a134981, /* 2144 */
128'h351703749b6300fb0cb300fa8db30034, /* 2145 */
128'h694670a67406962fd0eff02505130000, /* 2146 */
128'h86266da26d426ce27c027ba26a0669a6, /* 2147 */
128'he33ff06f61657ae285567b4264e685da, /* 2148 */
128'hc75fe0ef8d2ac7bfe0ef842ac81fe0ef, /* 2149 */
128'h1d1b0105151b0344f7b3c6ffe0ef892a, /* 2150 */
128'h91011402150201a4643300a96533010d, /* 2151 */
128'hf0ef4521ef8100adb02300acb0238d41, /* 2152 */
128'hf0ef0007c50397e20039f7930985b1ff, /* 2153 */
128'hf822fc06e032e42e7139b7ad0485b0ff, /* 2154 */
128'he0ef842ac19fe0ef89aaec4ef04af426, /* 2155 */
128'h151bc07fe0ef84aac0dfe0ef892ac13f, /* 2156 */
128'h65a2660215028fc18d450109179b0105, /* 2157 */
128'h00e588330037971347818d5d91011782, /* 2158 */
128'h854e790274a270e2744200c79c63974e, /* 2159 */
128'h8ea907856314d79ff06f6121863e69e2, /* 2160 */
128'h7139b7f100e830238f2900083703e314, /* 2161 */
128'h89aaec4ef04af426f822fc06e032e42e, /* 2162 */
128'hb95fe0ef892ab9bfe0ef842aba1fe0ef, /* 2163 */
128'h8d450109179b0105151bb8ffe0ef84aa, /* 2164 */
128'h47818d5d9101178265a2660215028fc1, /* 2165 */
128'h744200c79c63974e00e5883300379713, /* 2166 */
128'hf06f6121863e69e2854e790274a270e2, /* 2167 */
128'h8f0900083703e3148e8907856314d01f, /* 2168 */
128'hf822fc06e032e42e7139b7f100e83023, /* 2169 */
128'he0ef842ab29fe0ef89aaec4ef04af426, /* 2170 */
128'h151bb17fe0ef84aab1dfe0ef892ab23f, /* 2171 */
128'h65a2660215028fc18d450109179b0105, /* 2172 */
128'h00e588330037971347818d5d91011782, /* 2173 */
128'h854e790274a270e2744200c79c63974e, /* 2174 */
128'h86b307856314c89ff06f6121863e69e2, /* 2175 */
128'h00e8302302a7073300083703e31402a6, /* 2176 */
128'hf04af426f822fc06e032e42e7139b7e1, /* 2177 */
128'h892aaa7fe0ef842aaadfe0ef89aaec4e, /* 2178 */
128'h179b0105151ba9bfe0ef84aaaa1fe0ef, /* 2179 */
128'h9101178265a2660215028fc18d450109, /* 2180 */
128'h9c63974e00e588330037971347818d5d, /* 2181 */
128'h863e69e2854e790274a270e2744200c7, /* 2182 */
128'hd6b3078563144505e111c0dff06f6121, /* 2183 */
128'h00e8302302a7573300083703e31402a6, /* 2184 */
128'hf04af426f822fc06e032e42e7139b7d1, /* 2185 */
128'h892aa27fe0ef842aa2dfe0ef89aaec4e, /* 2186 */
128'h179b0105151ba1bfe0ef84aaa21fe0ef, /* 2187 */
128'h9101178265a2660215028fc18d450109, /* 2188 */
128'h9c63974e00e588330037971347818d5d, /* 2189 */
128'h863e69e2854e790274a270e2744200c7, /* 2190 */
128'h3703e3148ec907856314b8dff06f6121, /* 2191 */
128'he032e42e7139b7f100e830238f490008, /* 2192 */
128'h9b5fe0ef89aaec4ef04af426f822fc06, /* 2193 */
128'he0ef84aa9a9fe0ef892a9affe0ef842a, /* 2194 */
128'h15028fc18d450109179b0105151b9a3f, /* 2195 */
128'h0037971347818d5d9101178265a26602, /* 2196 */
128'h74a270e2744200c79c63974e00e58833, /* 2197 */
128'h6314b15ff06f6121863e69e2854e7902, /* 2198 */
128'h00e830238f6900083703e3148ee90785, /* 2199 */
128'hf04af426f822fc06e032e42e7139b7f1, /* 2200 */
128'h892a937fe0ef842a93dfe0ef89aaec4e, /* 2201 */
128'h179b0105151b92bfe0ef84aa931fe0ef, /* 2202 */
128'h9081178265a2660214828fc18cc90109, /* 2203 */
128'h1c6396ae00d988330037169347018fc5, /* 2204 */
128'h863a69e2854e790274a270e2744200c7, /* 2205 */
128'h00a83023e28800f70533a9dff06f6121, /* 2206 */
128'h051300003517892ae8ca7159bfc90705, /* 2207 */
128'hf062f45ef85afc56e0d2e4cef0a2a665, /* 2208 */
128'hd6dfc0ef44018b3289aeec66eca6f486, /* 2209 */
128'ha58b8b9300003b97a50a0a1300003a17, /* 2210 */
128'hc0ef855204000a93a60c0c1300003c17, /* 2211 */
128'hd3dfc0ef8885855e85a2fff44493d4bf, /* 2212 */
128'h00f905b30036179314fd460140900cb3, /* 2213 */
128'h85a2d1ffc0efe43285520566186397ce, /* 2214 */
128'ha03ff0ef854a85ce6622d17fc0ef8562, /* 2215 */
128'h051300003517fb541be32405e12984aa, /* 2216 */
128'h64e669468526740670a6cf7fc0efa6e5, /* 2217 */
128'h61656ce27c027ba27b427ae26a0669a6, /* 2218 */
128'he198e3988726c2918766001676938082, /* 2219 */
128'h351784aaeca67159bfc154fdbf590605, /* 2220 */
128'hfc56e0d2e4cee8caf0a2992505130000, /* 2221 */
128'h8ab2892ee86af486ec66f062f45ef85a, /* 2222 */
128'h3b1797a9899300003997c97fc0ef4401, /* 2223 */
128'h3c17c3ab8b9300003b97c3ab0b130000, /* 2224 */
128'h0a1397ac8c9300003c97972c0c130000, /* 2225 */
128'hbd03cba500147793c65fc0ef854e0400, /* 2226 */
128'hfffd45134601c53fc0ef856285a2000b, /* 2227 */
128'h854e05561c6397ca00f485b300361793, /* 2228 */
128'h6622c2ffc0ef856685a2c37fc0efe432, /* 2229 */
128'h1ae32405e5298d2a91bff0ef852685ca, /* 2230 */
128'h70a6c0ffc0ef9865051300003517fb44, /* 2231 */
128'h7b427ae26a0669a6694664e6856a7406, /* 2232 */
128'h000b3d03808261656d426ce27c027ba2, /* 2233 */
128'he198e398872ac291876a00167693bf49, /* 2234 */
128'h3517842ae8a2711db7e15d7db7790605, /* 2235 */
128'hf05af456f852e0cae4a68a2505130000, /* 2236 */
128'hc0ef4c018ab284aefc4eec86e862ec5e, /* 2237 */
128'h0b1300003b1788e9091300003917babf, /* 2238 */
128'h854a10000a1389eb8b9300003b97896b, /* 2239 */
128'hb7dfc0ef855a85ce000c099bb89fc0ef, /* 2240 */
128'h17130187e7b38fd9010c1793008c1713, /* 2241 */
128'h8fd9028c17138fd9020c17138fd9018c, /* 2242 */
128'h171346018fd9038c17138fd9030c1713, /* 2243 */
128'he432854a05561763972600e406b30036, /* 2244 */
128'h85a66622b31fc0ef855e85ceb39fc0ef, /* 2245 */
128'hf94c19e30c05e91d89aa81dff0ef8522, /* 2246 */
128'h644660e6b11fc0ef8885051300003517, /* 2247 */
128'h6be27b027aa27a4279e2690664a6854e, /* 2248 */
128'h59fdb74d0605e29ce31c808261256c42, /* 2249 */
128'h7b8505130000251784aaf4a67119bff1, /* 2250 */
128'hf862fc5ee0dae4d6e8d2eccef0caf8a2, /* 2251 */
128'hc0ef44018b32892eec6efc86f06af466, /* 2252 */
128'h8c9300002c9779ea0a1300002a17abbf, /* 2253 */
128'h00002d1703f00c13498507f00b937a6c, /* 2254 */
128'h85a2a8ffc0ef855208000a937a4d0d13, /* 2255 */
128'h95b300e99733408b873ba87fc0ef8566, /* 2256 */
128'h1a6397ca00f486b30036179346010089, /* 2257 */
128'hc0ef856a85a2a63fc0efe43285520566, /* 2258 */
128'he1398daaf46ff0ef852685ca6622a5bf, /* 2259 */
128'hc0ef7b25051300002517fb541be32405, /* 2260 */
128'h6a4669e6790674a6856e744670e6a3bf, /* 2261 */
128'h61096de27d027ca27c427be26b066aa6, /* 2262 */
128'he398bf610605e28ce38c008c66638082, /* 2263 */
128'h251784aaf4a67119b7f15dfdbfe5e298, /* 2264 */
128'he4d6e8d2eccef0caf8a26d2505130000, /* 2265 */
128'h892eec6efc86f06af466f862fc5ee0da, /* 2266 */
128'h6b8a0a1300002a179d5fc0ef44018b32, /* 2267 */
128'h0c13498507f00b936c0c8c9300002c97, /* 2268 */
128'h855208000a936bed0d1300002d1703f0, /* 2269 */
128'h408b87bb9a1fc0ef856685a29a9fc0ef, /* 2270 */
128'hfff6c693fff7c793008996b300f997b3, /* 2271 */
128'h05661a63974a00e485b3003617134601, /* 2272 */
128'h96dfc0ef856a85a2975fc0efe4328552, /* 2273 */
128'h2405e1398daae58ff0ef852685ca6622, /* 2274 */
128'h94dfc0ef6c45051300002517fb5417e3, /* 2275 */
128'h6aa66a4669e6790674a6856e744670e6, /* 2276 */
128'h808261096de27d027ca27c427be26b06, /* 2277 */
128'he19ce31cbf610605e194e314008c6663, /* 2278 */
128'h0000251784aaf4a67119b7f15dfdbfe5, /* 2279 */
128'he0dae4d6e8d2eccef0caf8a25e450513, /* 2280 */
128'h8a32892eec6efc86f06af466f862fc5e, /* 2281 */
128'h2c175ca98993000029978e7fc0ef4401, /* 2282 */
128'h08100b134d0507f00a935d2c0c130000, /* 2283 */
128'hc0ef854e5ccc8c9300002c9703f00b93, /* 2284 */
128'h07bb408a873b8b3fc0ef856285a28bbf, /* 2285 */
128'h0024079b8f5d00ed173300fd17b3408b, /* 2286 */
128'hc313fff748938fd5008d16b300fd17b3, /* 2287 */
128'h1c6396ca00d48533003616934601fff7, /* 2288 */
128'hc0ef856685a2873fc0efe432854e0546, /* 2289 */
128'hed298daad56ff0ef852685ca662286bf, /* 2290 */
128'h051300002517f8f41be3080007932405, /* 2291 */
128'h790674a6856e744670e6847fc0ef5be5, /* 2292 */
128'h7d027ca27c427be26b066aa66a4669e6, /* 2293 */
128'h859a008bea6300167813808261096de2, /* 2294 */
128'h85c6b7610605e10ce28c85be00081363, /* 2295 */
128'hf0ca7119bf755dfdbfc585bafe081be3, /* 2296 */
128'hfc5ee8d2ecce4ce5051300002517892a, /* 2297 */
128'he0dae4d6f4a6f8a2fc86ec6ef06af466, /* 2298 */
128'h00002a17fd0fc0ef4b81e03289aef862, /* 2299 */
128'h00002d174bcc8c9300002c974b4a0a13, /* 2300 */
128'h003b949b01779c3347854da14c4d0d13, /* 2301 */
128'h856685da00848b3bfa4fc0ef85524401, /* 2302 */
128'h0036171367824601fffc4a93f98fc0ef, /* 2303 */
128'hc0efe432855206f61063974e00e90833, /* 2304 */
128'h854a85ce6622f72fc0ef856a85daf7af, /* 2305 */
128'hfbb41be38c562405e9318b2ac5eff0ef, /* 2306 */
128'h051300002517fafb90e3040007932b85, /* 2307 */
128'h790674a6855a744670e6f46fc0ef4be5, /* 2308 */
128'h7d027ca27c427be26b066aa66a4669e6, /* 2309 */
128'h85d6e11185e200167513808261096de2, /* 2310 */
128'h7175b7e95b7db749060500b83023e30c, /* 2311 */
128'h698502000513892e84aaf4cef8cafca6, /* 2312 */
128'he122e506fc66e0e2e4dee8daecd6f0d2, /* 2313 */
128'h3c174a01904ff0ef4a81e032f46ef86a, /* 2314 */
128'h8c9300002c979c498993daac0c130000, /* 2315 */
128'h003d969367824d214d818bca8b2679ec, /* 2316 */
128'hba2ff0ef852685ca866e04fd956396da, /* 2317 */
128'h4385051300002517020a0863ed45842a, /* 2318 */
128'h79a6794674e6640a60aa8522e98fc0ef, /* 2319 */
128'h7da27d427ce26c066ba66b466ae67a06, /* 2320 */
128'he0efec36b7758ba68b4a4a0580826149, /* 2321 */
128'he42a9a6fe0efe82a9acfe0ef842a9b2f, /* 2322 */
128'h161b8d5d0105151b664267a29a0fe0ef, /* 2323 */
128'h37978d4166e29101140215028c510106, /* 2324 */
128'hc683018786b34781e288d0a7b5230000, /* 2325 */
128'h00d600230ff6f693078500fb86330006, /* 2326 */
128'hf0ef4521ef910ba1033df7b3ffa795e3, /* 2327 */
128'hc50397e68b8d00078a9b001a879b82ef, /* 2328 */
128'h7175bfa1547dbf0d0d8581aff0ef0007, /* 2329 */
128'h6a050200051389ae892af0d2f4cef8ca, /* 2330 */
128'he506f86afc66e0e2e4dee8daecd6fca6, /* 2331 */
128'h34974a81fe5fe0ef4b018cb2f46ee122, /* 2332 */
128'h0d1300002d179c4a0a13c92484930000, /* 2333 */
128'h00fc06b3003d97934d818c4e8bca67ed, /* 2334 */
128'ha82ff0ef854a85ce866e059d956397de, /* 2335 */
128'h3185051300002517020a8863e579842a, /* 2336 */
128'h79a6794674e6640a60aa8522d78fc0ef, /* 2337 */
128'h7da27d427ce26c066ba66b466ae67a06, /* 2338 */
128'he836ec3eb7758c4a8bce4a8580826149, /* 2339 */
128'h884fe0efe42a88afe0ef842a890fe0ef, /* 2340 */
128'h161b0105151b6702662287efe0efe02a, /* 2341 */
128'h37978d419101140215028c518d590106, /* 2342 */
128'h0004d783e38866c267e2bea7b9230000, /* 2343 */
128'h93c117c20024d78300f6902393c117c2, /* 2344 */
128'h00f6922393c117c20044d78300f69123, /* 2345 */
128'h034df7b300f6932393c117c20064d783, /* 2346 */
128'h00078b1b001b079bef9fe0ef4521ef91, /* 2347 */
128'hbf290d85ee5fe0ef0007c50397ea8b8d, /* 2348 */
128'h86138932f8ca717580826505b789547d, /* 2349 */
128'h251785aa962a84ae842afca6e122fff5, /* 2350 */
128'he4dee8daecd6f0d2f4ce23a505130000, /* 2351 */
128'hc7cfc0efec36e506f46ef86afc66e0e2, /* 2352 */
128'h99a20034d793e83e0014d9930044d793, /* 2353 */
128'h2b97222b0b1300002b1744854a81e43e, /* 2354 */
128'h2c97222c0c1300002c17222b8b930000, /* 2355 */
128'h2d9722ad0d1300002d17222c8c930000, /* 2356 */
128'h7863aeaa0a1300003a1722ad8d930000, /* 2357 */
128'h60aac1efc0ef21e50513000025170299, /* 2358 */
128'h6b466ae67a0679a6794674e68556640a, /* 2359 */
128'h85a6808261497da27d427ce26c066ba6, /* 2360 */
128'hc0ef855e85ca00090663bf6fc0ef855a, /* 2361 */
128'hbdcfc0ef856a85e6be4fc0ef8562beaf, /* 2362 */
128'hbccfc0ef856eed15920ff0ef852265a2, /* 2363 */
128'hc58d000a358302f749636762010a2783, /* 2364 */
128'h008a3783bb0fc0ef1a05051300002517, /* 2365 */
128'h19050513000025179782852285ce6642, /* 2366 */
128'hec05051300002517b7e94a89b98fc0ef, /* 2367 */
128'h0513000025177179bfa10485b88fc0ef, /* 2368 */
128'hc8bfe0efe44ee84aec26f022f40617e5, /* 2369 */
128'hb5cfc0ef17c505130000251704000593, /* 2370 */
128'h00002517b50fc0ef1985051300002517, /* 2371 */
128'he705051300002517b44fc0ef1bc50513, /* 2372 */
128'h95b3497901f499934441b36fc0ef4485, /* 2373 */
128'he6dff0ef240501358533460546850084, /* 2374 */
128'h614569a2694264e2740270a2ff2417e3, /* 2375 */
128'h46814881470100c5131b460580828082, /* 2376 */
128'h000780234000081387f245a901f61e13, /* 2377 */
128'h802397aa0007802397aa0007802397aa, /* 2378 */
128'h02b71d632705fe0813e397aa387d0007, /* 2379 */
128'h86b33e800513c00026f38e15c0202673, /* 2380 */
128'h45bb02c747334000059302a687334116, /* 2381 */
128'h05130000251702a7473302a767b302b3, /* 2382 */
128'h28f3c02026f3fac710e3a96fc06f1565, /* 2383 */
128'h4505f7bff0ef4501e4061141bf51c000, /* 2384 */
128'hf69ff0ef4511f6fff0ef4509f75ff0ef, /* 2385 */
128'h07b7bff1f5dff0ef4541f63ff0ef4521, /* 2386 */
128'h07b780824788400007b78082c3884000, /* 2387 */
128'h05130000251780824b880007a8234000, /* 2388 */
128'hec4ef04af426fc067139b55fe06f1be5, /* 2389 */
128'h00002517b0dfe0eff822e05ae456e852, /* 2390 */
128'h0b1300002b174901b33fe0ef11c50513, /* 2391 */
128'h2a17112a8a9300002a97400004b72e6b, /* 2392 */
128'h0007c783016907b34991122a0a130000, /* 2393 */
128'hc0ef862224014480448cc09c09058556, /* 2394 */
128'h1de39cefc0ef8552488c0004a8239daf, /* 2395 */
128'h02e78b634709006457930ff47413fd39, /* 2396 */
128'h0000251700e78c63470504e78163470d, /* 2397 */
128'ha001bfdfe0ef85229a4fc0ef0ec50513, /* 2398 */
128'he0dff0ef990fc0ef0e85051300002517, /* 2399 */
128'h80ef97efc0ef0e65051300002517b7fd, /* 2400 */
128'h96cfc0ef0e45051300002517bff1f7af, /* 2401 */
128'h00000000000000000000b7e9ee5ff0ef, /* 2402 */
128'h00000000000000000000000000000000, /* 2403 */
128'h00000000000000000000000000000000, /* 2404 */
128'h00000000000000000000000000000000, /* 2405 */
128'h00000000000000000000000000000000, /* 2406 */
128'h00000000000000000000000000000000, /* 2407 */
128'h00000000000000000000000000000000, /* 2408 */
128'h00000000000000000000000000000000, /* 2409 */
128'h00000000000000000000000000000000, /* 2410 */
128'h00000000000000000000000000000000, /* 2411 */
128'h00000000000000000000000000000000, /* 2412 */
128'h00000000000000000000000000000000, /* 2413 */
128'h00000000000000000000000000000000, /* 2414 */
128'h00000000000000000000000000000000, /* 2415 */
128'h08082828282828080808080808080808, /* 2416 */
128'h08080808080808080808080808080808, /* 2417 */
128'h101010101010101010101010101010a0, /* 2418 */
128'h10101010101004040404040404040404, /* 2419 */
128'h01010101010101010141414141414110, /* 2420 */
128'h10101010100101010101010101010101, /* 2421 */
128'h02020202020202020242424242424210, /* 2422 */
128'h08101010100202020202020202020202, /* 2423 */
128'h00000000000000000000000000000000, /* 2424 */
128'h00000000000000000000000000000000, /* 2425 */
128'h101010101010101010101010101010a0, /* 2426 */
128'h10101010101010101010101010101010, /* 2427 */
128'h01010101010101010101010101010101, /* 2428 */
128'h02010101010101011001010101010101, /* 2429 */
128'h02020202020202020202020202020202, /* 2430 */
128'h02020202020202021002020202020202, /* 2431 */
128'hc1bdceee242070dbe8c7b756d76aa478, /* 2432 */
128'hfd469501a83046134787c62af57c0faf, /* 2433 */
128'h895cd7beffff5bb18b44f7af698098d8, /* 2434 */
128'h49b40821a679438efd9871936b901122, /* 2435 */
128'he9b6c7aa265e5a51c040b340f61e2562, /* 2436 */
128'he7d3fbc8d8a1e68102441453d62f105d, /* 2437 */
128'h455a14edf4d50d87c33707d621e1cde6, /* 2438 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /* 2439 */
128'hfde5380c6d9d61228771f681fffa3942, /* 2440 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /* 2441 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /* 2442 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /* 2443 */
128'hfc93a039ab9423a7432aff97f4292244, /* 2444 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /* 2445 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /* 2446 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /* 2447 */
128'h0c07020d08030e09040f0a05000b0601, /* 2448 */
128'h020f0c090603000d0a0704010e0b0805, /* 2449 */
128'h09020b040d060f08010a030c050e0700, /* 2450 */
128'h6c5f7465735f64735f63736972776f6c, /* 2451 */
128'h6e67696c615f64730000000000006465, /* 2452 */
128'h645f6b6c635f64730000000000000000, /* 2453 */
128'h69747465735f64730000000000007669, /* 2454 */
128'h735f646d635f6473000000000000676e, /* 2455 */
128'h74657365725f64730000000074726174, /* 2456 */
128'h6e636b6c625f64730000000000000000, /* 2457 */
128'h69736b6c625f64730000000000000074, /* 2458 */
128'h6f656d69745f6473000000000000657a, /* 2459 */
128'h655f7172695f64730000000000007475, /* 2460 */
128'h5f63736972776f6c000000000000006e, /* 2461 */
128'h00000000646d635f74726174735f6473, /* 2462 */
128'h746e695f746961775f63736972776f6c, /* 2463 */
128'h000000000067616c665f747075727265, /* 2464 */
128'h00007172695f64735f63736972776f6c, /* 2465 */
128'h695f646d635f64735f63736972776f6c, /* 2466 */
128'h5f63736972776f6c0000000000007172, /* 2467 */
128'h007172695f646e655f617461645f6473, /* 2468 */
128'h00000000bffe9a8800000000bffead70, /* 2469 */
128'h004c4b40004c4b400030000020000000, /* 2470 */
128'h6d6d5f6472616f62000000020000ffff, /* 2471 */
128'h00000000bffe4e8c0064637465675f63, /* 2472 */
128'h00000000bffe4cf800000000bffe4a9a, /* 2473 */
128'h00000000000000000000000000000000, /* 2474 */
128'hffffbd6effffbd6affffbd6affffbd44, /* 2475 */
128'hffffbd72ffffbd72ffffbd72ffffbd72, /* 2476 */
128'h00000000bffeb09800000000bffeb088, /* 2477 */
128'h00000000bffeb0c000000000bffeb0a8, /* 2478 */
128'h00000000bffeb0f000000000bffeb0d8, /* 2479 */
128'h00000000bffeb12000000000bffeb108, /* 2480 */
128'h00000000bffeb15000000000bffeb138, /* 2481 */
128'h00000000bffeb18000000000bffeb168, /* 2482 */
128'h40040300400402004004010040040000, /* 2483 */
128'h40050000400405004004040140040400, /* 2484 */
128'h30000000000000030000000040050100, /* 2485 */
128'h60000000000000053000000000000001, /* 2486 */
128'h70000000000000027000000000000004, /* 2487 */
128'h00000001400000007000000000000000, /* 2488 */
128'h00000005000000012000000000000006, /* 2489 */
128'h20000000000000020000000040000000, /* 2490 */
128'h00000000100000000000000100000000, /* 2491 */
128'h1e19140f0d0c0a000000000000000000, /* 2492 */
128'h000186a00000271050463c37322d2823, /* 2493 */
128'h017d7840017d784000989680000f4240, /* 2494 */
128'h031975000319750002faf080018cba80, /* 2495 */
128'h02faf08005f5e10002faf080017d7840, /* 2496 */
128'h00000020000000000bebc2000c65d400, /* 2497 */
128'h00000200000001000000008000000040, /* 2498 */
128'h00002000000010000000080000000400, /* 2499 */
128'h0000c000000080000000600000004000, /* 2500 */
128'h37363534333231300002000000010000, /* 2501 */
128'h2043534952776f4c4645444342413938, /* 2502 */
128'h746f6f622d7520646573696d696e696d, /* 2503 */
128'h00000000647261432d445320726f6620, /* 2504 */
128'he00600003800000039080000edfe0dd0, /* 2505 */
128'h00000000100000001100000028000000, /* 2506 */
128'h0000000000000000a806000059010000, /* 2507 */
128'h00000000010000000000000000000000, /* 2508 */
128'h02000000000000000400000003000000, /* 2509 */
128'h020000000f0000000400000003000000, /* 2510 */
128'h2c6874651b0000001400000003000000, /* 2511 */
128'h007665642d657261622d656e61697261, /* 2512 */
128'h2c687465260000001000000003000000, /* 2513 */
128'h0100000000657261622d656e61697261, /* 2514 */
128'h1a0000000300000000006e65736f6863, /* 2515 */
128'h303140747261752f636f732f2c000000, /* 2516 */
128'h0000003030323531313a303030303030, /* 2517 */
128'h00000000737570630100000002000000, /* 2518 */
128'h01000000000000000400000003000000, /* 2519 */
128'h000000000f0000000400000003000000, /* 2520 */
128'h40787d01380000000400000003000000, /* 2521 */
128'h03000000000000304075706301000000, /* 2522 */
128'h0300000080f0fa024b00000004000000, /* 2523 */
128'h03000000007570635b00000004000000, /* 2524 */
128'h03000000000000006700000004000000, /* 2525 */
128'h0000000079616b6f6b00000005000000, /* 2526 */
128'h7a6874651b0000001300000003000000, /* 2527 */
128'h0000766373697200656e61697261202c, /* 2528 */
128'h34367672720000000b00000003000000, /* 2529 */
128'h0b000000030000000000636466616d69, /* 2530 */
128'h0000393376732c76637369727c000000, /* 2531 */
128'h01000000850000000000000003000000, /* 2532 */
128'h6f72746e6f632d747075727265746e69, /* 2533 */
128'h04000000030000000000000072656c6c, /* 2534 */
128'h0000000003000000010000008f000000, /* 2535 */
128'h1b0000000f00000003000000a0000000, /* 2536 */
128'h000063746e692d7570632c7663736972, /* 2537 */
128'h01000000b50000000400000003000000, /* 2538 */
128'h01000000bb0000000400000003000000, /* 2539 */
128'h01000000020000000200000002000000, /* 2540 */
128'h0030303030303030384079726f6d656d, /* 2541 */
128'h6f6d656d5b0000000700000003000000, /* 2542 */
128'h67000000100000000300000000007972, /* 2543 */
128'h00000040000000000000008000000000, /* 2544 */
128'h0300000000636f730100000002000000, /* 2545 */
128'h03000000020000000000000004000000, /* 2546 */
128'h03000000020000000f00000004000000, /* 2547 */
128'h616972612c6874651b0000001f000000, /* 2548 */
128'h706d697300636f732d657261622d656e, /* 2549 */
128'h000000000300000000007375622d656c, /* 2550 */
128'h303240746e696c6301000000c3000000, /* 2551 */
128'h0d000000030000000000003030303030, /* 2552 */
128'h30746e696c632c76637369721b000000, /* 2553 */
128'hca000000100000000300000000000000, /* 2554 */
128'h07000000010000000300000001000000, /* 2555 */
128'h00000000670000001000000003000000, /* 2556 */
128'h0300000000000c000000000000000002, /* 2557 */
128'h006c6f72746e6f63de00000008000000, /* 2558 */
128'h7075727265746e690100000002000000, /* 2559 */
128'h3030634072656c6c6f72746e6f632d74, /* 2560 */
128'h04000000030000000000000030303030, /* 2561 */
128'h04000000030000000000000000000000, /* 2562 */
128'h0c00000003000000010000008f000000, /* 2563 */
128'h003063696c702c76637369721b000000, /* 2564 */
128'h03000000a00000000000000003000000, /* 2565 */
128'h0b00000001000000ca00000010000000, /* 2566 */
128'h10000000030000000900000001000000, /* 2567 */
128'h000000000000000c0000000067000000, /* 2568 */
128'he8000000040000000300000000000004, /* 2569 */
128'hfb000000040000000300000007000000, /* 2570 */
128'hb5000000040000000300000003000000, /* 2571 */
128'hbb000000040000000300000002000000, /* 2572 */
128'h75626564010000000200000002000000, /* 2573 */
128'h0000304072656c6c6f72746e6f632d67, /* 2574 */
128'h637369721b0000001000000003000000, /* 2575 */
128'h03000000003331302d67756265642c76, /* 2576 */
128'hffff000001000000ca00000008000000, /* 2577 */
128'h00000000670000001000000003000000, /* 2578 */
128'h03000000001000000000000000000000, /* 2579 */
128'h006c6f72746e6f63de00000008000000, /* 2580 */
128'h30303140747261750100000002000000, /* 2581 */
128'h08000000030000000000003030303030, /* 2582 */
128'h03000000003035373631736e1b000000, /* 2583 */
128'h00000010000000006700000010000000, /* 2584 */
128'h04000000030000000010000000000000, /* 2585 */
128'h040000000300000080f0fa024b000000, /* 2586 */
128'h040000000300000000c2010006010000, /* 2587 */
128'h04000000030000000200000014010000, /* 2588 */
128'h04000000030000000100000025010000, /* 2589 */
128'h04000000030000000200000030010000, /* 2590 */
128'h0100000002000000040000003a010000, /* 2591 */
128'h3030303240636d6d2d63736972776f6c, /* 2592 */
128'h10000000030000000000000030303030, /* 2593 */
128'h00000000000000200000000067000000, /* 2594 */
128'h14010000040000000300000000000100, /* 2595 */
128'h25010000040000000300000002000000, /* 2596 */
128'h1b0000000c0000000300000002000000, /* 2597 */
128'h0200000000636d6d2d63736972776f6c, /* 2598 */
128'h406874652d63736972776f6c01000000, /* 2599 */
128'h03000000000000003030303030303033, /* 2600 */
128'h2d63736972776f6c1b0000000c000000, /* 2601 */
128'h5b000000080000000300000000687465, /* 2602 */
128'h0400000003000000006b726f7774656e, /* 2603 */
128'h04000000030000000200000014010000, /* 2604 */
128'h06000000030000000300000025010000, /* 2605 */
128'h0300000000007fe3023e180047010000, /* 2606 */
128'h00000030000000006700000010000000, /* 2607 */
128'h01000000020000000080000000000000, /* 2608 */
128'h303440646e7277682d63736972776f6c, /* 2609 */
128'h0e000000030000000000303030303030, /* 2610 */
128'h6e7277682d63736972776f6c1b000000, /* 2611 */
128'h67000000100000000300000000000064, /* 2612 */
128'h00100000000000000000004000000000, /* 2613 */
128'h09000000020000000200000002000000, /* 2614 */
128'h2300736c6c65632d7373657264646123, /* 2615 */
128'h61706d6f6300736c6c65632d657a6973, /* 2616 */
128'h6f647473006c65646f6d00656c626974, /* 2617 */
128'h65736162656d697400687461702d7475, /* 2618 */
128'h6b636f6c630079636e6575716572662d, /* 2619 */
128'h63697665640079636e6575716572662d, /* 2620 */
128'h75746174730067657200657079745f65, /* 2621 */
128'h2d756d6d006173692c76637369720073, /* 2622 */
128'h230074696c70732d626c740065707974, /* 2623 */
128'h00736c6c65632d747075727265746e69, /* 2624 */
128'h6f72746e6f632d747075727265746e69, /* 2625 */
128'h646e6168702c78756e696c0072656c6c, /* 2626 */
128'h727265746e69007365676e617200656c, /* 2627 */
128'h6572006465646e657478652d73747075, /* 2628 */
128'h616d2c76637369720073656d616e2d67, /* 2629 */
128'h766373697200797469726f6972702d78, /* 2630 */
128'h70732d746e6572727563007665646e2c, /* 2631 */
128'h61702d747075727265746e6900646565, /* 2632 */
128'h0073747075727265746e6900746e6572, /* 2633 */
128'h6f692d6765720074666968732d676572, /* 2634 */
128'h63616d2d6c61636f6c0068746469772d, /* 2635 */
128'h0000000000000000737365726464612d, /* 2636 */
128'h0000000000203a642520656369766544, /* 2637 */
128'h00203a6425206563697665642073250a, /* 2638 */
128'h00000000203a6425206563697665440a, /* 2639 */
128'h000a656369766564206e776f6e6b6e75, /* 2640 */
128'h00000a2973252c73252870756b6f6f6c, /* 2641 */
128'h7265206c616e7265746e692070636864, /* 2642 */
128'h00000000000000000a7025202c726f72, /* 2643 */
128'h5145525f5043484420676e69646e6553, /* 2644 */
128'h4b434120504348440000000a54534555, /* 2645 */
128'h696c432050434844000000000000000a, /* 2646 */
128'h203a7373657264644120504920746e65, /* 2647 */
128'h0000000a64252e64252e64252e642520, /* 2648 */
128'h73657264644120504920726576726553, /* 2649 */
128'h0a64252e64252e64252e642520203a73, /* 2650 */
128'h6120726574756f520000000000000000, /* 2651 */
128'h252e64252e642520203a737365726464, /* 2652 */
128'h6b73616d2074654e0000000a64252e64, /* 2653 */
128'h64252e642520203a7373657264646120, /* 2654 */
128'h697420657361654c000a64252e64252e, /* 2655 */
128'h00000000000000000a6425203d20656d, /* 2656 */
128'h00000a22732522203d206e69616d6f64, /* 2657 */
128'h00000a22732522203d20726576726573, /* 2658 */
128'h000000000a44455050494b53204b4341, /* 2659 */
128'h000000000000000a4b414e2050434844, /* 2660 */
128'h73657264646120646574736575716552, /* 2661 */
128'h0000000000000a646573756665722073, /* 2662 */
128'h000000000000000a732520726f727245, /* 2663 */
128'h6e6f6974706f2064656c646e61686e75, /* 2664 */
128'h656c646e61686e55000000000a642520, /* 2665 */
128'h64252065646f63706f20504348442064, /* 2666 */
128'h20676e69646e6553000000000000000a, /* 2667 */
128'h000a595245564f435349445f50434844, /* 2668 */
128'h00000000000a29732528726f72726570, /* 2669 */
128'h3a2043414d2073250000000030687465, /* 2670 */
128'h3a583230253a583230253a5832302520, /* 2671 */
128'h000a583230253a583230253a58323025, /* 2672 */
128'h484420646e65732074276e646c756f43, /* 2673 */
128'h206e6f20595245564f43534944205043, /* 2674 */
128'h00000a7325203a732520656369766564, /* 2675 */
128'h5043484420726f6620676e6974696157, /* 2676 */
128'h2020202020202020000a524546464f5f, /* 2677 */
128'h00000000000063250000000000000020, /* 2678 */
128'h0000005832302520000000000000002e, /* 2679 */
128'h00000000732573250000000000000a0a, /* 2680 */
128'h00000000007325203a646c697542202c, /* 2681 */
128'h73257a4820756c250000000000007325, /* 2682 */
128'h0000000000756c250000000000000000, /* 2683 */
128'h0073257a4863252000000000646c252e, /* 2684 */
128'h00000000007325736574794220756c25, /* 2685 */
128'h00003a786c3830250073254269632520, /* 2686 */
128'h000a73252020202000786c6c2a302520, /* 2687 */
128'h000000203a5d64255b6e6f6974636553, /* 2688 */
128'h25203d206465726975716572206e656c, /* 2689 */
128'h000a7825203d206c6175746361202c58, /* 2690 */
128'h302c782578302c7825287970636d656d, /* 2691 */
128'h25287465736d656d00000a3b29782578, /* 2692 */
128'h00000000000a3b29782578302c302c78, /* 2693 */
128'h0000000054455346464f5f4f4c43414d, /* 2694 */
128'h0000000054455346464f5f494843414d, /* 2695 */
128'h000000000054455346464f5f524c5054, /* 2696 */
128'h000000000054455346464f5f53434654, /* 2697 */
128'h0054455346464f5f4c5254434f49444d, /* 2698 */
128'h000000000054455346464f5f53434652, /* 2699 */
128'h00000000000054455346464f5f525352, /* 2700 */
128'h000000000054455346464f5f44414252, /* 2701 */
128'h000000000054455346464f5f524c5052, /* 2702 */
128'h46464f5f524c5052000000003f3f3f3f, /* 2703 */
128'h0000000000000047000064252b544553, /* 2704 */
128'h0a50495049203d206f746f7250205049, /* 2705 */
128'h00000000000000540000000000000000, /* 2706 */
128'h000a504745203d206f746f7250205049, /* 2707 */
128'h000a505550203d206f746f7250205049, /* 2708 */
128'h0000000a3a7265646165682074736574, /* 2709 */
128'h000a3a73746e65746e6f632074736574, /* 2710 */
128'h000a504449203d206f746f7250205049, /* 2711 */
128'h00000a5054203d206f746f7250205049, /* 2712 */
128'h0a50434344203d206f746f7250205049, /* 2713 */
128'h00000000000000360000000000000000, /* 2714 */
128'h0a50565352203d206f746f7250205049, /* 2715 */
128'h6f746f72502050490000000000000000, /* 2716 */
128'h6f746f7250205049000a455247203d20, /* 2717 */
128'h6f746f7250205049000a505345203d20, /* 2718 */
128'h6f746f725020504900000a4841203d20, /* 2719 */
128'h6f746f7250205049000a50544d203d20, /* 2720 */
128'h0000000000000a485054454542203d20, /* 2721 */
128'h5041434e45203d206f746f7250205049, /* 2722 */
128'h000000000000004d000000000000000a, /* 2723 */
128'h0a504d4f43203d206f746f7250205049, /* 2724 */
128'h6f746f72502050490000000000000000, /* 2725 */
128'h00000000000000000a50544353203d20, /* 2726 */
128'h494c504455203d206f746f7250205049, /* 2727 */
128'h6f746f725020504900000000000a4554, /* 2728 */
128'h00000000000000000a534c504d203d20, /* 2729 */
128'h000a574152203d206f746f7250205049, /* 2730 */
128'h7075736e75203d206f746f7270205049, /* 2731 */
128'h000000000a2978252820646574726f70, /* 2732 */
128'h257830203d20657079745f6f746f7270, /* 2733 */
128'h656c646e61686e750000000000000a78, /* 2734 */
128'h0000000a21747075727265746e692064, /* 2735 */
128'h000a726464612043414d207075746553, /* 2736 */
128'h00000a786c253a786c25203d2043414d, /* 2737 */
128'h3025203d20737365726464612043414d, /* 2738 */
128'h3230253a783230253a783230253a7832, /* 2739 */
128'h0000000a2e783230253a783230253a78, /* 2740 */
128'h75727265746e692074656e7265687445, /* 2741 */
128'h0a646c25203d20737574617473207470, /* 2742 */
128'h65687420746f6f420000000000000000, /* 2743 */
128'h2e6d6172676f727020646564616f6c20, /* 2744 */
128'h2c657962646f6f4700000000000a2e2e, /* 2745 */
128'h000000000a2e2e2e207265746f6f6220, /* 2746 */
128'h00007f7c5d5b3f3e3d3c3b3a2c2b2a22, /* 2747 */
128'h007f7c5d5b3f3e3d3c3b3a2e2c2b2a22, /* 2748 */
128'h66656463626139383736353433323130, /* 2749 */
128'h72776f6c2f6372730000000000000000, /* 2750 */
128'h00000000000000632e636d6d5f637369, /* 2751 */
128'h61625f6473203d3d20657361625f6473, /* 2752 */
128'h5f63736972776f6c00726464615f6573, /* 2753 */
128'h000a74756f656d6974207325203a6473, /* 2754 */
128'h616d202c6465766f6d65722064726143, /* 2755 */
128'h6425206f74206465676e616863206b73, /* 2756 */
128'h736e692064726143000000000000000a, /* 2757 */
128'h6e616863206b73616d202c6465747265, /* 2758 */
128'h0000000000000a6425206f7420646567, /* 2759 */
128'h25207461206465746165726320636d6d, /* 2760 */
128'h0000000a7825203d2074736f68202c78, /* 2761 */
128'h0000000000006f4e0000000000736559, /* 2762 */
128'h002020203a434d4d0000000052444420, /* 2763 */
128'h00000000000a7325203a656369766544, /* 2764 */
128'h3a4449207265727574636166756e614d, /* 2765 */
128'h0a7825203a4d454f000000000a782520, /* 2766 */
128'h6325203a656d614e0000000000000000, /* 2767 */
128'h0000000000000a206325632563256325, /* 2768 */
128'h00000a6425203a646565705320737542, /* 2769 */
128'h25203a79746963617061432068676948, /* 2770 */
128'h79746963617061430000000000000a73, /* 2771 */
128'h7464695720737542000000000000203a, /* 2772 */
128'h000000000a73257469622d6425203a68, /* 2773 */
128'h0000007825782520000000203a78250a, /* 2774 */
128'h00000000000064735f63736972776f6c, /* 2775 */
128'h0000000065646f6d206e776f6e6b6e55, /* 2776 */
128'h7830203a726f72724520737574617453, /* 2777 */
128'h2074756f656d69540000000a58383025, /* 2778 */
128'h616572206472616320676e6974696177, /* 2779 */
128'h6c69616620636d6d00000000000a7964, /* 2780 */
128'h6d6320706f747320646e6573206f7420, /* 2781 */
128'h6f6c62203a434d4d0000000000000a64, /* 2782 */
128'h20786c257830207265626d756e206b63, /* 2783 */
128'h6c2578302878616d2073646565637865, /* 2784 */
128'h203d3e20434d4d6500000000000a2978, /* 2785 */
128'h726f6620646572697571657220342e34, /* 2786 */
128'h642072657375206465636e61686e6520, /* 2787 */
128'h000000000000000a6165726120617461, /* 2788 */
128'h757320746f6e2073656f642064726143, /* 2789 */
128'h696e6f697469747261702074726f7070, /* 2790 */
128'h656f64206472614300000000000a676e, /* 2791 */
128'h20434820656e6966656420746f6e2073, /* 2792 */
128'h00000a657a69732070756f7267205057, /* 2793 */
128'h636e61686e6520617461642072657355, /* 2794 */
128'h5720434820746f6e2061657261206465, /* 2795 */
128'h696c6120657a69732070756f72672050, /* 2796 */
128'h72617020692550470000000a64656e67, /* 2797 */
128'h505720434820746f6e206e6f69746974, /* 2798 */
128'h67696c6120657a69732070756f726720, /* 2799 */
128'h656f642064726143000000000a64656e, /* 2800 */
128'h6e652074726f7070757320746f6e2073, /* 2801 */
128'h657475626972747461206465636e6168, /* 2802 */
128'h6e65206c61746f54000000000000000a, /* 2803 */
128'h6563786520657a6973206465636e6168, /* 2804 */
128'h20752528206d756d6978616d20736465, /* 2805 */
128'h656f64206472614300000a297525203e, /* 2806 */
128'h6f682074726f7070757320746f6e2073, /* 2807 */
128'h61702064656c6c6f72746e6f63207473, /* 2808 */
128'h6572206574697277206e6f6974697472, /* 2809 */
128'h6e6974746573207974696c696261696c, /* 2810 */
128'h726c61206472614300000000000a7367, /* 2811 */
128'h64656e6f697469747261702079646165, /* 2812 */
128'h206f6e203a434d4d000000000000000a, /* 2813 */
128'h0000000a746e65736572702064726163, /* 2814 */
128'h73657220746f6e206469642064726143, /* 2815 */
128'h20656761746c6f76206f7420646e6f70, /* 2816 */
128'h00000000000000000a217463656c6573, /* 2817 */
128'h7463656c6573206f7420656c62616e75, /* 2818 */
128'h00000000000000000a65646f6d206120, /* 2819 */
128'h646e756f66206473635f747865206f4e, /* 2820 */
128'h78363025206e614d0000000000000a21, /* 2821 */
128'h000000783430257834302520726e5320, /* 2822 */
128'h00000000632563256325632563256325, /* 2823 */
128'h6167656c20434d4d00000064252e6425, /* 2824 */
128'h636167654c2044530000000000007963, /* 2825 */
128'h6867694820434d4d0000000000000079, /* 2826 */
128'h0000297a484d36322820646565705320, /* 2827 */
128'h35282064656570532068676948204453, /* 2828 */
128'h6867694820434d4d000000297a484d30, /* 2829 */
128'h0000297a484d32352820646565705320, /* 2830 */
128'h7a484d32352820323552444420434d4d, /* 2831 */
128'h31524453205348550000000000000029, /* 2832 */
128'h00000000000000297a484d3532282032, /* 2833 */
128'h7a484d30352820353252445320534855, /* 2834 */
128'h35524453205348550000000000000029, /* 2835 */
128'h000000000000297a484d303031282030, /* 2836 */
128'h7a484d30352820303552444420534855, /* 2837 */
128'h31524453205348550000000000000029, /* 2838 */
128'h0000000000297a484d38303228203430, /* 2839 */
128'h0000297a484d30303228203030325348, /* 2840 */
128'h6f6e2064252065636976654420434d4d, /* 2841 */
128'h00000000000000000a646e756f662074, /* 2842 */
128'h000000000000445300000000434d4d65, /* 2843 */
128'h000000297325282000006425203a7325, /* 2844 */
128'h6e656c20656c69460000000000636d6d, /* 2845 */
128'h000000000000000a6425203d20687467, /* 2846 */
128'h0a7325203d202964252c70252835646d, /* 2847 */
128'h20747365757165520000000000000000, /* 2848 */
128'h25202e676e6f6c206f6f742068746170, /* 2849 */
128'h000000000000002f00000000000a646c, /* 2850 */
128'h6b636f6c62202c22732522203a717277, /* 2851 */
128'h00000000000000000a64253d657a6973, /* 2852 */
128'h646e6520656c69662065766965636552, /* 2853 */
128'h775f656c646e61680000000000000a2e, /* 2854 */
128'h00000000000a2e64656c6c6163207172, /* 2855 */
128'h65706f2050544654206c6167656c6c49, /* 2856 */
128'h00000000000000000a2e6e6f69746172, /* 2857 */
128'h445320746e756f6d206f74206c696146, /* 2858 */
128'h000000000000000a2172657669726420, /* 2859 */
128'h6e69206e69622e746f6f622064616f4c, /* 2860 */
128'h0000000000000a79726f6d656d206f74, /* 2861 */
128'h00000000000000006e69622e746f6f62, /* 2862 */
128'h62206e65706f206f742064656c696146, /* 2863 */
128'h206f74206c6961660000000a21746f6f, /* 2864 */
128'h000000000021656c69662065736f6c63, /* 2865 */
128'h6420746e756f6d75206f74206c696166, /* 2866 */
128'h2520646564616f4c00000000216b7369, /* 2867 */
128'h726f6d656d206f742073657479622064, /* 2868 */
128'h6f726620782520737365726464612079, /* 2869 */
128'h642520666f206e69622e746f6f62206d, /* 2870 */
128'h00000000000000000a2e736574796220, /* 2871 */
128'h20524444206f7420666c652064616f6c, /* 2872 */
128'h6461657220666c65000a79726f6d656d, /* 2873 */
128'h646f6320687469772064656c69616620, /* 2874 */
128'h000000005c2d2f7c0000000064252065, /* 2875 */
128'h696620646573616220746f6f622d750a, /* 2876 */
128'h6c20746f6f6220656761747320747372, /* 2877 */
128'h6f6974726573736100000a726564616f, /* 2878 */
128'h6c6966202c64656c696166207325206e, /* 2879 */
128'h66202c642520656e696c202c73252065, /* 2880 */
128'h00000000000a7325206e6f6974636e75, /* 2881 */
128'h3d212078257830203a4552554c494146, /* 2882 */
128'h2074657366666f207461207825783020, /* 2883 */
128'h2c7025203d20317000000a2e78257830, /* 2884 */
128'h000000000000000a7025203d20327020, /* 2885 */
128'h00000000002020202020202020202020, /* 2886 */
128'h00000000000808080808080808080808, /* 2887 */
128'h000000000000752520676e6974746573, /* 2888 */
128'h000000000000752520676e6974736574, /* 2889 */
128'h6c626973736f70203a4552554c494146, /* 2890 */
128'h696c2073736572646461206461622065, /* 2891 */
128'h2578302074657366666f20746120656e, /* 2892 */
128'h676e697070696b5300000000000a2e78, /* 2893 */
128'h2e2e2e74736574207478656e206f7420, /* 2894 */
128'h0808080808080808000000000000000a, /* 2895 */
128'h08082020202020202020202020080808, /* 2896 */
128'h00000000000000080808080808080808, /* 2897 */
128'h6e617220747365740000000000082008, /* 2898 */
128'h7830206f742070257830207369206567, /* 2899 */
128'h00752520706f6f4c00000000000a7025, /* 2900 */
128'h0000000000000a3a000000000075252f, /* 2901 */
128'h00000073736572646441206b63757453, /* 2902 */
128'h00000000000a6b6f0000203a73252020, /* 2903 */
128'h656d20657261420a00000a2e656e6f44, /* 2904 */
128'h00000a74736574204d415244206c6174, /* 2905 */
128'h6f6973726576207265747365746d656d, /* 2906 */
128'h297469622d64252820302e332e34206e, /* 2907 */
128'h6867697279706f43000000000000000a, /* 2908 */
128'h20323130322d31303032202943282074, /* 2909 */
128'h2e6e6f62617a61432073656c72616843, /* 2910 */
128'h6465736e6563694c000000000000000a, /* 2911 */
128'h4720554e4720656874207265646e7520, /* 2912 */
128'h694c2063696c627550206c6172656e65, /* 2913 */
128'h2032206e6f69737265762065736e6563, /* 2914 */
128'h00000000000000000a2e29796c6e6f28, /* 2915 */
128'h6425203d207465735f676e696b726f77, /* 2916 */
128'h7463757274736e6920646c25202c424b, /* 2917 */
128'h73656c63796320646c25202c736e6f69, /* 2918 */
128'h0a646c252e646c25203d20495043202c, /* 2919 */
128'h6f57206f6c6c65480000000000000000, /* 2920 */
128'h732068637469775300000a0d21646c72, /* 2921 */
128'h000a58252c5825203d20676e69747465, /* 2922 */
128'h5825203d2064656573206d6f646e6152, /* 2923 */
128'h0a746f6f62204453000000000000000a, /* 2924 */
128'h736574204d4152440000000000000000, /* 2925 */
128'h6f6f6220505446540000000000000a74, /* 2926 */
128'h65742065686361430000000000000a74, /* 2927 */
128'h00000a0d7061727400000000000a7473, /* 2928 */
128'hefcdab8967452301cccccccccccccccd, /* 2929 */
128'h10000000200000001032547698badcfe, /* 2930 */
128'h55555555555555555851f42d4c957f2d, /* 2931 */
128'h0000000000000000aaaaaaaaaaaaaaaa, /* 2932 */
128'h00000000000000000000000000000000, /* 2933 */
128'h00000000000000000000000000000000, /* 2934 */
128'h00000000000000000000000000000000, /* 2935 */
128'h00000000000000000000000000000000, /* 2936 */
128'h00000000000000000000000000000000, /* 2937 */
128'h00000000000000000000000000000000, /* 2938 */
128'h00000000000000000000000000000000, /* 2939 */
128'h00000000000000000000000000000000, /* 2940 */
128'h00000000000000000000000000000000, /* 2941 */
128'h00000000000000000000000000000000, /* 2942 */
128'h00000000000000000000000000000000, /* 2943 */
128'h00004b4d47545045000000030f060301, /* 2944 */
128'h000000003000000000000000004b4d47, /* 2945 */
128'h00000000ffffffff0000000000000000, /* 2946 */
128'h0000646d635f6473000000000c000000, /* 2947 */
128'h00000000ffffffff00006772615f6473, /* 2948 */
128'h000000002f7c5c2d00000000bffeb018, /* 2949 */
128'h0000000600000000bffeb1d0cc33aa55, /* 2950 */
128'hbffe70840000000000000000ffffffff, /* 2951 */
128'h00000000000000000000000000000000, /* 2952 */
128'h00000000000000000000000000000000, /* 2953 */
128'h00000000000000000000000000000000, /* 2954 */
128'h00000000000000000000000000000000, /* 2955 */
128'h00000000000000000000000000000000, /* 2956 */
128'h00000000000000000000000000000000, /* 2957 */
128'h00000000000000000000000000000000, /* 2958 */
128'h00000000000000000000000000000000, /* 2959 */
128'h00000000000000000000000000000000, /* 2960 */
128'h00000000000000000000000000000000, /* 2961 */
128'h00000000000000000000000000000000, /* 2962 */
128'h00000000000000000000000000000000, /* 2963 */
128'h00000000000000000000000000000000, /* 2964 */
128'h00000000000000000000000000000000, /* 2965 */
128'h00000000000000000000000000000000, /* 2966 */
128'h00000000000000000000000000000000, /* 2967 */
128'h00000000000000000000000000000000, /* 2968 */
128'h00000000000000000000000000000000, /* 2969 */
128'h00000000000000000000000000000000, /* 2970 */
128'h00000000000000000000000000000000, /* 2971 */
128'h00000000000000000000000000000000, /* 2972 */
128'h00000000000000000000000000000000, /* 2973 */
128'h00000000000000000000000000000000, /* 2974 */
128'h00000000000000000000000000000000, /* 2975 */
128'h00000000000000000000000000000000, /* 2976 */
128'h00000000000000000000000000000000, /* 2977 */
128'h00000000000000000000000000000000, /* 2978 */
128'h00000000000000000000000000000000, /* 2979 */
128'h00000000000000000000000000000000, /* 2980 */
128'h00000000000000000000000000000000, /* 2981 */
128'h00000000000000000000000000000000, /* 2982 */
128'h00000000000000000000000000000000, /* 2983 */
128'h00000000000000000000000000000000, /* 2984 */
128'h00000000000000000000000000000000, /* 2985 */
128'h00000000000000000000000000000000, /* 2986 */
128'h00000000000000000000000000000000, /* 2987 */
128'h00000000000000000000000000000000, /* 2988 */
128'h00000000000000000000000000000000, /* 2989 */
128'h00000000000000000000000000000000, /* 2990 */
128'h00000000000000000000000000000000, /* 2991 */
128'h00000000000000000000000000000000, /* 2992 */
128'h00000000000000000000000000000000, /* 2993 */
128'h00000000000000000000000000000000, /* 2994 */
128'h00000000000000000000000000000000, /* 2995 */
128'h00000000000000000000000000000000, /* 2996 */
128'h00000000000000000000000000000000, /* 2997 */
128'h00000000000000000000000000000000, /* 2998 */
128'h00000000000000000000000000000000, /* 2999 */
128'h00000000000000000000000000000000, /* 3000 */
128'h00000000000000000000000000000000, /* 3001 */
128'h00000000000000000000000000000000, /* 3002 */
128'h00000000000000000000000000000000, /* 3003 */
128'h00000000000000000000000000000000, /* 3004 */
128'h00000000000000000000000000000000, /* 3005 */
128'h00000000000000000000000000000000, /* 3006 */
128'h00000000000000000000000000000000, /* 3007 */
128'h00000000000000000000000000000000, /* 3008 */
128'h00000000000000000000000000000000, /* 3009 */
128'h00000000000000000000000000000000, /* 3010 */
128'h00000000000000000000000000000000, /* 3011 */
128'h00000000000000000000000000000000, /* 3012 */
128'h00000000000000000000000000000000, /* 3013 */
128'h00000000000000000000000000000000, /* 3014 */
128'h00000000000000000000000000000000, /* 3015 */
128'h00000000000000000000000000000000, /* 3016 */
128'h00000000000000000000000000000000, /* 3017 */
128'h00000000000000000000000000000000, /* 3018 */
128'h00000000000000000000000000000000, /* 3019 */
128'h00000000000000000000000000000000, /* 3020 */
128'h00000000000000000000000000000000, /* 3021 */
128'h00000000000000000000000000000000, /* 3022 */
128'h00000000000000000000000000000000, /* 3023 */
128'h00000000000000000000000000000000, /* 3024 */
128'h00000000000000000000000000000000, /* 3025 */
128'h00000000000000000000000000000000, /* 3026 */
128'h00000000000000000000000000000000, /* 3027 */
128'h00000000000000000000000000000000, /* 3028 */
128'h00000000000000000000000000000000, /* 3029 */
128'h00000000000000000000000000000000, /* 3030 */
128'h00000000000000000000000000000000, /* 3031 */
128'h00000000000000000000000000000000, /* 3032 */
128'h00000000000000000000000000000000, /* 3033 */
128'h00000000000000000000000000000000, /* 3034 */
128'h00000000000000000000000000000000, /* 3035 */
128'h00000000000000000000000000000000, /* 3036 */
128'h00000000000000000000000000000000, /* 3037 */
128'h00000000000000000000000000000000, /* 3038 */
128'h00000000000000000000000000000000, /* 3039 */
128'h00000000000000000000000000000000, /* 3040 */
128'h00000000000000000000000000000000, /* 3041 */
128'h00000000000000000000000000000000, /* 3042 */
128'h00000000000000000000000000000000, /* 3043 */
128'h00000000000000000000000000000000, /* 3044 */
128'h00000000000000000000000000000000, /* 3045 */
128'h00000000000000000000000000000000, /* 3046 */
128'h00000000000000000000000000000000, /* 3047 */
128'h00000000000000000000000000000000, /* 3048 */
128'h00000000000000000000000000000000, /* 3049 */
128'h00000000000000000000000000000000, /* 3050 */
128'h00000000000000000000000000000000, /* 3051 */
128'h00000000000000000000000000000000, /* 3052 */
128'h00000000000000000000000000000000, /* 3053 */
128'h00000000000000000000000000000000, /* 3054 */
128'h00000000000000000000000000000000, /* 3055 */
128'h00000000000000000000000000000000, /* 3056 */
128'h00000000000000000000000000000000, /* 3057 */
128'h00000000000000000000000000000000, /* 3058 */
128'h00000000000000000000000000000000, /* 3059 */
128'h00000000000000000000000000000000, /* 3060 */
128'h00000000000000000000000000000000, /* 3061 */
128'h00000000000000000000000000000000, /* 3062 */
128'h00000000000000000000000000000000, /* 3063 */
128'h00000000000000000000000000000000, /* 3064 */
128'h00000000000000000000000000000000, /* 3065 */
128'h00000000000000000000000000000000, /* 3066 */
128'h00000000000000000000000000000000, /* 3067 */
128'h00000000000000000000000000000000, /* 3068 */
128'h00000000000000000000000000000000, /* 3069 */
128'h00000000000000000000000000000000, /* 3070 */
128'h00000000000000000000000000000000, /* 3071 */
128'h00000000000000000000000000000000, /* 3072 */
128'h00000000000000000000000000000000, /* 3073 */
128'h00000000000000000000000000000000, /* 3074 */
128'h00000000000000000000000000000000, /* 3075 */
128'h00000000000000000000000000000000, /* 3076 */
128'h00000000000000000000000000000000, /* 3077 */
128'h00000000000000000000000000000000, /* 3078 */
128'h00000000000000000000000000000000, /* 3079 */
128'h00000000000000000000000000000000, /* 3080 */
128'h00000000000000000000000000000000, /* 3081 */
128'h00000000000000000000000000000000, /* 3082 */
128'h00000000000000000000000000000000, /* 3083 */
128'h00000000000000000000000000000000, /* 3084 */
128'h00000000000000000000000000000000, /* 3085 */
128'h00000000000000000000000000000000, /* 3086 */
128'h00000000000000000000000000000000, /* 3087 */
128'h00000000000000000000000000000000, /* 3088 */
128'h00000000000000000000000000000000, /* 3089 */
128'h00000000000000000000000000000000, /* 3090 */
128'h00000000000000000000000000000000, /* 3091 */
128'h00000000000000000000000000000000, /* 3092 */
128'h00000000000000000000000000000000, /* 3093 */
128'h00000000000000000000000000000000, /* 3094 */
128'h00000000000000000000000000000000, /* 3095 */
128'h00000000000000000000000000000000, /* 3096 */
128'h00000000000000000000000000000000, /* 3097 */
128'h00000000000000000000000000000000, /* 3098 */
128'h00000000000000000000000000000000, /* 3099 */
128'h00000000000000000000000000000000, /* 3100 */
128'h00000000000000000000000000000000, /* 3101 */
128'h00000000000000000000000000000000, /* 3102 */
128'h00000000000000000000000000000000, /* 3103 */
128'h00000000000000000000000000000000, /* 3104 */
128'h00000000000000000000000000000000, /* 3105 */
128'h00000000000000000000000000000000, /* 3106 */
128'h00000000000000000000000000000000, /* 3107 */
128'h00000000000000000000000000000000, /* 3108 */
128'h00000000000000000000000000000000, /* 3109 */
128'h00000000000000000000000000000000, /* 3110 */
128'h00000000000000000000000000000000, /* 3111 */
128'h00000000000000000000000000000000, /* 3112 */
128'h00000000000000000000000000000000, /* 3113 */
128'h00000000000000000000000000000000, /* 3114 */
128'h00000000000000000000000000000000, /* 3115 */
128'h00000000000000000000000000000000, /* 3116 */
128'h00000000000000000000000000000000, /* 3117 */
128'h00000000000000000000000000000000, /* 3118 */
128'h00000000000000000000000000000000, /* 3119 */
128'h00000000000000000000000000000000, /* 3120 */
128'h00000000000000000000000000000000, /* 3121 */
128'h00000000000000000000000000000000, /* 3122 */
128'h00000000000000000000000000000000, /* 3123 */
128'h00000000000000000000000000000000, /* 3124 */
128'h00000000000000000000000000000000, /* 3125 */
128'h00000000000000000000000000000000, /* 3126 */
128'h00000000000000000000000000000000, /* 3127 */
128'h00000000000000000000000000000000, /* 3128 */
128'h00000000000000000000000000000000, /* 3129 */
128'h00000000000000000000000000000000, /* 3130 */
128'h00000000000000000000000000000000, /* 3131 */
128'h00000000000000000000000000000000, /* 3132 */
128'h00000000000000000000000000000000, /* 3133 */
128'h00000000000000000000000000000000, /* 3134 */
128'h00000000000000000000000000000000, /* 3135 */
128'h00000000000000000000000000000000, /* 3136 */
128'h00000000000000000000000000000000, /* 3137 */
128'h00000000000000000000000000000000, /* 3138 */
128'h00000000000000000000000000000000, /* 3139 */
128'h00000000000000000000000000000000, /* 3140 */
128'h00000000000000000000000000000000, /* 3141 */
128'h00000000000000000000000000000000, /* 3142 */
128'h00000000000000000000000000000000, /* 3143 */
128'h00000000000000000000000000000000, /* 3144 */
128'h00000000000000000000000000000000, /* 3145 */
128'h00000000000000000000000000000000, /* 3146 */
128'h00000000000000000000000000000000, /* 3147 */
128'h00000000000000000000000000000000, /* 3148 */
128'h00000000000000000000000000000000, /* 3149 */
128'h00000000000000000000000000000000, /* 3150 */
128'h00000000000000000000000000000000, /* 3151 */
128'h00000000000000000000000000000000, /* 3152 */
128'h00000000000000000000000000000000, /* 3153 */
128'h00000000000000000000000000000000, /* 3154 */
128'h00000000000000000000000000000000, /* 3155 */
128'h00000000000000000000000000000000, /* 3156 */
128'h00000000000000000000000000000000, /* 3157 */
128'h00000000000000000000000000000000, /* 3158 */
128'h00000000000000000000000000000000, /* 3159 */
128'h00000000000000000000000000000000, /* 3160 */
128'h00000000000000000000000000000000, /* 3161 */
128'h00000000000000000000000000000000, /* 3162 */
128'h00000000000000000000000000000000, /* 3163 */
128'h00000000000000000000000000000000, /* 3164 */
128'h00000000000000000000000000000000, /* 3165 */
128'h00000000000000000000000000000000, /* 3166 */
128'h00000000000000000000000000000000, /* 3167 */
128'h00000000000000000000000000000000, /* 3168 */
128'h00000000000000000000000000000000, /* 3169 */
128'h00000000000000000000000000000000, /* 3170 */
128'h00000000000000000000000000000000, /* 3171 */
128'h00000000000000000000000000000000, /* 3172 */
128'h00000000000000000000000000000000, /* 3173 */
128'h00000000000000000000000000000000, /* 3174 */
128'h00000000000000000000000000000000, /* 3175 */
128'h00000000000000000000000000000000, /* 3176 */
128'h00000000000000000000000000000000, /* 3177 */
128'h00000000000000000000000000000000, /* 3178 */
128'h00000000000000000000000000000000, /* 3179 */
128'h00000000000000000000000000000000, /* 3180 */
128'h00000000000000000000000000000000, /* 3181 */
128'h00000000000000000000000000000000, /* 3182 */
128'h00000000000000000000000000000000, /* 3183 */
128'h00000000000000000000000000000000, /* 3184 */
128'h00000000000000000000000000000000, /* 3185 */
128'h00000000000000000000000000000000, /* 3186 */
128'h00000000000000000000000000000000, /* 3187 */
128'h00000000000000000000000000000000, /* 3188 */
128'h00000000000000000000000000000000, /* 3189 */
128'h00000000000000000000000000000000, /* 3190 */
128'h00000000000000000000000000000000, /* 3191 */
128'h00000000000000000000000000000000, /* 3192 */
128'h00000000000000000000000000000000, /* 3193 */
128'h00000000000000000000000000000000, /* 3194 */
128'h00000000000000000000000000000000, /* 3195 */
128'h00000000000000000000000000000000, /* 3196 */
128'h00000000000000000000000000000000, /* 3197 */
128'h00000000000000000000000000000000, /* 3198 */
128'h00000000000000000000000000000000, /* 3199 */
128'h00000000000000000000000000000000, /* 3200 */
128'h00000000000000000000000000000000, /* 3201 */
128'h00000000000000000000000000000000, /* 3202 */
128'h00000000000000000000000000000000, /* 3203 */
128'h00000000000000000000000000000000, /* 3204 */
128'h00000000000000000000000000000000, /* 3205 */
128'h00000000000000000000000000000000, /* 3206 */
128'h00000000000000000000000000000000, /* 3207 */
128'h00000000000000000000000000000000, /* 3208 */
128'h00000000000000000000000000000000, /* 3209 */
128'h00000000000000000000000000000000, /* 3210 */
128'h00000000000000000000000000000000, /* 3211 */
128'h00000000000000000000000000000000, /* 3212 */
128'h00000000000000000000000000000000, /* 3213 */
128'h00000000000000000000000000000000, /* 3214 */
128'h00000000000000000000000000000000, /* 3215 */
128'h00000000000000000000000000000000, /* 3216 */
128'h00000000000000000000000000000000, /* 3217 */
128'h00000000000000000000000000000000, /* 3218 */
128'h00000000000000000000000000000000, /* 3219 */
128'h00000000000000000000000000000000, /* 3220 */
128'h00000000000000000000000000000000, /* 3221 */
128'h00000000000000000000000000000000, /* 3222 */
128'h00000000000000000000000000000000, /* 3223 */
128'h00000000000000000000000000000000, /* 3224 */
128'h00000000000000000000000000000000, /* 3225 */
128'h00000000000000000000000000000000, /* 3226 */
128'h00000000000000000000000000000000, /* 3227 */
128'h00000000000000000000000000000000, /* 3228 */
128'h00000000000000000000000000000000, /* 3229 */
128'h00000000000000000000000000000000, /* 3230 */
128'h00000000000000000000000000000000, /* 3231 */
128'h00000000000000000000000000000000, /* 3232 */
128'h00000000000000000000000000000000, /* 3233 */
128'h00000000000000000000000000000000, /* 3234 */
128'h00000000000000000000000000000000, /* 3235 */
128'h00000000000000000000000000000000, /* 3236 */
128'h00000000000000000000000000000000, /* 3237 */
128'h00000000000000000000000000000000, /* 3238 */
128'h00000000000000000000000000000000, /* 3239 */
128'h00000000000000000000000000000000, /* 3240 */
128'h00000000000000000000000000000000, /* 3241 */
128'h00000000000000000000000000000000, /* 3242 */
128'h00000000000000000000000000000000, /* 3243 */
128'h00000000000000000000000000000000, /* 3244 */
128'h00000000000000000000000000000000, /* 3245 */
128'h00000000000000000000000000000000, /* 3246 */
128'h00000000000000000000000000000000, /* 3247 */
128'h00000000000000000000000000000000, /* 3248 */
128'h00000000000000000000000000000000, /* 3249 */
128'h00000000000000000000000000000000, /* 3250 */
128'h00000000000000000000000000000000, /* 3251 */
128'h00000000000000000000000000000000, /* 3252 */
128'h00000000000000000000000000000000, /* 3253 */
128'h00000000000000000000000000000000, /* 3254 */
128'h00000000000000000000000000000000, /* 3255 */
128'h00000000000000000000000000000000, /* 3256 */
128'h00000000000000000000000000000000, /* 3257 */
128'h00000000000000000000000000000000, /* 3258 */
128'h00000000000000000000000000000000, /* 3259 */
128'h00000000000000000000000000000000, /* 3260 */
128'h00000000000000000000000000000000, /* 3261 */
128'h00000000000000000000000000000000, /* 3262 */
128'h00000000000000000000000000000000, /* 3263 */
128'h00000000000000000000000000000000, /* 3264 */
128'h00000000000000000000000000000000, /* 3265 */
128'h00000000000000000000000000000000, /* 3266 */
128'h00000000000000000000000000000000, /* 3267 */
128'h00000000000000000000000000000000, /* 3268 */
128'h00000000000000000000000000000000, /* 3269 */
128'h00000000000000000000000000000000, /* 3270 */
128'h00000000000000000000000000000000, /* 3271 */
128'h00000000000000000000000000000000, /* 3272 */
128'h00000000000000000000000000000000, /* 3273 */
128'h00000000000000000000000000000000, /* 3274 */
128'h00000000000000000000000000000000, /* 3275 */
128'h00000000000000000000000000000000, /* 3276 */
128'h00000000000000000000000000000000, /* 3277 */
128'h00000000000000000000000000000000, /* 3278 */
128'h00000000000000000000000000000000, /* 3279 */
128'h00000000000000000000000000000000, /* 3280 */
128'h00000000000000000000000000000000, /* 3281 */
128'h00000000000000000000000000000000, /* 3282 */
128'h00000000000000000000000000000000, /* 3283 */
128'h00000000000000000000000000000000, /* 3284 */
128'h00000000000000000000000000000000, /* 3285 */
128'h00000000000000000000000000000000, /* 3286 */
128'h00000000000000000000000000000000, /* 3287 */
128'h00000000000000000000000000000000, /* 3288 */
128'h00000000000000000000000000000000, /* 3289 */
128'h00000000000000000000000000000000, /* 3290 */
128'h00000000000000000000000000000000, /* 3291 */
128'h00000000000000000000000000000000, /* 3292 */
128'h00000000000000000000000000000000, /* 3293 */
128'h00000000000000000000000000000000, /* 3294 */
128'h00000000000000000000000000000000, /* 3295 */
128'h00000000000000000000000000000000, /* 3296 */
128'h00000000000000000000000000000000, /* 3297 */
128'h00000000000000000000000000000000, /* 3298 */
128'h00000000000000000000000000000000, /* 3299 */
128'h00000000000000000000000000000000, /* 3300 */
128'h00000000000000000000000000000000, /* 3301 */
128'h00000000000000000000000000000000, /* 3302 */
128'h00000000000000000000000000000000, /* 3303 */
128'h00000000000000000000000000000000, /* 3304 */
128'h00000000000000000000000000000000, /* 3305 */
128'h00000000000000000000000000000000, /* 3306 */
128'h00000000000000000000000000000000, /* 3307 */
128'h00000000000000000000000000000000, /* 3308 */
128'h00000000000000000000000000000000, /* 3309 */
128'h00000000000000000000000000000000, /* 3310 */
128'h00000000000000000000000000000000, /* 3311 */
128'h00000000000000000000000000000000, /* 3312 */
128'h00000000000000000000000000000000, /* 3313 */
128'h00000000000000000000000000000000, /* 3314 */
128'h00000000000000000000000000000000, /* 3315 */
128'h00000000000000000000000000000000, /* 3316 */
128'h00000000000000000000000000000000, /* 3317 */
128'h00000000000000000000000000000000, /* 3318 */
128'h00000000000000000000000000000000, /* 3319 */
128'h00000000000000000000000000000000, /* 3320 */
128'h00000000000000000000000000000000, /* 3321 */
128'h00000000000000000000000000000000, /* 3322 */
128'h00000000000000000000000000000000, /* 3323 */
128'h00000000000000000000000000000000, /* 3324 */
128'h00000000000000000000000000000000, /* 3325 */
128'h00000000000000000000000000000000, /* 3326 */
128'h00000000000000000000000000000000, /* 3327 */
128'h00000000000000000000000000000000, /* 3328 */
128'h00000000000000000000000000000000, /* 3329 */
128'h00000000000000000000000000000000, /* 3330 */
128'h00000000000000000000000000000000, /* 3331 */
128'h00000000000000000000000000000000, /* 3332 */
128'h00000000000000000000000000000000, /* 3333 */
128'h00000000000000000000000000000000, /* 3334 */
128'h00000000000000000000000000000000, /* 3335 */
128'h00000000000000000000000000000000, /* 3336 */
128'h00000000000000000000000000000000, /* 3337 */
128'h00000000000000000000000000000000, /* 3338 */
128'h00000000000000000000000000000000, /* 3339 */
128'h00000000000000000000000000000000, /* 3340 */
128'h00000000000000000000000000000000, /* 3341 */
128'h00000000000000000000000000000000, /* 3342 */
128'h00000000000000000000000000000000, /* 3343 */
128'h00000000000000000000000000000000, /* 3344 */
128'h00000000000000000000000000000000, /* 3345 */
128'h00000000000000000000000000000000, /* 3346 */
128'h00000000000000000000000000000000, /* 3347 */
128'h00000000000000000000000000000000, /* 3348 */
128'h00000000000000000000000000000000, /* 3349 */
128'h00000000000000000000000000000000, /* 3350 */
128'h00000000000000000000000000000000, /* 3351 */
128'h00000000000000000000000000000000, /* 3352 */
128'h00000000000000000000000000000000, /* 3353 */
128'h00000000000000000000000000000000, /* 3354 */
128'h00000000000000000000000000000000, /* 3355 */
128'h00000000000000000000000000000000, /* 3356 */
128'h00000000000000000000000000000000, /* 3357 */
128'h00000000000000000000000000000000, /* 3358 */
128'h00000000000000000000000000000000, /* 3359 */
128'h00000000000000000000000000000000, /* 3360 */
128'h00000000000000000000000000000000, /* 3361 */
128'h00000000000000000000000000000000, /* 3362 */
128'h00000000000000000000000000000000, /* 3363 */
128'h00000000000000000000000000000000, /* 3364 */
128'h00000000000000000000000000000000, /* 3365 */
128'h00000000000000000000000000000000, /* 3366 */
128'h00000000000000000000000000000000, /* 3367 */
128'h00000000000000000000000000000000, /* 3368 */
128'h00000000000000000000000000000000, /* 3369 */
128'h00000000000000000000000000000000, /* 3370 */
128'h00000000000000000000000000000000, /* 3371 */
128'h00000000000000000000000000000000, /* 3372 */
128'h00000000000000000000000000000000, /* 3373 */
128'h00000000000000000000000000000000, /* 3374 */
128'h00000000000000000000000000000000, /* 3375 */
128'h00000000000000000000000000000000, /* 3376 */
128'h00000000000000000000000000000000, /* 3377 */
128'h00000000000000000000000000000000, /* 3378 */
128'h00000000000000000000000000000000, /* 3379 */
128'h00000000000000000000000000000000, /* 3380 */
128'h00000000000000000000000000000000, /* 3381 */
128'h00000000000000000000000000000000, /* 3382 */
128'h00000000000000000000000000000000, /* 3383 */
128'h00000000000000000000000000000000, /* 3384 */
128'h00000000000000000000000000000000, /* 3385 */
128'h00000000000000000000000000000000, /* 3386 */
128'h00000000000000000000000000000000, /* 3387 */
128'h00000000000000000000000000000000, /* 3388 */
128'h00000000000000000000000000000000, /* 3389 */
128'h00000000000000000000000000000000, /* 3390 */
128'h00000000000000000000000000000000, /* 3391 */
128'h00000000000000000000000000000000, /* 3392 */
128'h00000000000000000000000000000000, /* 3393 */
128'h00000000000000000000000000000000, /* 3394 */
128'h00000000000000000000000000000000, /* 3395 */
128'h00000000000000000000000000000000, /* 3396 */
128'h00000000000000000000000000000000, /* 3397 */
128'h00000000000000000000000000000000, /* 3398 */
128'h00000000000000000000000000000000, /* 3399 */
128'h00000000000000000000000000000000, /* 3400 */
128'h00000000000000000000000000000000, /* 3401 */
128'h00000000000000000000000000000000, /* 3402 */
128'h00000000000000000000000000000000, /* 3403 */
128'h00000000000000000000000000000000, /* 3404 */
128'h00000000000000000000000000000000, /* 3405 */
128'h00000000000000000000000000000000, /* 3406 */
128'h00000000000000000000000000000000, /* 3407 */
128'h00000000000000000000000000000000, /* 3408 */
128'h00000000000000000000000000000000, /* 3409 */
128'h00000000000000000000000000000000, /* 3410 */
128'h00000000000000000000000000000000, /* 3411 */
128'h00000000000000000000000000000000, /* 3412 */
128'h00000000000000000000000000000000, /* 3413 */
128'h00000000000000000000000000000000, /* 3414 */
128'h00000000000000000000000000000000, /* 3415 */
128'h00000000000000000000000000000000, /* 3416 */
128'h00000000000000000000000000000000, /* 3417 */
128'h00000000000000000000000000000000, /* 3418 */
128'h00000000000000000000000000000000, /* 3419 */
128'h00000000000000000000000000000000, /* 3420 */
128'h00000000000000000000000000000000, /* 3421 */
128'h00000000000000000000000000000000, /* 3422 */
128'h00000000000000000000000000000000, /* 3423 */
128'h00000000000000000000000000000000, /* 3424 */
128'h00000000000000000000000000000000, /* 3425 */
128'h00000000000000000000000000000000, /* 3426 */
128'h00000000000000000000000000000000, /* 3427 */
128'h00000000000000000000000000000000, /* 3428 */
128'h00000000000000000000000000000000, /* 3429 */
128'h00000000000000000000000000000000, /* 3430 */
128'h00000000000000000000000000000000, /* 3431 */
128'h00000000000000000000000000000000, /* 3432 */
128'h00000000000000000000000000000000, /* 3433 */
128'h00000000000000000000000000000000, /* 3434 */
128'h00000000000000000000000000000000, /* 3435 */
128'h00000000000000000000000000000000, /* 3436 */
128'h00000000000000000000000000000000, /* 3437 */
128'h00000000000000000000000000000000, /* 3438 */
128'h00000000000000000000000000000000, /* 3439 */
128'h00000000000000000000000000000000, /* 3440 */
128'h00000000000000000000000000000000, /* 3441 */
128'h00000000000000000000000000000000, /* 3442 */
128'h00000000000000000000000000000000, /* 3443 */
128'h00000000000000000000000000000000, /* 3444 */
128'h00000000000000000000000000000000, /* 3445 */
128'h00000000000000000000000000000000, /* 3446 */
128'h00000000000000000000000000000000, /* 3447 */
128'h00000000000000000000000000000000, /* 3448 */
128'h00000000000000000000000000000000, /* 3449 */
128'h00000000000000000000000000000000, /* 3450 */
128'h00000000000000000000000000000000, /* 3451 */
128'h00000000000000000000000000000000, /* 3452 */
128'h00000000000000000000000000000000, /* 3453 */
128'h00000000000000000000000000000000, /* 3454 */
128'h00000000000000000000000000000000, /* 3455 */
128'h00000000000000000000000000000000, /* 3456 */
128'h00000000000000000000000000000000, /* 3457 */
128'h00000000000000000000000000000000, /* 3458 */
128'h00000000000000000000000000000000, /* 3459 */
128'h00000000000000000000000000000000, /* 3460 */
128'h00000000000000000000000000000000, /* 3461 */
128'h00000000000000000000000000000000, /* 3462 */
128'h00000000000000000000000000000000, /* 3463 */
128'h00000000000000000000000000000000, /* 3464 */
128'h00000000000000000000000000000000, /* 3465 */
128'h00000000000000000000000000000000, /* 3466 */
128'h00000000000000000000000000000000, /* 3467 */
128'h00000000000000000000000000000000, /* 3468 */
128'h00000000000000000000000000000000, /* 3469 */
128'h00000000000000000000000000000000, /* 3470 */
128'h00000000000000000000000000000000, /* 3471 */
128'h00000000000000000000000000000000, /* 3472 */
128'h00000000000000000000000000000000, /* 3473 */
128'h00000000000000000000000000000000, /* 3474 */
128'h00000000000000000000000000000000, /* 3475 */
128'h00000000000000000000000000000000, /* 3476 */
128'h00000000000000000000000000000000, /* 3477 */
128'h00000000000000000000000000000000, /* 3478 */
128'h00000000000000000000000000000000, /* 3479 */
128'h00000000000000000000000000000000, /* 3480 */
128'h00000000000000000000000000000000, /* 3481 */
128'h00000000000000000000000000000000, /* 3482 */
128'h00000000000000000000000000000000, /* 3483 */
128'h00000000000000000000000000000000, /* 3484 */
128'h00000000000000000000000000000000, /* 3485 */
128'h00000000000000000000000000000000, /* 3486 */
128'h00000000000000000000000000000000, /* 3487 */
128'h00000000000000000000000000000000, /* 3488 */
128'h00000000000000000000000000000000, /* 3489 */
128'h00000000000000000000000000000000, /* 3490 */
128'h00000000000000000000000000000000, /* 3491 */
128'h00000000000000000000000000000000, /* 3492 */
128'h00000000000000000000000000000000, /* 3493 */
128'h00000000000000000000000000000000, /* 3494 */
128'h00000000000000000000000000000000, /* 3495 */
128'h00000000000000000000000000000000, /* 3496 */
128'h00000000000000000000000000000000, /* 3497 */
128'h00000000000000000000000000000000, /* 3498 */
128'h00000000000000000000000000000000, /* 3499 */
128'h00000000000000000000000000000000, /* 3500 */
128'h00000000000000000000000000000000, /* 3501 */
128'h00000000000000000000000000000000, /* 3502 */
128'h00000000000000000000000000000000, /* 3503 */
128'h00000000000000000000000000000000, /* 3504 */
128'h00000000000000000000000000000000, /* 3505 */
128'h00000000000000000000000000000000, /* 3506 */
128'h00000000000000000000000000000000, /* 3507 */
128'h00000000000000000000000000000000, /* 3508 */
128'h00000000000000000000000000000000, /* 3509 */
128'h00000000000000000000000000000000, /* 3510 */
128'h00000000000000000000000000000000, /* 3511 */
128'h00000000000000000000000000000000, /* 3512 */
128'h00000000000000000000000000000000, /* 3513 */
128'h00000000000000000000000000000000, /* 3514 */
128'h00000000000000000000000000000000, /* 3515 */
128'h00000000000000000000000000000000, /* 3516 */
128'h00000000000000000000000000000000, /* 3517 */
128'h00000000000000000000000000000000, /* 3518 */
128'h00000000000000000000000000000000, /* 3519 */
128'h00000000000000000000000000000000, /* 3520 */
128'h00000000000000000000000000000000, /* 3521 */
128'h00000000000000000000000000000000, /* 3522 */
128'h00000000000000000000000000000000, /* 3523 */
128'h00000000000000000000000000000000, /* 3524 */
128'h00000000000000000000000000000000, /* 3525 */
128'h00000000000000000000000000000000, /* 3526 */
128'h00000000000000000000000000000000, /* 3527 */
128'h00000000000000000000000000000000, /* 3528 */
128'h00000000000000000000000000000000, /* 3529 */
128'h00000000000000000000000000000000, /* 3530 */
128'h00000000000000000000000000000000, /* 3531 */
128'h00000000000000000000000000000000, /* 3532 */
128'h00000000000000000000000000000000, /* 3533 */
128'h00000000000000000000000000000000, /* 3534 */
128'h00000000000000000000000000000000, /* 3535 */
128'h00000000000000000000000000000000, /* 3536 */
128'h00000000000000000000000000000000, /* 3537 */
128'h00000000000000000000000000000000, /* 3538 */
128'h00000000000000000000000000000000, /* 3539 */
128'h00000000000000000000000000000000, /* 3540 */
128'h00000000000000000000000000000000, /* 3541 */
128'h00000000000000000000000000000000, /* 3542 */
128'h00000000000000000000000000000000, /* 3543 */
128'h00000000000000000000000000000000, /* 3544 */
128'h00000000000000000000000000000000, /* 3545 */
128'h00000000000000000000000000000000, /* 3546 */
128'h00000000000000000000000000000000, /* 3547 */
128'h00000000000000000000000000000000, /* 3548 */
128'h00000000000000000000000000000000, /* 3549 */
128'h00000000000000000000000000000000, /* 3550 */
128'h00000000000000000000000000000000, /* 3551 */
128'h00000000000000000000000000000000, /* 3552 */
128'h00000000000000000000000000000000, /* 3553 */
128'h00000000000000000000000000000000, /* 3554 */
128'h00000000000000000000000000000000, /* 3555 */
128'h00000000000000000000000000000000, /* 3556 */
128'h00000000000000000000000000000000, /* 3557 */
128'h00000000000000000000000000000000, /* 3558 */
128'h00000000000000000000000000000000, /* 3559 */
128'h00000000000000000000000000000000, /* 3560 */
128'h00000000000000000000000000000000, /* 3561 */
128'h00000000000000000000000000000000, /* 3562 */
128'h00000000000000000000000000000000, /* 3563 */
128'h00000000000000000000000000000000, /* 3564 */
128'h00000000000000000000000000000000, /* 3565 */
128'h00000000000000000000000000000000, /* 3566 */
128'h00000000000000000000000000000000, /* 3567 */
128'h00000000000000000000000000000000, /* 3568 */
128'h00000000000000000000000000000000, /* 3569 */
128'h00000000000000000000000000000000, /* 3570 */
128'h00000000000000000000000000000000, /* 3571 */
128'h00000000000000000000000000000000, /* 3572 */
128'h00000000000000000000000000000000, /* 3573 */
128'h00000000000000000000000000000000, /* 3574 */
128'h00000000000000000000000000000000, /* 3575 */
128'h00000000000000000000000000000000, /* 3576 */
128'h00000000000000000000000000000000, /* 3577 */
128'h00000000000000000000000000000000, /* 3578 */
128'h00000000000000000000000000000000, /* 3579 */
128'h00000000000000000000000000000000, /* 3580 */
128'h00000000000000000000000000000000, /* 3581 */
128'h00000000000000000000000000000000, /* 3582 */
128'h00000000000000000000000000000000, /* 3583 */
128'h00000000000000000000000000000000, /* 3584 */
128'h00000000000000000000000000000000, /* 3585 */
128'h00000000000000000000000000000000, /* 3586 */
128'h00000000000000000000000000000000, /* 3587 */
128'h00000000000000000000000000000000, /* 3588 */
128'h00000000000000000000000000000000, /* 3589 */
128'h00000000000000000000000000000000, /* 3590 */
128'h00000000000000000000000000000000, /* 3591 */
128'h00000000000000000000000000000000, /* 3592 */
128'h00000000000000000000000000000000, /* 3593 */
128'h00000000000000000000000000000000, /* 3594 */
128'h00000000000000000000000000000000, /* 3595 */
128'h00000000000000000000000000000000, /* 3596 */
128'h00000000000000000000000000000000, /* 3597 */
128'h00000000000000000000000000000000, /* 3598 */
128'h00000000000000000000000000000000, /* 3599 */
128'h00000000000000000000000000000000, /* 3600 */
128'h00000000000000000000000000000000, /* 3601 */
128'h00000000000000000000000000000000, /* 3602 */
128'h00000000000000000000000000000000, /* 3603 */
128'h00000000000000000000000000000000, /* 3604 */
128'h00000000000000000000000000000000, /* 3605 */
128'h00000000000000000000000000000000, /* 3606 */
128'h00000000000000000000000000000000, /* 3607 */
128'h00000000000000000000000000000000, /* 3608 */
128'h00000000000000000000000000000000, /* 3609 */
128'h00000000000000000000000000000000, /* 3610 */
128'h00000000000000000000000000000000, /* 3611 */
128'h00000000000000000000000000000000, /* 3612 */
128'h00000000000000000000000000000000, /* 3613 */
128'h00000000000000000000000000000000, /* 3614 */
128'h00000000000000000000000000000000, /* 3615 */
128'h00000000000000000000000000000000, /* 3616 */
128'h00000000000000000000000000000000, /* 3617 */
128'h00000000000000000000000000000000, /* 3618 */
128'h00000000000000000000000000000000, /* 3619 */
128'h00000000000000000000000000000000, /* 3620 */
128'h00000000000000000000000000000000, /* 3621 */
128'h00000000000000000000000000000000, /* 3622 */
128'h00000000000000000000000000000000, /* 3623 */
128'h00000000000000000000000000000000, /* 3624 */
128'h00000000000000000000000000000000, /* 3625 */
128'h00000000000000000000000000000000, /* 3626 */
128'h00000000000000000000000000000000, /* 3627 */
128'h00000000000000000000000000000000, /* 3628 */
128'h00000000000000000000000000000000, /* 3629 */
128'h00000000000000000000000000000000, /* 3630 */
128'h00000000000000000000000000000000, /* 3631 */
128'h00000000000000000000000000000000, /* 3632 */
128'h00000000000000000000000000000000, /* 3633 */
128'h00000000000000000000000000000000, /* 3634 */
128'h00000000000000000000000000000000, /* 3635 */
128'h00000000000000000000000000000000, /* 3636 */
128'h00000000000000000000000000000000, /* 3637 */
128'h00000000000000000000000000000000, /* 3638 */
128'h00000000000000000000000000000000, /* 3639 */
128'h00000000000000000000000000000000, /* 3640 */
128'h00000000000000000000000000000000, /* 3641 */
128'h00000000000000000000000000000000, /* 3642 */
128'h00000000000000000000000000000000, /* 3643 */
128'h00000000000000000000000000000000, /* 3644 */
128'h00000000000000000000000000000000, /* 3645 */
128'h00000000000000000000000000000000, /* 3646 */
128'h00000000000000000000000000000000, /* 3647 */
128'h00000000000000000000000000000000, /* 3648 */
128'h00000000000000000000000000000000, /* 3649 */
128'h00000000000000000000000000000000, /* 3650 */
128'h00000000000000000000000000000000, /* 3651 */
128'h00000000000000000000000000000000, /* 3652 */
128'h00000000000000000000000000000000, /* 3653 */
128'h00000000000000000000000000000000, /* 3654 */
128'h00000000000000000000000000000000, /* 3655 */
128'h00000000000000000000000000000000, /* 3656 */
128'h00000000000000000000000000000000, /* 3657 */
128'h00000000000000000000000000000000, /* 3658 */
128'h00000000000000000000000000000000, /* 3659 */
128'h00000000000000000000000000000000, /* 3660 */
128'h00000000000000000000000000000000, /* 3661 */
128'h00000000000000000000000000000000, /* 3662 */
128'h00000000000000000000000000000000, /* 3663 */
128'h00000000000000000000000000000000, /* 3664 */
128'h00000000000000000000000000000000, /* 3665 */
128'h00000000000000000000000000000000, /* 3666 */
128'h00000000000000000000000000000000, /* 3667 */
128'h00000000000000000000000000000000, /* 3668 */
128'h00000000000000000000000000000000, /* 3669 */
128'h00000000000000000000000000000000, /* 3670 */
128'h00000000000000000000000000000000, /* 3671 */
128'h00000000000000000000000000000000, /* 3672 */
128'h00000000000000000000000000000000, /* 3673 */
128'h00000000000000000000000000000000, /* 3674 */
128'h00000000000000000000000000000000, /* 3675 */
128'h00000000000000000000000000000000, /* 3676 */
128'h00000000000000000000000000000000, /* 3677 */
128'h00000000000000000000000000000000, /* 3678 */
128'h00000000000000000000000000000000, /* 3679 */
128'h00000000000000000000000000000000, /* 3680 */
128'h00000000000000000000000000000000, /* 3681 */
128'h00000000000000000000000000000000, /* 3682 */
128'h00000000000000000000000000000000, /* 3683 */
128'h00000000000000000000000000000000, /* 3684 */
128'h00000000000000000000000000000000, /* 3685 */
128'h00000000000000000000000000000000, /* 3686 */
128'h00000000000000000000000000000000, /* 3687 */
128'h00000000000000000000000000000000, /* 3688 */
128'h00000000000000000000000000000000, /* 3689 */
128'h00000000000000000000000000000000, /* 3690 */
128'h00000000000000000000000000000000, /* 3691 */
128'h00000000000000000000000000000000, /* 3692 */
128'h00000000000000000000000000000000, /* 3693 */
128'h00000000000000000000000000000000, /* 3694 */
128'h00000000000000000000000000000000, /* 3695 */
128'h00000000000000000000000000000000, /* 3696 */
128'h00000000000000000000000000000000, /* 3697 */
128'h00000000000000000000000000000000, /* 3698 */
128'h00000000000000000000000000000000, /* 3699 */
128'h00000000000000000000000000000000, /* 3700 */
128'h00000000000000000000000000000000, /* 3701 */
128'h00000000000000000000000000000000, /* 3702 */
128'h00000000000000000000000000000000, /* 3703 */
128'h00000000000000000000000000000000, /* 3704 */
128'h00000000000000000000000000000000, /* 3705 */
128'h00000000000000000000000000000000, /* 3706 */
128'h00000000000000000000000000000000, /* 3707 */
128'h00000000000000000000000000000000, /* 3708 */
128'h00000000000000000000000000000000, /* 3709 */
128'h00000000000000000000000000000000, /* 3710 */
128'h00000000000000000000000000000000, /* 3711 */
128'h00000000000000000000000000000000, /* 3712 */
128'h00000000000000000000000000000000, /* 3713 */
128'h00000000000000000000000000000000, /* 3714 */
128'h00000000000000000000000000000000, /* 3715 */
128'h00000000000000000000000000000000, /* 3716 */
128'h00000000000000000000000000000000, /* 3717 */
128'h00000000000000000000000000000000, /* 3718 */
128'h00000000000000000000000000000000, /* 3719 */
128'h00000000000000000000000000000000, /* 3720 */
128'h00000000000000000000000000000000, /* 3721 */
128'h00000000000000000000000000000000, /* 3722 */
128'h00000000000000000000000000000000, /* 3723 */
128'h00000000000000000000000000000000, /* 3724 */
128'h00000000000000000000000000000000, /* 3725 */
128'h00000000000000000000000000000000, /* 3726 */
128'h00000000000000000000000000000000, /* 3727 */
128'h00000000000000000000000000000000, /* 3728 */
128'h00000000000000000000000000000000, /* 3729 */
128'h00000000000000000000000000000000, /* 3730 */
128'h00000000000000000000000000000000, /* 3731 */
128'h00000000000000000000000000000000, /* 3732 */
128'h00000000000000000000000000000000, /* 3733 */
128'h00000000000000000000000000000000, /* 3734 */
128'h00000000000000000000000000000000, /* 3735 */
128'h00000000000000000000000000000000, /* 3736 */
128'h00000000000000000000000000000000, /* 3737 */
128'h00000000000000000000000000000000, /* 3738 */
128'h00000000000000000000000000000000, /* 3739 */
128'h00000000000000000000000000000000, /* 3740 */
128'h00000000000000000000000000000000, /* 3741 */
128'h00000000000000000000000000000000, /* 3742 */
128'h00000000000000000000000000000000, /* 3743 */
128'h00000000000000000000000000000000, /* 3744 */
128'h00000000000000000000000000000000, /* 3745 */
128'h00000000000000000000000000000000, /* 3746 */
128'h00000000000000000000000000000000, /* 3747 */
128'h00000000000000000000000000000000, /* 3748 */
128'h00000000000000000000000000000000, /* 3749 */
128'h00000000000000000000000000000000, /* 3750 */
128'h00000000000000000000000000000000, /* 3751 */
128'h00000000000000000000000000000000, /* 3752 */
128'h00000000000000000000000000000000, /* 3753 */
128'h00000000000000000000000000000000, /* 3754 */
128'h00000000000000000000000000000000, /* 3755 */
128'h00000000000000000000000000000000, /* 3756 */
128'h00000000000000000000000000000000, /* 3757 */
128'h00000000000000000000000000000000, /* 3758 */
128'h00000000000000000000000000000000, /* 3759 */
128'h00000000000000000000000000000000, /* 3760 */
128'h00000000000000000000000000000000, /* 3761 */
128'h00000000000000000000000000000000, /* 3762 */
128'h00000000000000000000000000000000, /* 3763 */
128'h00000000000000000000000000000000, /* 3764 */
128'h00000000000000000000000000000000, /* 3765 */
128'h00000000000000000000000000000000, /* 3766 */
128'h00000000000000000000000000000000, /* 3767 */
128'h00000000000000000000000000000000, /* 3768 */
128'h00000000000000000000000000000000, /* 3769 */
128'h00000000000000000000000000000000, /* 3770 */
128'h00000000000000000000000000000000, /* 3771 */
128'h00000000000000000000000000000000, /* 3772 */
128'h00000000000000000000000000000000, /* 3773 */
128'h00000000000000000000000000000000, /* 3774 */
128'h00000000000000000000000000000000, /* 3775 */
128'h00000000000000000000000000000000, /* 3776 */
128'h00000000000000000000000000000000, /* 3777 */
128'h00000000000000000000000000000000, /* 3778 */
128'h00000000000000000000000000000000, /* 3779 */
128'h00000000000000000000000000000000, /* 3780 */
128'h00000000000000000000000000000000, /* 3781 */
128'h00000000000000000000000000000000, /* 3782 */
128'h00000000000000000000000000000000, /* 3783 */
128'h00000000000000000000000000000000, /* 3784 */
128'h00000000000000000000000000000000, /* 3785 */
128'h00000000000000000000000000000000, /* 3786 */
128'h00000000000000000000000000000000, /* 3787 */
128'h00000000000000000000000000000000, /* 3788 */
128'h00000000000000000000000000000000, /* 3789 */
128'h00000000000000000000000000000000, /* 3790 */
128'h00000000000000000000000000000000, /* 3791 */
128'h00000000000000000000000000000000, /* 3792 */
128'h00000000000000000000000000000000, /* 3793 */
128'h00000000000000000000000000000000, /* 3794 */
128'h00000000000000000000000000000000, /* 3795 */
128'h00000000000000000000000000000000, /* 3796 */
128'h00000000000000000000000000000000, /* 3797 */
128'h00000000000000000000000000000000, /* 3798 */
128'h00000000000000000000000000000000, /* 3799 */
128'h00000000000000000000000000000000, /* 3800 */
128'h00000000000000000000000000000000, /* 3801 */
128'h00000000000000000000000000000000, /* 3802 */
128'h00000000000000000000000000000000, /* 3803 */
128'h00000000000000000000000000000000, /* 3804 */
128'h00000000000000000000000000000000, /* 3805 */
128'h00000000000000000000000000000000, /* 3806 */
128'h00000000000000000000000000000000, /* 3807 */
128'h00000000000000000000000000000000, /* 3808 */
128'h00000000000000000000000000000000, /* 3809 */
128'h00000000000000000000000000000000, /* 3810 */
128'h00000000000000000000000000000000, /* 3811 */
128'h00000000000000000000000000000000, /* 3812 */
128'h00000000000000000000000000000000, /* 3813 */
128'h00000000000000000000000000000000, /* 3814 */
128'h00000000000000000000000000000000, /* 3815 */
128'h00000000000000000000000000000000, /* 3816 */
128'h00000000000000000000000000000000, /* 3817 */
128'h00000000000000000000000000000000, /* 3818 */
128'h00000000000000000000000000000000, /* 3819 */
128'h00000000000000000000000000000000, /* 3820 */
128'h00000000000000000000000000000000, /* 3821 */
128'h00000000000000000000000000000000, /* 3822 */
128'h00000000000000000000000000000000, /* 3823 */
128'h00000000000000000000000000000000, /* 3824 */
128'h00000000000000000000000000000000, /* 3825 */
128'h00000000000000000000000000000000, /* 3826 */
128'h00000000000000000000000000000000, /* 3827 */
128'h00000000000000000000000000000000, /* 3828 */
128'h00000000000000000000000000000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00000000000000000000000000000000, /* 3840 */
128'h00000000000000000000000000000000, /* 3841 */
128'h00000000000000000000000000000000, /* 3842 */
128'h00000000000000000000000000000000, /* 3843 */
128'h00000000000000000000000000000000, /* 3844 */
128'h00000000000000000000000000000000, /* 3845 */
128'h00000000000000000000000000000000, /* 3846 */
128'h00000000000000000000000000000000, /* 3847 */
128'h00000000000000000000000000000000, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule

