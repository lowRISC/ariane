/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'h00004617fec58593000005970d249263, /*    1 */
128'h010696937ff6869b000086b7de460613, /*    2 */
128'h0085b70300e6b0230005b70300d007b3, /*    3 */
128'h0185b70300e6b8230105b70300e6b423, /*    4 */
128'hfcc5cce3020686930205859300e6bc23, /*    5 */
128'h40b787b300d787b30147879300000797, /*    6 */
128'h305790730b8787930000079700078067, /*    7 */
128'h00004597010111137ff1011b00008137, /*    8 */
128'h0005b023fb06061300004617d7458593, /*    9 */
128'h020585930005bc230005b8230005b423, /*   10 */
128'h00100913020004b7003020effec5c6e3, /*   11 */
128'h4009091b02000937004484930124a023, /*   12 */
128'h008979133440297310500073ff24c6e3, /*   13 */
128'h00291913f1402973020004b7fe090ae3, /*   14 */
128'hfe091ee30004a9030009202300990933, /*   15 */
128'hff24c6e34009091b0200093700448493, /*   16 */
128'h000084b792c5859300003597f1402573, /*   17 */
128'h342022f300048067010494937ff4849b, /*   18 */
128'h00000000ffdff06f1050007334102373, /*   19 */
128'h00000000000000000000000000000000, /*   20 */
128'h00000000000000000000000000000000, /*   21 */
128'h00000000000000000000000000000000, /*   22 */
128'h00000000000000000000000000000000, /*   23 */
128'h00000000000000000000000000000000, /*   24 */
128'h00000000000000000000000000000000, /*   25 */
128'h00000000000000000000000000000000, /*   26 */
128'h00000000000000000000000000000000, /*   27 */
128'h00000000000000000000000000000000, /*   28 */
128'h00000000000000000000000000000000, /*   29 */
128'h00000000000000000000000000000000, /*   30 */
128'h00000000000000000000000000000000, /*   31 */
128'h00b500230640006f4605051300003517, /*   32 */
128'h0147c503100007b78082000545038082, /*   33 */
128'hf7930147478310000737808202057513, /*   34 */
128'h8223100007b7808200a70023dfe50207, /*   35 */
128'h00e78023476d00e78623f80007130007, /*   36 */
128'h8423fc70071300e78623470d00078223, /*   37 */
128'he0221141808200e788230200071300e7, /*   38 */
128'h0141640260a2e50900044503842ae406, /*   39 */
128'h879300002797b7f50405fa5ff0ef8082, /*   40 */
128'h0007470397aa973e811100f577136767, /*   41 */
128'h1101808200f5802300e580a30007c783, /*   42 */
128'h4503fd1ff0efec068121842a002ce822, /*   43 */
128'h002cf5dff0ef00914503f65ff0ef0081, /*   44 */
128'hf4bff0ef00814503fb7ff0ef0ff47513, /*   45 */
128'h80826105644260e2f43ff0ef00914503, /*   46 */
128'h54e14461892af406e84aec26f0227179, /*   47 */
128'h4503f81ff0ef0ff57513002c0089553b, /*   48 */
128'hf0bff0ef00914503f13ff0ef34610081, /*   49 */
128'h80826145694264e2740270a2fe9410e3, /*   50 */
128'h03800413892af406e84aec26f0227179, /*   51 */
128'hf3fff0ef0ff57513002c0089553354e1, /*   52 */
128'hf0ef00914503ed1ff0ef346100814503, /*   53 */
128'h6145694264e2740270a2fe9410e3ec9f, /*   54 */
128'h00814503f13ff0efec06002c11018082, /*   55 */
128'h610560e2e9fff0ef00914503ea7ff0ef, /*   56 */
128'h47178082400005378082057e45058082, /*   57 */
128'h869300756513157d631ccea707130000, /*   58 */
128'h057e450597aa20000537e30895360017, /*   59 */
128'h862a0ce507638207871367858082953e, /*   60 */
128'h2a050513000035178087871308a74463, /*   61 */
128'h000035178006079b04c7496306e60b63, /*   62 */
128'h0000351787f787936785c3ad27c50513, /*   63 */
128'h11417c07879b77fd04c7c9632fc50513, /*   64 */
128'h0513000045172ee58593000035979e3d, /*   65 */
128'h05130000451760a2696010efe4069e65, /*   66 */
128'h05130000351781078713808201419d65, /*   67 */
128'h0513000035178187879300e60a6324e5, /*   68 */
128'h00003517830787138082faf612e324e5, /*   69 */
128'h8287879300c74963fee609e326c50513, /*   70 */
128'h351783878713bfe92485051300003517, /*   71 */
128'h351784078793fce608e325a505130000, /*   72 */
128'h2105051300003517bf7525a505130000, /*   73 */
128'h440184aaf406e84aec26f02271798082, /*   74 */
128'h0104551302f04463409907bb00a5893b, /*   75 */
128'h740270a2952201045513942a90411442, /*   76 */
128'h808261459141694264e21542fff54513, /*   77 */
128'h048900c157835f9010ef0068460985a6, /*   78 */
128'h17c200f117238fd90087979b0087d71b, /*   79 */
128'hfc26e486e0a26785715dbf45943e93c1, /*   80 */
128'h67a13cf50463842e80678793f44ef84a, /*   81 */
128'h440799638005079b0af50e636dd78793, /*   82 */
128'h006409135a7010ef4611082884b205e9, /*   83 */
128'h593010efb3c5051300004517461985ca, /*   84 */
128'h08b7e76332f5886302e0079301744583, /*   85 */
128'h1af58263479104b7e5631cf5816347b1, /*   86 */
128'h00003517478910f58463478502b7e363, /*   87 */
128'h330505130000351702f5836319450513, /*   88 */
128'h351747a118f581634799a41554e010ef, /*   89 */
128'ha429534010effef591e319a505130000, /*   90 */
128'h16f5896347c500b7ed632cf5816347f5, /*   91 */
128'hbf6dfef580e31b6505130000351747d9, /*   92 */
128'hfaf596e3029007932af5856302100793, /*   93 */
128'h816306200793b7c91d05051300003517, /*   94 */
128'hef632af581630330079304b7e2632cf5, /*   95 */
128'h35170320079328f5866302f0079300b7, /*   96 */
128'h05c00793b7bdf8f58ae31d2505130000, /*   97 */
128'h1e8505130000351705e0079328f58363, /*   98 */
128'hef6328f5856308400793bf91f6f58de3, /*   99 */
128'h351706c0079326f58a630670079300b7, /*  100 */
128'h08900793b73df4f58ae31fa505130000, /*  101 */
128'h0880079326f588630ff0079326f58763, /*  102 */
128'h5703b73d2045051300003517f0f59ce3, /*  103 */
128'h8993000049979ee7d7830000479701e4, /*  104 */
128'hd783000047970204570312f713639e69, /*  105 */
128'h433010ef852285ca461910f71b639d87, /*  106 */
128'h423010ef854a9a658593000045974619, /*  107 */
128'h00f41f23020412230204012301a45783, /*  108 */
128'h02f4102302240513fde4859b01c45783, /*  109 */
128'h00f41e230029d78300f41d230009d783, /*  110 */
128'h00a11e238d5d05220085579bdb3ff0ef, /*  111 */
128'ha06d7bc000ef450185a2862602a41223, /*  112 */
128'h051300003517bd490085051300003517, /*  113 */
128'h4783bdbd0245051300003517b5610165, /*  114 */
128'h0e230254478300f10ea3026447030244, /*  115 */
128'h27810274470300e10ea301c1178300f1, /*  116 */
128'h00e10ea301c119030224470300e10e23, /*  117 */
128'h01c156830450071300e10e2302344703, /*  118 */
128'h461947e292d794230000479704e79b63, /*  119 */
128'h90850513000045179005859300004597, /*  120 */
128'h4762345010efe43690f7242300004717, /*  121 */
128'h0593ff89061b8de787930000479766a2, /*  122 */
128'h794274e2640660a6096020ef450102a4, /*  123 */
128'h47e204e69463043007138082616179a2, /*  124 */
128'h8cc78793000047978cf7242300004717, /*  125 */
128'hf7e9439c8bc7879300004797c799439c, /*  126 */
128'h8ac60613000046178b06869300004697, /*  127 */
128'h762000ef02a405138505859300004597, /*  128 */
128'h05130000351702e798634d200713b765, /*  129 */
128'h351769b000ef852285a62bc010eff3e5, /*  130 */
128'h02a4051385ca2a8010eff3a505130000, /*  131 */
128'h5703f6e787e35fe00713bf95685000ef, /*  132 */
128'h0de302045703f6f701e317fd67c101e4, /*  133 */
128'h10ef086880c58593000045974611f4f7, /*  134 */
128'h3517b33df145051300003517b7992710, /*  135 */
128'hf305051300003517b315f1a505130000, /*  136 */
128'h00003517bb01f3e5051300003517bb29, /*  137 */
128'hb9f5f5a5051300003517b319f5450513, /*  138 */
128'h051300003517b9cdf785051300003517, /*  139 */
128'h3517b9f9f9c5051300003517b1e5f865, /*  140 */
128'hfd05051300003517b9d1fc2505130000, /*  141 */
128'h349778a7d783000037970265d703b1e9, /*  142 */
128'h37970285d703ecf711e3782484930000, /*  143 */
128'h891320000793eaf719e37747d7830000, /*  144 */
128'h854a85ce461900f59a23016589930205, /*  145 */
128'h854e732585930000359746191bf010ef, /*  146 */
128'h0513722585930000359746191af010ef, /*  147 */
128'h193010ef852285ca461919d010ef0064, /*  148 */
128'h01e4578302f4132302a0061301c45783, /*  149 */
128'h0024d78300f41e230004d78302f41423, /*  150 */
128'h85aab36900f416236080079300f41f23, /*  151 */
128'hbba54601156010eff585051300003517, /*  152 */
128'h608130239f0101138307b603300017b7, /*  153 */
128'h0034179b66858387b70300f674132601, /*  154 */
128'h97ae300005b79fad8406879b0387f593, /*  155 */
128'hfee7881b2781601134235e913c23639c, /*  156 */
128'h05138a1d09056c63ffc7849b5f200513, /*  157 */
128'hc34927018f71fff7471300c5163b1010, /*  158 */
128'h0084171beb3d43186587071300003717, /*  159 */
128'h45d495ba070e9f318006871b70077613, /*  160 */
128'h0086d69b0106d69b0106969b00d100a3, /*  161 */
128'h6685c6918005069b0001550300d10023, /*  162 */
128'h27850077e79337ed02d51e6380668693, /*  163 */
128'h974285b246814037d79b30000837860a, /*  164 */
128'h3c230621068500083803983a00369813, /*  165 */
128'ha9bff0ef8626fef845e30006881bff06, /*  166 */
128'h3403608130838287b823300017b70405, /*  167 */
128'h11018082610101135f81348385266001, /*  168 */
128'h47812401ec06e42643c0e8220c2007b7, /*  169 */
128'h0206c163033716938304b703300014b7, /*  170 */
128'h07b7024010efe3e5051300003517e799, /*  171 */
128'hf0ef8082610564a2644260e2c3c00c20, /*  172 */
128'h84ae8432ec26f0227179bfc14785ec3f, /*  173 */
128'h10eff406006858e58593000035974611, /*  174 */
128'h47b20007a8035a678793000037977f00, /*  175 */
128'h0000371758c888930000389785a68622, /*  176 */
128'h53850513000035170450069359075703, /*  177 */
128'h8082614564e2740270a285222b1000ef, /*  178 */
128'h171b8082914115428d5d05220085579b, /*  179 */
128'h571bf00686938fd966c10185579b0185, /*  180 */
128'h8d7900ff07370085151b8fd98f750085, /*  181 */
128'hda05051300003517715d808225018d5d, /*  182 */
128'he85aec56f052f44ef84afc26e0a2e486, /*  183 */
128'h371747e14c0786230000379775f000ef, /*  184 */
128'h0c230000371703e007934cf701a30000, /*  185 */
128'h3717578d4af707a30000371747894af7, /*  186 */
128'h0000359707f0079346114af703230000, /*  187 */
128'h371748a4041300003417002849658593, /*  188 */
128'h006885a24609708010ef48f703a30000, /*  189 */
128'h4b09899300003997448145226fe010ef, /*  190 */
128'h971bf00606130100063746b2f4fff0ef, /*  191 */
128'h17b715028f558f710ff6f69382a10086, /*  192 */
128'h80e7b423934180a7b023174291013000, /*  193 */
128'hcf050513000035178087b7038007b703, /*  194 */
128'h07378087b5838007b60382e7b4234721, /*  195 */
128'h8f4d91c115c245ea0a1300003a170080, /*  196 */
128'h3fb747030000371768b000ef80e7b423, /*  197 */
128'h3ed84803000038173f47c78300003797, /*  198 */
128'h3d964603000036173e26c68300003697, /*  199 */
128'hca050513000035173d05c58300003597, /*  200 */
128'h371700989b376a890004478364f000ef, /*  201 */
128'h371730001937001447833af70d230000, /*  202 */
128'h002300003717002447833af705a30000, /*  203 */
128'h478338f70aa300003717003447833af7, /*  204 */
128'h37170054478338f70523000037170044, /*  205 */
128'h37973a079b230000379736f70fa30000, /*  206 */
128'h37973407a923000037973a07a5230000, /*  207 */
128'he4a93807ad23000037973a07a3230000, /*  208 */
128'h680b0493139000ef8522e78d0009a783, /*  209 */
128'h83093783020745630337971383093783, /*  210 */
128'h2783bfc5c59ff0effc075de303379713, /*  211 */
128'h710a8493355010ef4501dff154fd000a, /*  212 */
128'h300017b7b7d914fdb7e9c3fff0efbfc1, /*  213 */
128'h8f75e40616fd1141ff8006b78087b703, /*  214 */
128'hb58382e7b823f0070713670580e7b423, /*  215 */
128'h3517555000efbd650513000035178307, /*  216 */
128'h6709300027f3549000efbf2505130000, /*  217 */
128'h907307fe4785300790738fd988070713, /*  218 */
128'h100f525000efbee50513000035173417, /*  219 */
128'hf713419c8082014160a2302000730000, /*  220 */
128'h06220086571b419cc19c2785c3190017, /*  221 */
128'h0087d7138ed906a20086d71b8e5927a1, /*  222 */
128'h00c510238fd90087979b0ff77713c19c, /*  223 */
128'h419c80820005132300f5122300d51123, /*  224 */
128'h0457879b6785c19c27d1f022f4067179, /*  225 */
128'h77130087d713c632842a419c00f51023, /*  226 */
128'h57fd460900f11a238fd90087979b0ff7, /*  227 */
128'h4609494010ef00f11b23c4360509084c, /*  228 */
128'h462147c1486010ef0044051301610593, /*  229 */
128'h472010efec3e0084051300041323082c, /*  230 */
128'h051300041523006c461100f404a347c5, /*  231 */
128'h10ef01040513002c461145c010ef00c4, /*  232 */
128'hffe7d6030789470187a2014406934500, /*  233 */
128'h9fb9934117424107579bfed79ce39f31, /*  234 */
128'h70a200f41523fff7c7939fb94107d71b, /*  235 */
128'h6394e027879300003797808261457402, /*  236 */
128'he793fff6079b8007bc2397b647216785, /*  237 */
128'h0005071b6805450102e7c7bb27850077, /*  238 */
128'h1713808280c6b82396be678500f74763, /*  239 */
128'h3023973697420008b88300e588b30035, /*  240 */
128'h86220005841be0221141bfe105050117, /*  241 */
128'h640260a28522fa1ff0efe406450185aa, /*  242 */
128'h051984b2842aec26f022717980820141, /*  243 */
128'h4619852266a2398010efe436f4064619, /*  244 */
128'h7402852200f4162347a138c010ef85b6, /*  245 */
128'h0113fadff06f614564e200e4859b70a2, /*  246 */
128'h3423392138233a8130236785737dc501, /*  247 */
128'h3c23394130233931342338913c233a11, /*  248 */
128'h3c233781302337713423376138233751, /*  249 */
128'h747d978a911a3507879335a138233591, /*  250 */
128'h0023ca040b23ce042023d00007b7943e, /*  251 */
128'h5800073797aad0040023f0040023e004, /*  252 */
128'h9e0505130000351785aa00e7ea63892a, /*  253 */
128'h24f71c63478900054703a0012ff000ef, /*  254 */
128'h9abacd848a93970a3507871374fd6785, /*  255 */
128'h8baed0048c13cb848b13970a35078713, /*  256 */
128'h95ca0f0985939c3a9b3a49818a368cb2, /*  257 */
128'h071329890f07c7830015cd03013907b3, /*  258 */
128'h04f76b6326e78a6301a989bb058902a0, /*  259 */
128'h2ae78863470502f7626322e78e634719, /*  260 */
128'h0000351785be22e78663cc848513470d, /*  261 */
128'h22e782634731bf4d27b000efad450513, /*  262 */
128'h8513978a350787936785fee794e3473d, /*  263 */
128'he00d0023256010ef9d22953e866ae004, /*  264 */
128'h071300f76e6322e7806303600713b769, /*  265 */
128'h8513fae798e30350071320e78d630330, /*  266 */
128'h071324e7846303800713aac14605cb64, /*  267 */
128'h8263747d479500614583f8e79ce30ff0, /*  268 */
128'ha7833af59163478936f58563479924f5, /*  269 */
128'h4985978a350a87936a8516079163000c, /*  270 */
128'h013ca023953e461101090593ce440513, /*  271 */
128'h0593ce840513978a350a87931de010ef, /*  272 */
128'h0513000035171c8010ef953e46110149, /*  273 */
128'h350a87931b7000efde0254e25a528be5, /*  274 */
128'h122300f9202357fd993e978acf840913, /*  275 */
128'h46f115231350079300f103a3478d00f9, /*  276 */
128'h460594becb740493c2a6978a350a8793, /*  277 */
128'h03200793176010efc0d246c1051385a6, /*  278 */
128'h95becf040593978a350a879346f106a3, /*  279 */
128'h152010ef4741072346f1051346114a11, /*  280 */
128'h0593978a350a879346f109a303600793, /*  281 */
128'h10ef47410a2347510513461195becf44, /*  282 */
128'h46f10ca347b1051385a6460557fd1300, /*  283 */
128'h10200793116010ef47310d23000103a3, /*  284 */
128'h07930b6010efde3e1ee845810ee00613, /*  285 */
128'h3961051385de4799464136f11d231010, /*  286 */
128'h13232637879377e10ea010ef36f10e23, /*  287 */
128'h350a879346f1142335378793679946f1, /*  288 */
128'h0440061304300693943ecec40413978a, /*  289 */
128'h85a2460156fdba7ff0ef3721051385a2, /*  290 */
128'h0e8885de86ca5672bdbff0ef35e10513, /*  291 */
128'h3a0134033a813083911a6305cf5ff0ef, /*  292 */
128'h38013a03388139833901390339813483, /*  293 */
128'h36013c0336813b8337013b0337813a83, /*  294 */
128'h851380823b01011335013d0335813c83, /*  295 */
128'ha00d953e978a3507879367854611cd04, /*  296 */
128'h953e866af0048513978a350787936785, /*  297 */
128'h85564611bb85f00d002303c010ef9d22, /*  298 */
128'h87936785bfdd855a4611b39d02e010ef, /*  299 */
128'h012010ef4611953ece048513978a3507, /*  300 */
128'h11238fd90087979b0087d71bce045783, /*  301 */
128'h8fd90087979b0087d71bce24578300f4, /*  302 */
128'hcc048513b305cef42023401c00f41023, /*  303 */
128'hd00d00237d7000ef9d228562866ab749, /*  304 */
128'h00fa2023478510079d63000a2783b329, /*  305 */
128'h059346117b6000ef6d05051300002517, /*  306 */
128'h978a3504879364857ab000ef0e880109, /*  307 */
128'h793000ef014905934611953ecb840513, /*  308 */
128'h35014583351146033521468335314703, /*  309 */
128'h35015783776000ef6a05051300002517, /*  310 */
128'hcef71c23000037170091460300a14683, /*  311 */
128'h6a050513000025170081458335215783, /*  312 */
128'h742000ef00b14703cef7112300003717, /*  313 */
128'h018145830191460301a1468301b14703, /*  314 */
128'h01314703726000ef6a05051300002517, /*  315 */
128'h00002517010145830111460301214683, /*  316 */
128'h251755c20101578370a000ef6a450513, /*  317 */
128'h5783c8f71123000037176b2505130000, /*  318 */
128'h87936e4000efc6f71c23000037170121, /*  319 */
128'h05130000251795bee0040593978a3504, /*  320 */
128'h978af0040593350487936cc000ef69e5, /*  321 */
128'hbd196b4000ef696505130000251795be, /*  322 */
128'h2783b5216a6000ef6985051300002517, /*  323 */
128'h0000251700fa20234785e00791e3000a, /*  324 */
128'h690505130000251768a000ef68c50513, /*  325 */
128'h978ad004059335078793678567e000ef, /*  326 */
128'h00002517bf45696505130000251795be, /*  327 */
128'hec86711d737dbb7565a000ef69c50513, /*  328 */
128'h911a89aaf456f852fc4ee0cae4a6e8a2, /*  329 */
128'h632000efca026a856b05051300002517, /*  330 */
128'h57fd94beff840493978a020a8793747d, /*  331 */
128'h439c822787930000379700f49223c09c, /*  332 */
128'h12f11d2313500793c83e4a05fef40913, /*  333 */
128'h07a31a68460585ca993e978a020a8793, /*  334 */
128'h479112f10ea3037007935ed000ef0141, /*  335 */
128'h95beff040593978a020a879312f10f23, /*  336 */
128'h460585ca57fd5c9000ef13f105134611, /*  337 */
128'h000107a31541022314f101a314510513, /*  338 */
128'h00e845810ee006130fc007935af000ef, /*  339 */
128'h85ce04f115231010079354f000efca3e, /*  340 */
128'h583000ef04f106230661051346414799, /*  341 */
128'h35378793679912f11b232637879377e1, /*  342 */
128'h85a2943e1451978a020a879312f11c23, /*  343 */
128'h841ff0ef044006130430069304210513, /*  344 */
128'h4652875ff0ef460156fd02e1051385a2, /*  345 */
128'h60e6911a630598fff0ef85ce86a61008, /*  346 */
128'h61257aa27a4279e2690664a664464501, /*  347 */
128'h5120006f5a4505130000251785aa8082, /*  348 */
128'h81010113e4cee8caeca6f0a2f4867159, /*  349 */
128'hec3ae442893689b2e04605a1051384aa, /*  350 */
128'h81078793101867854eb000efd602e83e, /*  351 */
128'h864a86ba943e7fc404136762747d97ba, /*  352 */
128'h67c26822fb4ff0efd64e0521051385a2, /*  353 */
128'h6882fe4ff0ef03e10513863e86c285a2, /*  354 */
128'h7f0101138fdff0ef86c685a618085632, /*  355 */
128'h8082616569a6694664e67406450170a6, /*  356 */
128'h47830045480300554883e222e606716d, /*  357 */
128'h842a0005460300154683002547030035, /*  358 */
128'h50850513000025175085859300002597, /*  359 */
128'h860ac10d842ae05ff0ef852245e000ef, /*  360 */
128'h51050513000025174e85859300002597, /*  361 */
128'h251780826151641260b2852243e000ef, /*  362 */
128'h00ef9a07af230000379752a505130000, /*  363 */
128'hf85afc56e0d2e4ceeca67159b7cd4200, /*  364 */
128'he46ee8caf0a2f486e86aec66f062f45e, /*  365 */
128'h2b17532a0a1300002a1744818aae89aa, /*  366 */
128'h0c1300002c1706000b93502b0b130000, /*  367 */
128'h841bfff58d1b4fec8c9300002c9750ec, /*  368 */
128'h69a6694664e6740670a6035441630004, /*  369 */
128'h6da26d426ce27c027ba27b427ae26a06, /*  370 */
128'h00ef855ae39d00f47793c01d80826165, /*  371 */
128'h251702879d630009079bff0489133a00, /*  372 */
128'h382000ef8552388000ef392505130000, /*  373 */
128'h4a850513000025170007c583009987b3, /*  374 */
128'h79134d81fffd4913068d126336e000ef, /*  375 */
128'hfe05879b0007c583012987b3a80500f9, /*  376 */
128'h0905344000ef856600fbe7630ff7f793, /*  377 */
128'h332000ef8552bfdd33a000ef8562b75d, /*  378 */
128'h322000ef00f4f913855aff2dcce32d85, /*  379 */
128'h0000251700f45a630009079b4124093b, /*  380 */
128'h012987b3bf15048530a000ef31450513, /*  381 */
128'h00fbe7630ff7f793fe05879b0007c583, /*  382 */
128'h2e2000ef8562b7f109052ec000ef8566, /*  383 */
128'h07b30003b6830083b7830103b703bfdd, /*  384 */
128'h0017079300d7fe6393811782278540f7, /*  385 */
128'h802345050103b78300a7002300f3b823, /*  386 */
128'h0103b7830083b7038082450180820007, /*  387 */
128'hfff706930003b7038f99920102059613, /*  388 */
128'h869b47819d9dfff7059b00c6f5638e9d, /*  389 */
128'h852e0007002300b6e6630103b7030007, /*  390 */
128'hc68300f506b300d3b823001706938082, /*  391 */
128'h000556634301bfd900d7002307850006, /*  392 */
128'h0693c21906100693430540a0053be681, /*  393 */
128'h0005089b385986ba4e250ff6f8130410, /*  394 */
128'h0306061b04ae6a630ff5761302b8f53b, /*  395 */
128'hffe302b8d53bfec68fa306850ff67613, /*  396 */
128'h00a606bb0300059340e0063b8536fcb8, /*  397 */
128'h00f5002302d007930003076302f6e963, /*  398 */
128'h081b46810015559b9d19000500230505, /*  399 */
128'h00c8063b808200b7ea630006879bfff5, /*  400 */
128'h178240f807bbb7d1feb50fa30505bf45, /*  401 */
128'h000648830007c30300d7063397ba9381, /*  402 */
128'hf0ca7119b7e101178023006600230685, /*  403 */
128'hfc86e4d6e8d2eccef4a6f8a2597d011c, /*  404 */
128'h0993f82af02ef42afc3e843684b2e0da, /*  405 */
128'h77420209591303000a9306c00a130250, /*  406 */
128'h76820017079bc52d8f1d0004c50377a2, /*  407 */
128'h039304850135086304d7ff6393811782, /*  408 */
128'h05450f630014c503bfe1e71ff0ef0201, /*  409 */
128'h879bcb9d0004c7830355106347810489, /*  410 */
128'hc503478100f6f36346a50ff7f793fd07, /*  411 */
128'h02a6eb6306d50f630640069304890014, /*  412 */
128'h08f509630630079304d50f6305800693, /*  413 */
128'h6aa66a4669e6790674a6744670e6f55d, /*  414 */
128'h048d0024c503808261090007051b6b06, /*  415 */
128'h071300a76c6306e50e6307300713b74d, /*  416 */
128'h46014685003800840b13f6e51ee30700, /*  417 */
128'h10e30780071302e5006307500713a00d, /*  418 */
128'h36134685003800840b13fa850613f6e5, /*  419 */
128'h003800840b13f8b50693a81145c10016, /*  420 */
128'h059be31ff0ef400845a946010016b693, /*  421 */
128'h4503a809dd1ff0ef0028020103930005, /*  422 */
128'h845ad89ff0ef00840b13020103930004, /*  423 */
128'h00ef852201247433600000840b13b5fd, /*  424 */
128'h715db7f18522020103930005059b6920, /*  425 */
128'he436e4c6e0c2fc3ef83aec061034f436, /*  426 */
128'hf436f032715d8082616160e2e8dff0ef, /*  427 */
128'he0c2fc3ef83aec06100005931014862e, /*  428 */
128'h710d8082616160e2e69ff0efe436e4c6, /*  429 */
128'h0808100005931234862afe36fa32f62e, /*  430 */
128'hf0efe436eec6eac2e6bee2baea22ee06, /*  431 */
128'h645260f28522f66fe0ef0808842ae3ff, /*  432 */
128'h0585230305452e0305052e8380826135, /*  433 */
128'h02938f2ae44ae826ec22110105c52883, /*  434 */
128'h8f9300001f97887687f2869a86460405, /*  435 */
128'h000fa38300b647338dfd00c6c5b3dd6f, /*  436 */
128'h9db9007585bb0fc1008fa403000f2583, /*  437 */
128'h0078159b0105883b004f2703ff4fa383, /*  438 */
128'h00f805bb0077073b0105e8330198581b, /*  439 */
128'h9e39008f23838e358e6d00f6c6339f31, /*  440 */
128'h873b008383bb8e590146561b00c6171b, /*  441 */
128'h00cf24038ef900b7c6b300d383bb00c5, /*  442 */
128'he6b30116969b00f6d39b007686bb8ebd, /*  443 */
128'h0007061b00d703bbffcfa4039fa100d3, /*  444 */
128'h00a7579b9f3d8f2d9fa1007777338f2d, /*  445 */
128'h0003869b0005881b0f418f5d0167171b, /*  446 */
128'he18f0f1300001f17f45f17e300e387bb, /*  447 */
128'he182829300001297d50f8f9300001f97, /*  448 */
128'h4383000fa58300b6c7338df100d7c5b3, /*  449 */
128'h93aa038a000f47039db9002f4403001f, /*  450 */
128'h004fa7039db9942a040a4318972a070a, /*  451 */
128'ha70301b8581b9e390058159b0105883b, /*  452 */
128'h00b7c6339f3100f805bb0105e8330003, /*  453 */
128'h561b0096139b008fa7039e398e3d8e75, /*  454 */
128'h9f3500c583bb00c3e63340189eb90176, /*  455 */
128'h0fc18eadffff44838efd0075c6b30f11, /*  456 */
128'h9fb900e6941b94aa048affcfa7039eb9, /*  457 */
128'hc7339fb900d3843b8ec140980126d69b, /*  458 */
128'h171b00c7579b9f3d007747338f6d0083, /*  459 */
128'h0004069b0003861b0005881b8f5d0147, /*  460 */
128'hd38f8f9300001f97f25f1ee300e407bb, /*  461 */
128'ha7030102c403cae383930000139782fe, /*  462 */
128'h400000c5c4b3942a040a00d7c5b30003, /*  463 */
128'h94aa048a0043a4039f210112c4839f25, /*  464 */
128'h0048171b0122c4830107083b40809e21, /*  465 */
128'h073b0083a4039e210107683301c8581b, /*  466 */
128'h159b40809e2d9ea194aa8db9048a00f8, /*  467 */
128'h05bb03c18e4d0156561b0132c90300b6, /*  468 */
128'h090a8ead00e7c6b3ffc3a4839c3500c7, /*  469 */
128'h24830106d69b9fa50106941b992a9ea1, /*  470 */
128'h9fa58f2d0007081b00d5843b8ec10009, /*  471 */
128'h02918f5d0177171b0097579b9f3d8f21, /*  472 */
128'hf45f17e300e407bb0004069b0005861b, /*  473 */
128'h45b38f5dfff64713c302829300001297, /*  474 */
128'h9f2d022fc403021fc3830002a70300d7, /*  475 */
128'h040a418c95aa058a93aa038a020fc583, /*  476 */
128'h0068171b0107083b0042a5839f2d942a, /*  477 */
128'h073b0107683301a8581b0003a5839e2d, /*  478 */
128'ha5839e2d8e3d8e59fff6c6139db100f8, /*  479 */
128'he633400c9ead0166561b00a6139b0082, /*  480 */
128'hfff7c593023fc4839ead00c703bb00c3, /*  481 */
128'h048a9db5ffc2a4038db902c10075e5b3, /*  482 */
128'h40809fa18dd50115d59b94aa00f5969b, /*  483 */
128'h9fa18f4dfff747130007081b00b385bb, /*  484 */
128'h8f5d0157171b00b7579b9f3d00774733, /*  485 */
128'h1de300e587bb0005869b0003861b0f91, /*  486 */
128'h00d306bb00fe07bb010e883b6462f3ff, /*  487 */
128'h64c2cd70cd34c97c0505282300c8863b, /*  488 */
128'hf84afc26e0a2715d653c808261056922, /*  489 */
128'h03f7f413ec56f052e486e45ee85af44e, /*  490 */
128'h0b9304000b13e53c893289ae84aa97b2, /*  491 */
128'h74639381178200078a1b408b07bb0400, /*  492 */
128'h85ce020ada93020a1a9300090a1b00f9, /*  493 */
128'h09333f4000ef0144043b865600848533, /*  494 */
128'h97824401852660bc0174176399d64159, /*  495 */
128'h6ae27a0279a2794274e2640660a6b7c9, /*  496 */
128'hf793f0227179653c808261616ba26b42, /*  497 */
128'h00178513e84af406e44eec26842a03f7, /*  498 */
128'h449d0400099300e7802397a2f8000713, /*  499 */
128'h95224581920116020006091b40a9863b, /*  500 */
128'h603cfc1c078e643c0124f563340000ef, /*  501 */
128'h64e2740270a2fd24fde3450197828522, /*  502 */
128'hd8078793000027978082614569a26942, /*  503 */
128'hd787879300002797e93c04053423639c, /*  504 */
128'h8082e13cb807879300000797ed3c639c, /*  505 */
128'h332000efec06850a4641050505931101, /*  506 */
128'h859300002597e6668693000026974701, /*  507 */
128'h070506890007c78300e107b34541c665, /*  508 */
128'hc78397ae000646038bbd962e0047d613, /*  509 */
128'h60e2fca71de3fef68fa3fec68f230007, /*  510 */
128'he122717580826105e285051300002517, /*  511 */
128'h85a26622f71ff0efe42ee5060808842a, /*  512 */
128'hf0ef0808f01ff0ef0808e85ff0ef0808, /*  513 */
128'hc703058587aa80826149640a60aaf83f, /*  514 */
128'h8c6347818082fb75fee78fa30785fff5, /*  515 */
128'h078500f506b30007470300f5873300c7, /*  516 */
128'h86930007c70387aa8082f76d00e68023, /*  517 */
128'hfee78fa30785fff5c7030585eb090017, /*  518 */
128'h87b68082e21987aab7d587b68082fb75, /*  519 */
128'hc7030585963efb7d001786930007c703, /*  520 */
128'h8023fec799e3d375fee78fa30785fff5, /*  521 */
128'h07bbfff5c78300054703058580820007, /*  522 */
128'hf37d0505e3994187d79b0187979b40f7, /*  523 */
128'h07b3a015478100e6146347018082853e, /*  524 */
128'h87bb0007c78300e587b30007c68300e5, /*  525 */
128'hfee10705e3994187d79b0187979b40f6, /*  526 */
128'h00b79363000547830ff5f5938082853e, /*  527 */
128'h0ff5f59380824501bfcd0505c3998082, /*  528 */
128'hbfcd0505dffd808200b7936300054783, /*  529 */
128'h0785808240a78533e7010007c70387aa, /*  530 */
128'hfe5ff0efec06842ae42ee8221101bfcd, /*  531 */
128'h00b78663000547830ff5f593952265a2, /*  532 */
128'h80826105644260e24501fe857be3157d, /*  533 */
128'h8533e7010007c70300b7856387aa95aa, /*  534 */
128'h468300f507334781b7fd0785808240a7, /*  535 */
128'h46030705fed60ee38082853eea990007, /*  536 */
128'h07334781bfd5872eb7d50785fa7d0007, /*  537 */
128'h00d60863a021872eca890007468300f5, /*  538 */
128'hb7c507858082853efa7d000746030705, /*  539 */
128'h0785fee68fe380824501eb1900054703, /*  540 */
128'h1101bfd587aeb7e50505fafd0007c683, /*  541 */
128'h00002797e519842a84aeec06e426e822, /*  542 */
128'hfa1ff0ef85a68522cc116380e8c78793, /*  543 */
128'he607b82300002797ef8100044783942a, /*  544 */
128'h85a68082610564a2644260e285224401, /*  545 */
128'h0023c78100054783c519f9fff0ef8522, /*  546 */
128'h1101bfd9e4a7b2230000279705050005, /*  547 */
128'hf0ef8526842ac891e822ec066104e426, /*  548 */
128'h644260e2e008050500050023c501f73f, /*  549 */
128'hcf9900054783c11d8082610564a28526, /*  550 */
128'h8082e3110017c703ce810007c68387aa, /*  551 */
128'h80824501b7e5078900d780a300e78023, /*  552 */
128'h07220ff5f69347a1eb0587aa00757713, /*  553 */
128'h8833469d00c508b387aaffed8f5537fd, /*  554 */
128'h02e787335761003657930106ee6340f8, /*  555 */
128'h07a1808200c79763963e963a97aa078e, /*  556 */
128'h0463b7f5feb78fa30785bfe9fee7bc23, /*  557 */
128'h471d4781eb9d872a8b9d00b567b304b5, /*  558 */
128'h07a100f506b30006b80300f586b3a811, /*  559 */
128'h00365793fed765e340f606b30106b023, /*  560 */
128'h00f50733963a95be078e02e787335761, /*  561 */
128'h0006c80300f586b3808200f613634781, /*  562 */
128'hf0227179b7e501068023078500f706b3, /*  563 */
128'hf0efe02ee84af406e432ec26852e842a, /*  564 */
128'h00c564636582892ace1184aa6622dd3f, /*  565 */
128'h0023f75ff0ef944a864a8522fff60913, /*  566 */
128'h8082614564e269428526740270a20004, /*  567 */
128'hf53ff0ef00a5e963842ae406e0221141, /*  568 */
128'h461386ae883280820141640260a28522, /*  569 */
128'h85b300f80733fef605e317fd4781fff6, /*  570 */
128'h4701b7e500b7002397220005c58300e6, /*  571 */
128'h00e586b300e507b3a821478100e61463, /*  572 */
128'h853ed3f59f9507050006c6830007c783, /*  573 */
128'h8de300054783808200c51363962a8082, /*  574 */
128'hec26852e842af0227179bfc50505feb7, /*  575 */
128'h0005049bd19ff0ef892ee44ef406e84a, /*  576 */
128'h408987bb008509bbd0dff0ef8522c899, /*  577 */
128'h694264e2740270a2852244010097db63, /*  578 */
128'hf83ff0ef852285ca86268082614569a2, /*  579 */
128'h00c514630ff5f593962abfe10405d17d, /*  580 */
128'hfeb70be3001507930005470380824501, /*  581 */
128'h260100c7ef630ff5f59347c1b7ed853e, /*  582 */
128'h1ce30007c7038082853e4781e60187aa, /*  583 */
128'h4721c39d00757793b7f5367d0785feb7, /*  584 */
128'hfcb69de30007c68387aa00a7083b9f1d, /*  585 */
128'h953a93011702fed819e30007869b0785, /*  586 */
128'h8fd90107179300b7e733008597938e19, /*  587 */
128'heb1187aa27018edd0036571302079693, /*  588 */
128'h367d0785f8b71fe30007c703d24d8a1d, /*  589 */
128'hc70300d80a63008785130007b803bfcd, /*  590 */
128'h87aabfa5fef51be30785f8b712e30007, /*  591 */
128'h154211418d5d05220085579bb7f1377d, /*  592 */
128'h00054703462946a54781808201419141, /*  593 */
128'h00b6e763fd07059b27018082853ee319, /*  594 */
128'h1141b7c50505fd07879b9fb902f607bb, /*  595 */
128'h00b7f86347a500a04563842ee406e022, /*  596 */
128'h753b4529fe7ff0ef357d02b455bb45a9, /*  597 */
128'hcbbfd06f03050513014160a2640202a4, /*  598 */
128'h00002717b2f73e230000271707fe4785, /*  599 */
128'h041300002417e82211018082b2f73e23, /*  600 */
128'hf0efec06600885aa84ae862ee426b2e4, /*  601 */
128'h610564a26442e00c95a660e2600cd41f, /*  602 */
128'h6380e022afc787930000279711418082, /*  603 */
128'h051300001517638caf87879300002797, /*  604 */
128'h83220000100fd08ff0ef9d81e40666e5, /*  605 */
128'h8432e406e02211418302014160a26402, /*  606 */
128'h640260a28522547d00850363ce6fe0ef, /*  607 */
128'h01258493ee2671698082450180820141, /*  608 */
128'hf0ef892eea4af222f606852689aae64e, /*  609 */
128'h0505af7ff0ef852200a484330505b03f, /*  610 */
128'hec631ff00793fff5071bee5ff0ef9522, /*  611 */
128'h458110000613a6a7a323000027970ae7, /*  612 */
128'h850a66a5859300001597c3fff0ef850a, /*  613 */
128'h00f7096302f00793012947039cbff0ef, /*  614 */
128'h85a69dfff0ef850a5e05859300001597, /*  615 */
128'h4390a2278793000027979d7ff0ef850a, /*  616 */
128'h4405c44ff0ef5c65051300001517858a, /*  617 */
128'h2717a0f7352300002717451101f41793, /*  618 */
128'h932300001797e4fff0efa0f735230000, /*  619 */
128'h76a79d2300001797e41ff0ef450178a7, /*  620 */
128'hf0dff0ef76c5859300001597854e4611, /*  621 */
128'h695264f274129c8795230000279770b2, /*  622 */
128'h272300002717200007938082615569b2, /*  623 */
128'h478de04ae426ec06e8221101b7a19af7, /*  624 */
128'hde9ff0ef84ae450d892a08c7df638432, /*  625 */
128'h55030000251708a7956325010004d783, /*  626 */
128'h06a79a6325010024d783dd3ff0ef9825, /*  627 */
128'hf0ef4511e3fff0ef00448513ffc4059b, /*  628 */
128'h5503000025176ea7972300001797db7f, /*  629 */
128'h6ca79d23000017974611da3ff0ef9525, /*  630 */
128'h4535e6fff0ef854a6d05859300001597, /*  631 */
128'hf0ef45159285d58300002597aa7fd0ef, /*  632 */
128'h879300002797a91fd0ef02000513db1f, /*  633 */
128'h90f712230000271727850007d7839127, /*  634 */
128'h0087cf63278d439c8f87879300002797, /*  635 */
128'h60e26442b16ff0ef4b85051300001517, /*  636 */
128'h64a2644260e2dddff06f6105690264a2, /*  637 */
128'h0105c703f022f4067179808261056902, /*  638 */
128'h570300e10f230115c70300e10fa34689, /*  639 */
128'h70a2740202f70a63478d00d70e6301e1, /*  640 */
128'h842aac4ff06f61454985051300001517, /*  641 */
128'h8522ab4ff0efe42e4705051300001517, /*  642 */
128'h41907402dd1ff06f614570a265a27402, /*  643 */
128'h3823dc010113ebfff06f614505c170a2, /*  644 */
128'h893284ae842a23213023229134232281, /*  645 */
128'ha25ff0ef22113c230028218006134581, /*  646 */
128'h002ca65ff0efc44a08282040061385a6, /*  647 */
128'h34832301340323813083f65ff0ef8522, /*  648 */
128'h00002797808224010113220139032281, /*  649 */
128'h59858593000015974611cb818107d783, /*  650 */
128'h1517981fd0efe40611418082d39ff06f, /*  651 */
128'ha001a9cfe0ef9a7fd0efd92505130000, /*  652 */
128'h00000000000000000000000000000000, /*  653 */
128'h00000000000000000000000000000000, /*  654 */
128'h00000000000000000000000000000000, /*  655 */
128'h46454443424139383736353433323130, /*  656 */
128'hc1bdceee242070dbe8c7b756d76aa478, /*  657 */
128'hfd469501a83046134787c62af57c0faf, /*  658 */
128'h895cd7beffff5bb18b44f7af698098d8, /*  659 */
128'h49b40821a679438efd9871936b901122, /*  660 */
128'he9b6c7aa265e5a51c040b340f61e2562, /*  661 */
128'he7d3fbc8d8a1e68102441453d62f105d, /*  662 */
128'h455a14edf4d50d87c33707d621e1cde6, /*  663 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /*  664 */
128'hfde5380c6d9d61228771f681fffa3942, /*  665 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /*  666 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /*  667 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /*  668 */
128'hfc93a039ab9423a7432aff97f4292244, /*  669 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /*  670 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /*  671 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /*  672 */
128'h0c07020d08030e09040f0a05000b0601, /*  673 */
128'h020f0c090603000d0a0704010e0b0805, /*  674 */
128'h09020b040d060f08010a030c050e0700, /*  675 */
128'h3809000038000000100c0000edfe0dd0, /*  676 */
128'h00000000100000001100000028000000, /*  677 */
128'h000000000000000000090000d8020000, /*  678 */
128'h00000000010000000000000000000000, /*  679 */
128'h02000000000000000400000003000000, /*  680 */
128'h020000000f0000000400000003000000, /*  681 */
128'h2c6874651b0000001400000003000000, /*  682 */
128'h007665642d657261622d656e61697261, /*  683 */
128'h2c687465260000001000000003000000, /*  684 */
128'h0100000000657261622d656e61697261, /*  685 */
128'h1a0000000300000000006e65736f6863, /*  686 */
128'h303140747261752f636f732f2c000000, /*  687 */
128'h0000003030323531313a303030303030, /*  688 */
128'h00000000737570630100000002000000, /*  689 */
128'h01000000000000000400000003000000, /*  690 */
128'h000000000f0000000400000003000000, /*  691 */
128'h40787d01380000000400000003000000, /*  692 */
128'h03000000000000304075706301000000, /*  693 */
128'h0300000080f0fa024b00000004000000, /*  694 */
128'h03000000007570635b00000004000000, /*  695 */
128'h03000000000000006700000004000000, /*  696 */
128'h0000000079616b6f6b00000005000000, /*  697 */
128'h2c6874651b0000001200000003000000, /*  698 */
128'h000000766373697200656e6169726120, /*  699 */
128'h34367672720000000b00000003000000, /*  700 */
128'h0b000000030000000000757363616d69, /*  701 */
128'h0000393376732c76637369727c000000, /*  702 */
128'h01000000850000000000000003000000, /*  703 */
128'h6f72746e6f632d747075727265746e69, /*  704 */
128'h04000000030000000000000072656c6c, /*  705 */
128'h0000000003000000010000008f000000, /*  706 */
128'h1b0000000f00000003000000a0000000, /*  707 */
128'h000063746e692d7570632c7663736972, /*  708 */
128'h02000000b50000000400000003000000, /*  709 */
128'h02000000bb0000000400000003000000, /*  710 */
128'h01000000020000000200000002000000, /*  711 */
128'h0030303030303030384079726f6d656d, /*  712 */
128'h6f6d656d5b0000000700000003000000, /*  713 */
128'h67000000100000000300000000007972, /*  714 */
128'h00000040000000000000008000000000, /*  715 */
128'h000000007364656c0100000002000000, /*  716 */
128'h6f6970671b0000000a00000003000000, /*  717 */
128'h72616568010000000000007364656c2d, /*  718 */
128'h0300000000000064656c2d7461656274, /*  719 */
128'h0100000001000000c30000000c000000, /*  720 */
128'hc90000000a0000000300000000000000, /*  721 */
128'h03000000000000746165627472616568, /*  722 */
128'h0200000002000000df00000000000000, /*  723 */
128'h040000000300000000636f7301000000, /*  724 */
128'h04000000030000000200000000000000, /*  725 */
128'h1f00000003000000020000000f000000, /*  726 */
128'h622d656e616972612c6874651b000000, /*  727 */
128'h622d656c706d697300636f732d657261, /*  728 */
128'hf6000000000000000300000000007375, /*  729 */
128'h30303030303240746e696c6301000000, /*  730 */
128'h1b0000000d0000000300000000000030, /*  731 */
128'h0000000030746e696c632c7663736972, /*  732 */
128'h02000000fd0000001000000003000000, /*  733 */
128'h03000000070000000200000003000000, /*  734 */
128'h00000002000000006700000010000000, /*  735 */
128'h080000000300000000000c0000000000, /*  736 */
128'h02000000006c6f72746e6f6311010000, /*  737 */
128'h6f632d747075727265746e6901000000, /*  738 */
128'h303030303030634072656c6c6f72746e, /*  739 */
128'h00000000040000000300000000000000, /*  740 */
128'h8f000000040000000300000000000000, /*  741 */
128'h1b0000000c0000000300000001000000, /*  742 */
128'h03000000003063696c702c7663736972, /*  743 */
128'h1000000003000000a000000000000000, /*  744 */
128'h020000000b00000002000000fd000000, /*  745 */
128'h67000000100000000300000009000000, /*  746 */
128'h00000004000000000000000c00000000, /*  747 */
128'h070000001b0100000400000003000000, /*  748 */
128'h030000002e0100000400000003000000, /*  749 */
128'h03000000b50000000400000003000000, /*  750 */
128'h03000000bb0000000400000003000000, /*  751 */
128'h6f632d67756265640100000002000000, /*  752 */
128'h030000000000304072656c6c6f72746e, /*  753 */
128'h65642c76637369721b00000010000000, /*  754 */
128'h0800000003000000003331302d677562, /*  755 */
128'h03000000ffff000002000000fd000000, /*  756 */
128'h00000000000000006700000010000000, /*  757 */
128'h08000000030000000010000000000000, /*  758 */
128'h02000000006c6f72746e6f6311010000, /*  759 */
128'h30303030303031407472617501000000, /*  760 */
128'h1b000000080000000300000000000030, /*  761 */
128'h1000000003000000003035373631736e, /*  762 */
128'h00000000000000100000000067000000, /*  763 */
128'h4b000000040000000300000000100000, /*  764 */
128'h39010000040000000300000080f0fa02, /*  765 */
128'h47010000040000000300000000c20100, /*  766 */
128'h58010000040000000300000003000000, /*  767 */
128'h63010000040000000300000001000000, /*  768 */
128'h6d010000040000000300000002000000, /*  769 */
128'h2d737078010000000200000004000000, /*  770 */
128'h00000000303030303030303240697073, /*  771 */
128'h786e6c781b0000002800000003000000, /*  772 */
128'h00622e30302e322d6970732d7370782c, /*  773 */
128'h302e322d6970732d7370782c786e6c78, /*  774 */
128'h00000000040000000300000000612e30, /*  775 */
128'h0f000000040000000300000001000000, /*  776 */
128'h47010000040000000300000000000000, /*  777 */
128'h58010000080000000300000003000000, /*  778 */
128'h10000000030000000200000002000000, /*  779 */
128'h00000000000000200000000067000000, /*  780 */
128'h7a010000080000000300000000100000, /*  781 */
128'h040000000300000000377865746e696b, /*  782 */
128'h04000000030000000100000086010000, /*  783 */
128'h04000000030000000100000096010000, /*  784 */
128'h040000000300000008000000a7010000, /*  785 */
128'h40636d6d0100000004000000be010000, /*  786 */
128'h1b0000000d0000000300000000000030, /*  787 */
128'h00000000746f6c732d6970732d636d6d, /*  788 */
128'h00000000670000000400000003000000, /*  789 */
128'h20bcbe00cd0100000400000003000000, /*  790 */
128'he40c0000df0100000800000003000000, /*  791 */
128'hee0100000000000003000000e40c0000, /*  792 */
128'h72776f6c010000000200000002000000, /*  793 */
128'h3030303030303033406874652d637369, /*  794 */
128'h1b0000000c0000000300000000000000, /*  795 */
128'h03000000006874652d63736972776f6c, /*  796 */
128'h006b726f7774656e5b00000008000000, /*  797 */
128'h03000000470100000400000003000000, /*  798 */
128'h03000000580100000800000003000000, /*  799 */
128'hf9010000060000000300000000000000, /*  800 */
128'h100000000300000000007fe3023e1800, /*  801 */
128'h00000000000000300000000067000000, /*  802 */
128'h6f697067010000000200000000800000, /*  803 */
128'h03000000000000303030303030303440, /*  804 */
128'h03000000020000000b02000004000000, /*  805 */
128'h7370782c786e6c781b00000015000000, /*  806 */
128'h00000000612e30302e312d6f6970672d, /*  807 */
128'h03000000170200000000000003000000, /*  808 */
128'h00000040000000006700000010000000, /*  809 */
128'h04000000030000000000010000000000, /*  810 */
128'h04000000030000000000000027020000, /*  811 */
128'h04000000030000000000000037020000, /*  812 */
128'h04000000030000000000000049020000, /*  813 */
128'h0400000003000000000000005b020000, /*  814 */
128'h0400000003000000080000006f020000, /*  815 */
128'h0400000003000000080000007f020000, /*  816 */
128'h04000000030000000000000090020000, /*  817 */
128'h040000000300000001000000a7020000, /*  818 */
128'h0400000003000000ffffffffb4020000, /*  819 */
128'h0400000003000000ffffffffc5020000, /*  820 */
128'h040000000300000001000000b5000000, /*  821 */
128'h020000000200000001000000bb000000, /*  822 */
128'h73736572646461230900000002000000, /*  823 */
128'h6c65632d657a69732300736c6c65632d, /*  824 */
128'h6f6d00656c62697461706d6f6300736c, /*  825 */
128'h00687461702d74756f647473006c6564, /*  826 */
128'h6e6575716572662d65736162656d6974, /*  827 */
128'h6e6575716572662d6b636f6c63007963, /*  828 */
128'h7200657079745f656369766564007963, /*  829 */
128'h2c766373697200737574617473006765, /*  830 */
128'h626c7400657079742d756d6d00617369, /*  831 */
128'h7075727265746e69230074696c70732d, /*  832 */
128'h7075727265746e6900736c6c65632d74, /*  833 */
128'h6e696c0072656c6c6f72746e6f632d74, /*  834 */
128'h736f69706700656c646e6168702c7875, /*  835 */
128'h742d746c75616665642c78756e696c00, /*  836 */
128'h74732d6e696174657200726567676972, /*  837 */
128'h6172006465646e65707375732d657461, /*  838 */
128'h2d73747075727265746e69007365676e, /*  839 */
128'h6d616e2d676572006465646e65747865, /*  840 */
128'h6972702d78616d2c7663736972007365, /*  841 */
128'h7665646e2c766373697200797469726f, /*  842 */
128'h690064656570732d746e657272756300, /*  843 */
128'h00746e657261702d747075727265746e, /*  844 */
128'h732d6765720073747075727265746e69, /*  845 */
128'h746469772d6f692d6765720074666968, /*  846 */
128'h6c7800796c696d61662c786e6c780068, /*  847 */
128'h6c780074736978652d6f6669662c786e, /*  848 */
128'h7800737469622d73732d6d756e2c786e, /*  849 */
128'h726566736e6172742d6d756e2c786e6c, /*  850 */
128'h722d6b63732c786e6c7800737469622d, /*  851 */
128'h6572662d78616d2d697073006f697461, /*  852 */
128'h722d656761746c6f760079636e657571, /*  853 */
128'h70772d656c6261736964007365676e61, /*  854 */
128'h65726464612d63616d2d6c61636f6c00, /*  855 */
128'h6700736c6c65632d6f69706723007373, /*  856 */
128'h780072656c6c6f72746e6f632d6f6970, /*  857 */
128'h7800737475706e692d6c6c612c786e6c, /*  858 */
128'h322d737475706e692d6c6c612c786e6c, /*  859 */
128'h75616665642d74756f642c786e6c7800, /*  860 */
128'h6665642d74756f642c786e6c7800746c, /*  861 */
128'h6f6970672c786e6c7800322d746c7561, /*  862 */
128'h6f6970672c786e6c780068746469772d, /*  863 */
128'h746e692c786e6c780068746469772d32, /*  864 */
128'h7800746e65736572702d747075727265, /*  865 */
128'h786e6c78006c6175642d73692c786e6c, /*  866 */
128'h6e6c7800746c75616665642d6972742c, /*  867 */
128'h00322d746c75616665642d6972742c78, /*  868 */
128'h00000a0d21646c726f57206f6c6c6548, /*  869 */
128'h464f5f4f4c43414d00000a0d70617274, /*  870 */
128'h464f5f494843414d0000000054455346, /*  871 */
128'h46464f5f524c50540000000054455346, /*  872 */
128'h46464f5f534346540000000000544553, /*  873 */
128'h4c5254434f49444d0000000000544553, /*  874 */
128'h46464f5f534346520054455346464f5f, /*  875 */
128'h5346464f5f5253520000000000544553, /*  876 */
128'h46464f5f444142520000000000005445, /*  877 */
128'h46464f5f524c50520000000000544553, /*  878 */
128'h000000003f3f3f3f0000000000544553, /*  879 */
128'h000064252b54455346464f5f524c5052, /*  880 */
128'h6f746f72502050490000000000000047, /*  881 */
128'h00000000000000000a50495049203d20, /*  882 */
128'h6f746f72502050490000000000000054, /*  883 */
128'h6f746f7250205049000a504745203d20, /*  884 */
128'h6165682074736574000a505550203d20, /*  885 */
128'h6e6f6320747365740000000a3a726564, /*  886 */
128'h6f746f7250205049000a3a73746e6574, /*  887 */
128'h6f746f7250205049000a504449203d20, /*  888 */
128'h6f746f725020504900000a5054203d20, /*  889 */
128'h00000000000000000a50434344203d20, /*  890 */
128'h6f746f72502050490000000000000036, /*  891 */
128'h00000000000000000a50565352203d20, /*  892 */
128'h000a455247203d206f746f7250205049, /*  893 */
128'h000a505345203d206f746f7250205049, /*  894 */
128'h00000a4841203d206f746f7250205049, /*  895 */
128'h000a50544d203d206f746f7250205049, /*  896 */
128'h5054454542203d206f746f7250205049, /*  897 */
128'h6f746f72502050490000000000000a48, /*  898 */
128'h000000000000000a5041434e45203d20, /*  899 */
128'h6f746f7250205049000000000000004d, /*  900 */
128'h00000000000000000a504d4f43203d20, /*  901 */
128'h0a50544353203d206f746f7250205049, /*  902 */
128'h6f746f72502050490000000000000000, /*  903 */
128'h00000000000a4554494c504455203d20, /*  904 */
128'h0a534c504d203d206f746f7250205049, /*  905 */
128'h6f746f72502050490000000000000000, /*  906 */
128'h6f746f7270205049000a574152203d20, /*  907 */
128'h2820646574726f707075736e75203d20, /*  908 */
128'h79745f6f746f7270000000000a297825, /*  909 */
128'h0000000000000a78257830203d206570, /*  910 */
128'h727265746e692064656c646e61686e75, /*  911 */
128'h414d2070757465530000000a21747075, /*  912 */
128'h6c25203d2043414d000a726464612043, /*  913 */
128'h726464612043414d00000a786c253a78, /*  914 */
128'h3a783230253a78323025203d20737365, /*  915 */
128'h253a783230253a783230253a78323025, /*  916 */
128'h74656e72656874450000000a2e783230, /*  917 */
128'h757461747320747075727265746e6920, /*  918 */
128'h00000000000000000a646c25203d2073, /*  919 */
128'h20646564616f6c2065687420746f6f42, /*  920 */
128'h00000000000a2e2e2e6d6172676f7270, /*  921 */
128'h207265746f6f62202c657962646f6f47, /*  922 */
128'h746e692070636864000000000a2e2e2e, /*  923 */
128'h0a7025202c726f727265206c616e7265, /*  924 */
128'h20676e69646e65530000000000000000, /*  925 */
128'h0000000a545345555145525f50434844, /*  926 */
128'h000000000000000a4b43412050434844, /*  927 */
128'h4120504920746e65696c432050434844, /*  928 */
128'h252e64252e642520203a737365726464, /*  929 */
128'h49207265767265530000000a64252e64, /*  930 */
128'h252e642520203a737365726464412050, /*  931 */
128'h00000000000000000a64252e64252e64, /*  932 */
128'h203a7373657264646120726574756f52, /*  933 */
128'h0000000a64252e64252e64252e642520, /*  934 */
128'h73736572646461206b73616d2074654e, /*  935 */
128'h000a64252e64252e64252e642520203a, /*  936 */
128'h0a6425203d20656d697420657361654c, /*  937 */
128'h3d206e69616d6f640000000000000000, /*  938 */
128'h3d2072657672657300000a2273252220, /*  939 */
128'h50494b53204b434100000a2273252220, /*  940 */
128'h4b414e2050434844000000000a444550, /*  941 */
128'h6574736575716552000000000000000a, /*  942 */
128'h65737566657220737365726464612064, /*  943 */
128'h732520726f7272450000000000000a64, /*  944 */
128'h656c646e61686e75000000000000000a, /*  945 */
128'h000000000a6425206e6f6974706f2064, /*  946 */
128'h6f20504348442064656c646e61686e55, /*  947 */
128'h000000000000000a64252065646f6370, /*  948 */
128'h5349445f5043484420676e69646e6553, /*  949 */
128'h2528726f72726570000a595245564f43, /*  950 */
128'h000000003068746500000000000a2973, /*  951 */
128'h30253a58323025203a2043414d207325, /*  952 */
128'h3230253a583230253a583230253a5832, /*  953 */
128'h74276e646c756f43000a583230253a58, /*  954 */
128'h4f43534944205043484420646e657320, /*  955 */
128'h2520656369766564206e6f2059524556, /*  956 */
128'h20676e697469615700000a7325203a73, /*  957 */
128'h000a524546464f5f5043484420726f66, /*  958 */
128'h00000000000000202020202020202020, /*  959 */
128'h000000000000002e0000000000006325, /*  960 */
128'h00000000002020200000005832302520, /*  961 */
128'h66656463626139383736353433323130, /*  962 */
128'h6e656c20656c69460000000000000000, /*  963 */
128'h000000000000000a6425203d20687467, /*  964 */
128'h732522203a717277000000000000002f, /*  965 */
128'h0a64253d657a69736b636f6c62202c22, /*  966 */
128'h20657669656365520000000000000000, /*  967 */
128'h0000000000000a2e646e6520656c6966, /*  968 */
128'h656c6c6163207172775f656c646e6168, /*  969 */
128'h206c6167656c6c4900000000000a2e64, /*  970 */
128'h0a2e6e6f6974617265706f2050544654, /*  971 */
128'h00000000300000000000000000000000, /*  972 */
128'h00000000ffffffff0000000000000000, /*  973 */
128'h000000030f060301000000000c000000, /*  974 */
128'hefcdab89674523010000000087ff3cc0, /*  975 */
128'h000000000000000000000000000000fe, /*  976 */
128'h00000000000000000000000000000000, /*  977 */
128'h00000000000000000000000000000000, /*  978 */
128'h00000000000000000000000000000000, /*  979 */
128'h00000000000000000000000000000000, /*  980 */
128'h00000000000000000000000000000000, /*  981 */
128'h00000000000000000000000000000000, /*  982 */
128'h00000000000000000000000000000000, /*  983 */
128'h00000000000000000000000000000000, /*  984 */
128'h00000000000000000000000000000000, /*  985 */
128'h00000000000000000000000000000000, /*  986 */
128'h00000000000000000000000000000000, /*  987 */
128'h00000000000000000000000000000000, /*  988 */
128'h00000000000000000000000000000000, /*  989 */
128'h00000000000000000000000000000000, /*  990 */
128'h00000000000000000000000000000000, /*  991 */
128'h00000000000000000000000000000000, /*  992 */
128'h00000000000000000000000000000000, /*  993 */
128'h00000000000000000000000000000000, /*  994 */
128'h00000000000000000000000000000000, /*  995 */
128'h00000000000000000000000000000000, /*  996 */
128'h00000000000000000000000000000000, /*  997 */
128'h00000000000000000000000000000000, /*  998 */
128'h00000000000000000000000000000000, /*  999 */
128'h00000000000000000000000000000000, /* 1000 */
128'h00000000000000000000000000000000, /* 1001 */
128'h00000000000000000000000000000000, /* 1002 */
128'h00000000000000000000000000000000, /* 1003 */
128'h00000000000000000000000000000000, /* 1004 */
128'h00000000000000000000000000000000, /* 1005 */
128'h00000000000000000000000000000000, /* 1006 */
128'h00000000000000000000000000000000, /* 1007 */
128'h00000000000000000000000000000000, /* 1008 */
128'h00000000000000000000000000000000, /* 1009 */
128'h00000000000000000000000000000000, /* 1010 */
128'h00000000000000000000000000000000, /* 1011 */
128'h00000000000000000000000000000000, /* 1012 */
128'h00000000000000000000000000000000, /* 1013 */
128'h00000000000000000000000000000000, /* 1014 */
128'h00000000000000000000000000000000, /* 1015 */
128'h00000000000000000000000000000000, /* 1016 */
128'h00000000000000000000000000000000, /* 1017 */
128'h00000000000000000000000000000000, /* 1018 */
128'h00000000000000000000000000000000, /* 1019 */
128'h00000000000000000000000000000000, /* 1020 */
128'h00000000000000000000000000000000, /* 1021 */
128'h00000000000000000000000000000000, /* 1022 */
128'h00000000000000000000000000000000, /* 1023 */
128'h00000000000000000000000000000000, /* 1024 */
128'h00000000000000000000000000000000, /* 1025 */
128'h00000000000000000000000000000000, /* 1026 */
128'h00000000000000000000000000000000, /* 1027 */
128'h00000000000000000000000000000000, /* 1028 */
128'h00000000000000000000000000000000, /* 1029 */
128'h00000000000000000000000000000000, /* 1030 */
128'h00000000000000000000000000000000, /* 1031 */
128'h00000000000000000000000000000000, /* 1032 */
128'h00000000000000000000000000000000, /* 1033 */
128'h00000000000000000000000000000000, /* 1034 */
128'h00000000000000000000000000000000, /* 1035 */
128'h00000000000000000000000000000000, /* 1036 */
128'h00000000000000000000000000000000, /* 1037 */
128'h00000000000000000000000000000000, /* 1038 */
128'h00000000000000000000000000000000, /* 1039 */
128'h00000000000000000000000000000000, /* 1040 */
128'h00000000000000000000000000000000, /* 1041 */
128'h00000000000000000000000000000000, /* 1042 */
128'h00000000000000000000000000000000, /* 1043 */
128'h00000000000000000000000000000000, /* 1044 */
128'h00000000000000000000000000000000, /* 1045 */
128'h00000000000000000000000000000000, /* 1046 */
128'h00000000000000000000000000000000, /* 1047 */
128'h00000000000000000000000000000000, /* 1048 */
128'h00000000000000000000000000000000, /* 1049 */
128'h00000000000000000000000000000000, /* 1050 */
128'h00000000000000000000000000000000, /* 1051 */
128'h00000000000000000000000000000000, /* 1052 */
128'h00000000000000000000000000000000, /* 1053 */
128'h00000000000000000000000000000000, /* 1054 */
128'h00000000000000000000000000000000, /* 1055 */
128'h00000000000000000000000000000000, /* 1056 */
128'h00000000000000000000000000000000, /* 1057 */
128'h00000000000000000000000000000000, /* 1058 */
128'h00000000000000000000000000000000, /* 1059 */
128'h00000000000000000000000000000000, /* 1060 */
128'h00000000000000000000000000000000, /* 1061 */
128'h00000000000000000000000000000000, /* 1062 */
128'h00000000000000000000000000000000, /* 1063 */
128'h00000000000000000000000000000000, /* 1064 */
128'h00000000000000000000000000000000, /* 1065 */
128'h00000000000000000000000000000000, /* 1066 */
128'h00000000000000000000000000000000, /* 1067 */
128'h00000000000000000000000000000000, /* 1068 */
128'h00000000000000000000000000000000, /* 1069 */
128'h00000000000000000000000000000000, /* 1070 */
128'h00000000000000000000000000000000, /* 1071 */
128'h00000000000000000000000000000000, /* 1072 */
128'h00000000000000000000000000000000, /* 1073 */
128'h00000000000000000000000000000000, /* 1074 */
128'h00000000000000000000000000000000, /* 1075 */
128'h00000000000000000000000000000000, /* 1076 */
128'h00000000000000000000000000000000, /* 1077 */
128'h00000000000000000000000000000000, /* 1078 */
128'h00000000000000000000000000000000, /* 1079 */
128'h00000000000000000000000000000000, /* 1080 */
128'h00000000000000000000000000000000, /* 1081 */
128'h00000000000000000000000000000000, /* 1082 */
128'h00000000000000000000000000000000, /* 1083 */
128'h00000000000000000000000000000000, /* 1084 */
128'h00000000000000000000000000000000, /* 1085 */
128'h00000000000000000000000000000000, /* 1086 */
128'h00000000000000000000000000000000, /* 1087 */
128'h00000000000000000000000000000000, /* 1088 */
128'h00000000000000000000000000000000, /* 1089 */
128'h00000000000000000000000000000000, /* 1090 */
128'h00000000000000000000000000000000, /* 1091 */
128'h00000000000000000000000000000000, /* 1092 */
128'h00000000000000000000000000000000, /* 1093 */
128'h00000000000000000000000000000000, /* 1094 */
128'h00000000000000000000000000000000, /* 1095 */
128'h00000000000000000000000000000000, /* 1096 */
128'h00000000000000000000000000000000, /* 1097 */
128'h00000000000000000000000000000000, /* 1098 */
128'h00000000000000000000000000000000, /* 1099 */
128'h00000000000000000000000000000000, /* 1100 */
128'h00000000000000000000000000000000, /* 1101 */
128'h00000000000000000000000000000000, /* 1102 */
128'h00000000000000000000000000000000, /* 1103 */
128'h00000000000000000000000000000000, /* 1104 */
128'h00000000000000000000000000000000, /* 1105 */
128'h00000000000000000000000000000000, /* 1106 */
128'h00000000000000000000000000000000, /* 1107 */
128'h00000000000000000000000000000000, /* 1108 */
128'h00000000000000000000000000000000, /* 1109 */
128'h00000000000000000000000000000000, /* 1110 */
128'h00000000000000000000000000000000, /* 1111 */
128'h00000000000000000000000000000000, /* 1112 */
128'h00000000000000000000000000000000, /* 1113 */
128'h00000000000000000000000000000000, /* 1114 */
128'h00000000000000000000000000000000, /* 1115 */
128'h00000000000000000000000000000000, /* 1116 */
128'h00000000000000000000000000000000, /* 1117 */
128'h00000000000000000000000000000000, /* 1118 */
128'h00000000000000000000000000000000, /* 1119 */
128'h00000000000000000000000000000000, /* 1120 */
128'h00000000000000000000000000000000, /* 1121 */
128'h00000000000000000000000000000000, /* 1122 */
128'h00000000000000000000000000000000, /* 1123 */
128'h00000000000000000000000000000000, /* 1124 */
128'h00000000000000000000000000000000, /* 1125 */
128'h00000000000000000000000000000000, /* 1126 */
128'h00000000000000000000000000000000, /* 1127 */
128'h00000000000000000000000000000000, /* 1128 */
128'h00000000000000000000000000000000, /* 1129 */
128'h00000000000000000000000000000000, /* 1130 */
128'h00000000000000000000000000000000, /* 1131 */
128'h00000000000000000000000000000000, /* 1132 */
128'h00000000000000000000000000000000, /* 1133 */
128'h00000000000000000000000000000000, /* 1134 */
128'h00000000000000000000000000000000, /* 1135 */
128'h00000000000000000000000000000000, /* 1136 */
128'h00000000000000000000000000000000, /* 1137 */
128'h00000000000000000000000000000000, /* 1138 */
128'h00000000000000000000000000000000, /* 1139 */
128'h00000000000000000000000000000000, /* 1140 */
128'h00000000000000000000000000000000, /* 1141 */
128'h00000000000000000000000000000000, /* 1142 */
128'h00000000000000000000000000000000, /* 1143 */
128'h00000000000000000000000000000000, /* 1144 */
128'h00000000000000000000000000000000, /* 1145 */
128'h00000000000000000000000000000000, /* 1146 */
128'h00000000000000000000000000000000, /* 1147 */
128'h00000000000000000000000000000000, /* 1148 */
128'h00000000000000000000000000000000, /* 1149 */
128'h00000000000000000000000000000000, /* 1150 */
128'h00000000000000000000000000000000, /* 1151 */
128'h00000000000000000000000000000000, /* 1152 */
128'h00000000000000000000000000000000, /* 1153 */
128'h00000000000000000000000000000000, /* 1154 */
128'h00000000000000000000000000000000, /* 1155 */
128'h00000000000000000000000000000000, /* 1156 */
128'h00000000000000000000000000000000, /* 1157 */
128'h00000000000000000000000000000000, /* 1158 */
128'h00000000000000000000000000000000, /* 1159 */
128'h00000000000000000000000000000000, /* 1160 */
128'h00000000000000000000000000000000, /* 1161 */
128'h00000000000000000000000000000000, /* 1162 */
128'h00000000000000000000000000000000, /* 1163 */
128'h00000000000000000000000000000000, /* 1164 */
128'h00000000000000000000000000000000, /* 1165 */
128'h00000000000000000000000000000000, /* 1166 */
128'h00000000000000000000000000000000, /* 1167 */
128'h00000000000000000000000000000000, /* 1168 */
128'h00000000000000000000000000000000, /* 1169 */
128'h00000000000000000000000000000000, /* 1170 */
128'h00000000000000000000000000000000, /* 1171 */
128'h00000000000000000000000000000000, /* 1172 */
128'h00000000000000000000000000000000, /* 1173 */
128'h00000000000000000000000000000000, /* 1174 */
128'h00000000000000000000000000000000, /* 1175 */
128'h00000000000000000000000000000000, /* 1176 */
128'h00000000000000000000000000000000, /* 1177 */
128'h00000000000000000000000000000000, /* 1178 */
128'h00000000000000000000000000000000, /* 1179 */
128'h00000000000000000000000000000000, /* 1180 */
128'h00000000000000000000000000000000, /* 1181 */
128'h00000000000000000000000000000000, /* 1182 */
128'h00000000000000000000000000000000, /* 1183 */
128'h00000000000000000000000000000000, /* 1184 */
128'h00000000000000000000000000000000, /* 1185 */
128'h00000000000000000000000000000000, /* 1186 */
128'h00000000000000000000000000000000, /* 1187 */
128'h00000000000000000000000000000000, /* 1188 */
128'h00000000000000000000000000000000, /* 1189 */
128'h00000000000000000000000000000000, /* 1190 */
128'h00000000000000000000000000000000, /* 1191 */
128'h00000000000000000000000000000000, /* 1192 */
128'h00000000000000000000000000000000, /* 1193 */
128'h00000000000000000000000000000000, /* 1194 */
128'h00000000000000000000000000000000, /* 1195 */
128'h00000000000000000000000000000000, /* 1196 */
128'h00000000000000000000000000000000, /* 1197 */
128'h00000000000000000000000000000000, /* 1198 */
128'h00000000000000000000000000000000, /* 1199 */
128'h00000000000000000000000000000000, /* 1200 */
128'h00000000000000000000000000000000, /* 1201 */
128'h00000000000000000000000000000000, /* 1202 */
128'h00000000000000000000000000000000, /* 1203 */
128'h00000000000000000000000000000000, /* 1204 */
128'h00000000000000000000000000000000, /* 1205 */
128'h00000000000000000000000000000000, /* 1206 */
128'h00000000000000000000000000000000, /* 1207 */
128'h00000000000000000000000000000000, /* 1208 */
128'h00000000000000000000000000000000, /* 1209 */
128'h00000000000000000000000000000000, /* 1210 */
128'h00000000000000000000000000000000, /* 1211 */
128'h00000000000000000000000000000000, /* 1212 */
128'h00000000000000000000000000000000, /* 1213 */
128'h00000000000000000000000000000000, /* 1214 */
128'h00000000000000000000000000000000, /* 1215 */
128'h00000000000000000000000000000000, /* 1216 */
128'h00000000000000000000000000000000, /* 1217 */
128'h00000000000000000000000000000000, /* 1218 */
128'h00000000000000000000000000000000, /* 1219 */
128'h00000000000000000000000000000000, /* 1220 */
128'h00000000000000000000000000000000, /* 1221 */
128'h00000000000000000000000000000000, /* 1222 */
128'h00000000000000000000000000000000, /* 1223 */
128'h00000000000000000000000000000000, /* 1224 */
128'h00000000000000000000000000000000, /* 1225 */
128'h00000000000000000000000000000000, /* 1226 */
128'h00000000000000000000000000000000, /* 1227 */
128'h00000000000000000000000000000000, /* 1228 */
128'h00000000000000000000000000000000, /* 1229 */
128'h00000000000000000000000000000000, /* 1230 */
128'h00000000000000000000000000000000, /* 1231 */
128'h00000000000000000000000000000000, /* 1232 */
128'h00000000000000000000000000000000, /* 1233 */
128'h00000000000000000000000000000000, /* 1234 */
128'h00000000000000000000000000000000, /* 1235 */
128'h00000000000000000000000000000000, /* 1236 */
128'h00000000000000000000000000000000, /* 1237 */
128'h00000000000000000000000000000000, /* 1238 */
128'h00000000000000000000000000000000, /* 1239 */
128'h00000000000000000000000000000000, /* 1240 */
128'h00000000000000000000000000000000, /* 1241 */
128'h00000000000000000000000000000000, /* 1242 */
128'h00000000000000000000000000000000, /* 1243 */
128'h00000000000000000000000000000000, /* 1244 */
128'h00000000000000000000000000000000, /* 1245 */
128'h00000000000000000000000000000000, /* 1246 */
128'h00000000000000000000000000000000, /* 1247 */
128'h00000000000000000000000000000000, /* 1248 */
128'h00000000000000000000000000000000, /* 1249 */
128'h00000000000000000000000000000000, /* 1250 */
128'h00000000000000000000000000000000, /* 1251 */
128'h00000000000000000000000000000000, /* 1252 */
128'h00000000000000000000000000000000, /* 1253 */
128'h00000000000000000000000000000000, /* 1254 */
128'h00000000000000000000000000000000, /* 1255 */
128'h00000000000000000000000000000000, /* 1256 */
128'h00000000000000000000000000000000, /* 1257 */
128'h00000000000000000000000000000000, /* 1258 */
128'h00000000000000000000000000000000, /* 1259 */
128'h00000000000000000000000000000000, /* 1260 */
128'h00000000000000000000000000000000, /* 1261 */
128'h00000000000000000000000000000000, /* 1262 */
128'h00000000000000000000000000000000, /* 1263 */
128'h00000000000000000000000000000000, /* 1264 */
128'h00000000000000000000000000000000, /* 1265 */
128'h00000000000000000000000000000000, /* 1266 */
128'h00000000000000000000000000000000, /* 1267 */
128'h00000000000000000000000000000000, /* 1268 */
128'h00000000000000000000000000000000, /* 1269 */
128'h00000000000000000000000000000000, /* 1270 */
128'h00000000000000000000000000000000, /* 1271 */
128'h00000000000000000000000000000000, /* 1272 */
128'h00000000000000000000000000000000, /* 1273 */
128'h00000000000000000000000000000000, /* 1274 */
128'h00000000000000000000000000000000, /* 1275 */
128'h00000000000000000000000000000000, /* 1276 */
128'h00000000000000000000000000000000, /* 1277 */
128'h00000000000000000000000000000000, /* 1278 */
128'h00000000000000000000000000000000, /* 1279 */
128'h00000000000000000000000000000000, /* 1280 */
128'h00000000000000000000000000000000, /* 1281 */
128'h00000000000000000000000000000000, /* 1282 */
128'h00000000000000000000000000000000, /* 1283 */
128'h00000000000000000000000000000000, /* 1284 */
128'h00000000000000000000000000000000, /* 1285 */
128'h00000000000000000000000000000000, /* 1286 */
128'h00000000000000000000000000000000, /* 1287 */
128'h00000000000000000000000000000000, /* 1288 */
128'h00000000000000000000000000000000, /* 1289 */
128'h00000000000000000000000000000000, /* 1290 */
128'h00000000000000000000000000000000, /* 1291 */
128'h00000000000000000000000000000000, /* 1292 */
128'h00000000000000000000000000000000, /* 1293 */
128'h00000000000000000000000000000000, /* 1294 */
128'h00000000000000000000000000000000, /* 1295 */
128'h00000000000000000000000000000000, /* 1296 */
128'h00000000000000000000000000000000, /* 1297 */
128'h00000000000000000000000000000000, /* 1298 */
128'h00000000000000000000000000000000, /* 1299 */
128'h00000000000000000000000000000000, /* 1300 */
128'h00000000000000000000000000000000, /* 1301 */
128'h00000000000000000000000000000000, /* 1302 */
128'h00000000000000000000000000000000, /* 1303 */
128'h00000000000000000000000000000000, /* 1304 */
128'h00000000000000000000000000000000, /* 1305 */
128'h00000000000000000000000000000000, /* 1306 */
128'h00000000000000000000000000000000, /* 1307 */
128'h00000000000000000000000000000000, /* 1308 */
128'h00000000000000000000000000000000, /* 1309 */
128'h00000000000000000000000000000000, /* 1310 */
128'h00000000000000000000000000000000, /* 1311 */
128'h00000000000000000000000000000000, /* 1312 */
128'h00000000000000000000000000000000, /* 1313 */
128'h00000000000000000000000000000000, /* 1314 */
128'h00000000000000000000000000000000, /* 1315 */
128'h00000000000000000000000000000000, /* 1316 */
128'h00000000000000000000000000000000, /* 1317 */
128'h00000000000000000000000000000000, /* 1318 */
128'h00000000000000000000000000000000, /* 1319 */
128'h00000000000000000000000000000000, /* 1320 */
128'h00000000000000000000000000000000, /* 1321 */
128'h00000000000000000000000000000000, /* 1322 */
128'h00000000000000000000000000000000, /* 1323 */
128'h00000000000000000000000000000000, /* 1324 */
128'h00000000000000000000000000000000, /* 1325 */
128'h00000000000000000000000000000000, /* 1326 */
128'h00000000000000000000000000000000, /* 1327 */
128'h00000000000000000000000000000000, /* 1328 */
128'h00000000000000000000000000000000, /* 1329 */
128'h00000000000000000000000000000000, /* 1330 */
128'h00000000000000000000000000000000, /* 1331 */
128'h00000000000000000000000000000000, /* 1332 */
128'h00000000000000000000000000000000, /* 1333 */
128'h00000000000000000000000000000000, /* 1334 */
128'h00000000000000000000000000000000, /* 1335 */
128'h00000000000000000000000000000000, /* 1336 */
128'h00000000000000000000000000000000, /* 1337 */
128'h00000000000000000000000000000000, /* 1338 */
128'h00000000000000000000000000000000, /* 1339 */
128'h00000000000000000000000000000000, /* 1340 */
128'h00000000000000000000000000000000, /* 1341 */
128'h00000000000000000000000000000000, /* 1342 */
128'h00000000000000000000000000000000, /* 1343 */
128'h00000000000000000000000000000000, /* 1344 */
128'h00000000000000000000000000000000, /* 1345 */
128'h00000000000000000000000000000000, /* 1346 */
128'h00000000000000000000000000000000, /* 1347 */
128'h00000000000000000000000000000000, /* 1348 */
128'h00000000000000000000000000000000, /* 1349 */
128'h00000000000000000000000000000000, /* 1350 */
128'h00000000000000000000000000000000, /* 1351 */
128'h00000000000000000000000000000000, /* 1352 */
128'h00000000000000000000000000000000, /* 1353 */
128'h00000000000000000000000000000000, /* 1354 */
128'h00000000000000000000000000000000, /* 1355 */
128'h00000000000000000000000000000000, /* 1356 */
128'h00000000000000000000000000000000, /* 1357 */
128'h00000000000000000000000000000000, /* 1358 */
128'h00000000000000000000000000000000, /* 1359 */
128'h00000000000000000000000000000000, /* 1360 */
128'h00000000000000000000000000000000, /* 1361 */
128'h00000000000000000000000000000000, /* 1362 */
128'h00000000000000000000000000000000, /* 1363 */
128'h00000000000000000000000000000000, /* 1364 */
128'h00000000000000000000000000000000, /* 1365 */
128'h00000000000000000000000000000000, /* 1366 */
128'h00000000000000000000000000000000, /* 1367 */
128'h00000000000000000000000000000000, /* 1368 */
128'h00000000000000000000000000000000, /* 1369 */
128'h00000000000000000000000000000000, /* 1370 */
128'h00000000000000000000000000000000, /* 1371 */
128'h00000000000000000000000000000000, /* 1372 */
128'h00000000000000000000000000000000, /* 1373 */
128'h00000000000000000000000000000000, /* 1374 */
128'h00000000000000000000000000000000, /* 1375 */
128'h00000000000000000000000000000000, /* 1376 */
128'h00000000000000000000000000000000, /* 1377 */
128'h00000000000000000000000000000000, /* 1378 */
128'h00000000000000000000000000000000, /* 1379 */
128'h00000000000000000000000000000000, /* 1380 */
128'h00000000000000000000000000000000, /* 1381 */
128'h00000000000000000000000000000000, /* 1382 */
128'h00000000000000000000000000000000, /* 1383 */
128'h00000000000000000000000000000000, /* 1384 */
128'h00000000000000000000000000000000, /* 1385 */
128'h00000000000000000000000000000000, /* 1386 */
128'h00000000000000000000000000000000, /* 1387 */
128'h00000000000000000000000000000000, /* 1388 */
128'h00000000000000000000000000000000, /* 1389 */
128'h00000000000000000000000000000000, /* 1390 */
128'h00000000000000000000000000000000, /* 1391 */
128'h00000000000000000000000000000000, /* 1392 */
128'h00000000000000000000000000000000, /* 1393 */
128'h00000000000000000000000000000000, /* 1394 */
128'h00000000000000000000000000000000, /* 1395 */
128'h00000000000000000000000000000000, /* 1396 */
128'h00000000000000000000000000000000, /* 1397 */
128'h00000000000000000000000000000000, /* 1398 */
128'h00000000000000000000000000000000, /* 1399 */
128'h00000000000000000000000000000000, /* 1400 */
128'h00000000000000000000000000000000, /* 1401 */
128'h00000000000000000000000000000000, /* 1402 */
128'h00000000000000000000000000000000, /* 1403 */
128'h00000000000000000000000000000000, /* 1404 */
128'h00000000000000000000000000000000, /* 1405 */
128'h00000000000000000000000000000000, /* 1406 */
128'h00000000000000000000000000000000, /* 1407 */
128'h00000000000000000000000000000000, /* 1408 */
128'h00000000000000000000000000000000, /* 1409 */
128'h00000000000000000000000000000000, /* 1410 */
128'h00000000000000000000000000000000, /* 1411 */
128'h00000000000000000000000000000000, /* 1412 */
128'h00000000000000000000000000000000, /* 1413 */
128'h00000000000000000000000000000000, /* 1414 */
128'h00000000000000000000000000000000, /* 1415 */
128'h00000000000000000000000000000000, /* 1416 */
128'h00000000000000000000000000000000, /* 1417 */
128'h00000000000000000000000000000000, /* 1418 */
128'h00000000000000000000000000000000, /* 1419 */
128'h00000000000000000000000000000000, /* 1420 */
128'h00000000000000000000000000000000, /* 1421 */
128'h00000000000000000000000000000000, /* 1422 */
128'h00000000000000000000000000000000, /* 1423 */
128'h00000000000000000000000000000000, /* 1424 */
128'h00000000000000000000000000000000, /* 1425 */
128'h00000000000000000000000000000000, /* 1426 */
128'h00000000000000000000000000000000, /* 1427 */
128'h00000000000000000000000000000000, /* 1428 */
128'h00000000000000000000000000000000, /* 1429 */
128'h00000000000000000000000000000000, /* 1430 */
128'h00000000000000000000000000000000, /* 1431 */
128'h00000000000000000000000000000000, /* 1432 */
128'h00000000000000000000000000000000, /* 1433 */
128'h00000000000000000000000000000000, /* 1434 */
128'h00000000000000000000000000000000, /* 1435 */
128'h00000000000000000000000000000000, /* 1436 */
128'h00000000000000000000000000000000, /* 1437 */
128'h00000000000000000000000000000000, /* 1438 */
128'h00000000000000000000000000000000, /* 1439 */
128'h00000000000000000000000000000000, /* 1440 */
128'h00000000000000000000000000000000, /* 1441 */
128'h00000000000000000000000000000000, /* 1442 */
128'h00000000000000000000000000000000, /* 1443 */
128'h00000000000000000000000000000000, /* 1444 */
128'h00000000000000000000000000000000, /* 1445 */
128'h00000000000000000000000000000000, /* 1446 */
128'h00000000000000000000000000000000, /* 1447 */
128'h00000000000000000000000000000000, /* 1448 */
128'h00000000000000000000000000000000, /* 1449 */
128'h00000000000000000000000000000000, /* 1450 */
128'h00000000000000000000000000000000, /* 1451 */
128'h00000000000000000000000000000000, /* 1452 */
128'h00000000000000000000000000000000, /* 1453 */
128'h00000000000000000000000000000000, /* 1454 */
128'h00000000000000000000000000000000, /* 1455 */
128'h00000000000000000000000000000000, /* 1456 */
128'h00000000000000000000000000000000, /* 1457 */
128'h00000000000000000000000000000000, /* 1458 */
128'h00000000000000000000000000000000, /* 1459 */
128'h00000000000000000000000000000000, /* 1460 */
128'h00000000000000000000000000000000, /* 1461 */
128'h00000000000000000000000000000000, /* 1462 */
128'h00000000000000000000000000000000, /* 1463 */
128'h00000000000000000000000000000000, /* 1464 */
128'h00000000000000000000000000000000, /* 1465 */
128'h00000000000000000000000000000000, /* 1466 */
128'h00000000000000000000000000000000, /* 1467 */
128'h00000000000000000000000000000000, /* 1468 */
128'h00000000000000000000000000000000, /* 1469 */
128'h00000000000000000000000000000000, /* 1470 */
128'h00000000000000000000000000000000, /* 1471 */
128'h00000000000000000000000000000000, /* 1472 */
128'h00000000000000000000000000000000, /* 1473 */
128'h00000000000000000000000000000000, /* 1474 */
128'h00000000000000000000000000000000, /* 1475 */
128'h00000000000000000000000000000000, /* 1476 */
128'h00000000000000000000000000000000, /* 1477 */
128'h00000000000000000000000000000000, /* 1478 */
128'h00000000000000000000000000000000, /* 1479 */
128'h00000000000000000000000000000000, /* 1480 */
128'h00000000000000000000000000000000, /* 1481 */
128'h00000000000000000000000000000000, /* 1482 */
128'h00000000000000000000000000000000, /* 1483 */
128'h00000000000000000000000000000000, /* 1484 */
128'h00000000000000000000000000000000, /* 1485 */
128'h00000000000000000000000000000000, /* 1486 */
128'h00000000000000000000000000000000, /* 1487 */
128'h00000000000000000000000000000000, /* 1488 */
128'h00000000000000000000000000000000, /* 1489 */
128'h00000000000000000000000000000000, /* 1490 */
128'h00000000000000000000000000000000, /* 1491 */
128'h00000000000000000000000000000000, /* 1492 */
128'h00000000000000000000000000000000, /* 1493 */
128'h00000000000000000000000000000000, /* 1494 */
128'h00000000000000000000000000000000, /* 1495 */
128'h00000000000000000000000000000000, /* 1496 */
128'h00000000000000000000000000000000, /* 1497 */
128'h00000000000000000000000000000000, /* 1498 */
128'h00000000000000000000000000000000, /* 1499 */
128'h00000000000000000000000000000000, /* 1500 */
128'h00000000000000000000000000000000, /* 1501 */
128'h00000000000000000000000000000000, /* 1502 */
128'h00000000000000000000000000000000, /* 1503 */
128'h00000000000000000000000000000000, /* 1504 */
128'h00000000000000000000000000000000, /* 1505 */
128'h00000000000000000000000000000000, /* 1506 */
128'h00000000000000000000000000000000, /* 1507 */
128'h00000000000000000000000000000000, /* 1508 */
128'h00000000000000000000000000000000, /* 1509 */
128'h00000000000000000000000000000000, /* 1510 */
128'h00000000000000000000000000000000, /* 1511 */
128'h00000000000000000000000000000000, /* 1512 */
128'h00000000000000000000000000000000, /* 1513 */
128'h00000000000000000000000000000000, /* 1514 */
128'h00000000000000000000000000000000, /* 1515 */
128'h00000000000000000000000000000000, /* 1516 */
128'h00000000000000000000000000000000, /* 1517 */
128'h00000000000000000000000000000000, /* 1518 */
128'h00000000000000000000000000000000, /* 1519 */
128'h00000000000000000000000000000000, /* 1520 */
128'h00000000000000000000000000000000, /* 1521 */
128'h00000000000000000000000000000000, /* 1522 */
128'h00000000000000000000000000000000, /* 1523 */
128'h00000000000000000000000000000000, /* 1524 */
128'h00000000000000000000000000000000, /* 1525 */
128'h00000000000000000000000000000000, /* 1526 */
128'h00000000000000000000000000000000, /* 1527 */
128'h00000000000000000000000000000000, /* 1528 */
128'h00000000000000000000000000000000, /* 1529 */
128'h00000000000000000000000000000000, /* 1530 */
128'h00000000000000000000000000000000, /* 1531 */
128'h00000000000000000000000000000000, /* 1532 */
128'h00000000000000000000000000000000, /* 1533 */
128'h00000000000000000000000000000000, /* 1534 */
128'h00000000000000000000000000000000, /* 1535 */
128'h00000000000000000000000000000000, /* 1536 */
128'h00000000000000000000000000000000, /* 1537 */
128'h00000000000000000000000000000000, /* 1538 */
128'h00000000000000000000000000000000, /* 1539 */
128'h00000000000000000000000000000000, /* 1540 */
128'h00000000000000000000000000000000, /* 1541 */
128'h00000000000000000000000000000000, /* 1542 */
128'h00000000000000000000000000000000, /* 1543 */
128'h00000000000000000000000000000000, /* 1544 */
128'h00000000000000000000000000000000, /* 1545 */
128'h00000000000000000000000000000000, /* 1546 */
128'h00000000000000000000000000000000, /* 1547 */
128'h00000000000000000000000000000000, /* 1548 */
128'h00000000000000000000000000000000, /* 1549 */
128'h00000000000000000000000000000000, /* 1550 */
128'h00000000000000000000000000000000, /* 1551 */
128'h00000000000000000000000000000000, /* 1552 */
128'h00000000000000000000000000000000, /* 1553 */
128'h00000000000000000000000000000000, /* 1554 */
128'h00000000000000000000000000000000, /* 1555 */
128'h00000000000000000000000000000000, /* 1556 */
128'h00000000000000000000000000000000, /* 1557 */
128'h00000000000000000000000000000000, /* 1558 */
128'h00000000000000000000000000000000, /* 1559 */
128'h00000000000000000000000000000000, /* 1560 */
128'h00000000000000000000000000000000, /* 1561 */
128'h00000000000000000000000000000000, /* 1562 */
128'h00000000000000000000000000000000, /* 1563 */
128'h00000000000000000000000000000000, /* 1564 */
128'h00000000000000000000000000000000, /* 1565 */
128'h00000000000000000000000000000000, /* 1566 */
128'h00000000000000000000000000000000, /* 1567 */
128'h00000000000000000000000000000000, /* 1568 */
128'h00000000000000000000000000000000, /* 1569 */
128'h00000000000000000000000000000000, /* 1570 */
128'h00000000000000000000000000000000, /* 1571 */
128'h00000000000000000000000000000000, /* 1572 */
128'h00000000000000000000000000000000, /* 1573 */
128'h00000000000000000000000000000000, /* 1574 */
128'h00000000000000000000000000000000, /* 1575 */
128'h00000000000000000000000000000000, /* 1576 */
128'h00000000000000000000000000000000, /* 1577 */
128'h00000000000000000000000000000000, /* 1578 */
128'h00000000000000000000000000000000, /* 1579 */
128'h00000000000000000000000000000000, /* 1580 */
128'h00000000000000000000000000000000, /* 1581 */
128'h00000000000000000000000000000000, /* 1582 */
128'h00000000000000000000000000000000, /* 1583 */
128'h00000000000000000000000000000000, /* 1584 */
128'h00000000000000000000000000000000, /* 1585 */
128'h00000000000000000000000000000000, /* 1586 */
128'h00000000000000000000000000000000, /* 1587 */
128'h00000000000000000000000000000000, /* 1588 */
128'h00000000000000000000000000000000, /* 1589 */
128'h00000000000000000000000000000000, /* 1590 */
128'h00000000000000000000000000000000, /* 1591 */
128'h00000000000000000000000000000000, /* 1592 */
128'h00000000000000000000000000000000, /* 1593 */
128'h00000000000000000000000000000000, /* 1594 */
128'h00000000000000000000000000000000, /* 1595 */
128'h00000000000000000000000000000000, /* 1596 */
128'h00000000000000000000000000000000, /* 1597 */
128'h00000000000000000000000000000000, /* 1598 */
128'h00000000000000000000000000000000, /* 1599 */
128'h00000000000000000000000000000000, /* 1600 */
128'h00000000000000000000000000000000, /* 1601 */
128'h00000000000000000000000000000000, /* 1602 */
128'h00000000000000000000000000000000, /* 1603 */
128'h00000000000000000000000000000000, /* 1604 */
128'h00000000000000000000000000000000, /* 1605 */
128'h00000000000000000000000000000000, /* 1606 */
128'h00000000000000000000000000000000, /* 1607 */
128'h00000000000000000000000000000000, /* 1608 */
128'h00000000000000000000000000000000, /* 1609 */
128'h00000000000000000000000000000000, /* 1610 */
128'h00000000000000000000000000000000, /* 1611 */
128'h00000000000000000000000000000000, /* 1612 */
128'h00000000000000000000000000000000, /* 1613 */
128'h00000000000000000000000000000000, /* 1614 */
128'h00000000000000000000000000000000, /* 1615 */
128'h00000000000000000000000000000000, /* 1616 */
128'h00000000000000000000000000000000, /* 1617 */
128'h00000000000000000000000000000000, /* 1618 */
128'h00000000000000000000000000000000, /* 1619 */
128'h00000000000000000000000000000000, /* 1620 */
128'h00000000000000000000000000000000, /* 1621 */
128'h00000000000000000000000000000000, /* 1622 */
128'h00000000000000000000000000000000, /* 1623 */
128'h00000000000000000000000000000000, /* 1624 */
128'h00000000000000000000000000000000, /* 1625 */
128'h00000000000000000000000000000000, /* 1626 */
128'h00000000000000000000000000000000, /* 1627 */
128'h00000000000000000000000000000000, /* 1628 */
128'h00000000000000000000000000000000, /* 1629 */
128'h00000000000000000000000000000000, /* 1630 */
128'h00000000000000000000000000000000, /* 1631 */
128'h00000000000000000000000000000000, /* 1632 */
128'h00000000000000000000000000000000, /* 1633 */
128'h00000000000000000000000000000000, /* 1634 */
128'h00000000000000000000000000000000, /* 1635 */
128'h00000000000000000000000000000000, /* 1636 */
128'h00000000000000000000000000000000, /* 1637 */
128'h00000000000000000000000000000000, /* 1638 */
128'h00000000000000000000000000000000, /* 1639 */
128'h00000000000000000000000000000000, /* 1640 */
128'h00000000000000000000000000000000, /* 1641 */
128'h00000000000000000000000000000000, /* 1642 */
128'h00000000000000000000000000000000, /* 1643 */
128'h00000000000000000000000000000000, /* 1644 */
128'h00000000000000000000000000000000, /* 1645 */
128'h00000000000000000000000000000000, /* 1646 */
128'h00000000000000000000000000000000, /* 1647 */
128'h00000000000000000000000000000000, /* 1648 */
128'h00000000000000000000000000000000, /* 1649 */
128'h00000000000000000000000000000000, /* 1650 */
128'h00000000000000000000000000000000, /* 1651 */
128'h00000000000000000000000000000000, /* 1652 */
128'h00000000000000000000000000000000, /* 1653 */
128'h00000000000000000000000000000000, /* 1654 */
128'h00000000000000000000000000000000, /* 1655 */
128'h00000000000000000000000000000000, /* 1656 */
128'h00000000000000000000000000000000, /* 1657 */
128'h00000000000000000000000000000000, /* 1658 */
128'h00000000000000000000000000000000, /* 1659 */
128'h00000000000000000000000000000000, /* 1660 */
128'h00000000000000000000000000000000, /* 1661 */
128'h00000000000000000000000000000000, /* 1662 */
128'h00000000000000000000000000000000, /* 1663 */
128'h00000000000000000000000000000000, /* 1664 */
128'h00000000000000000000000000000000, /* 1665 */
128'h00000000000000000000000000000000, /* 1666 */
128'h00000000000000000000000000000000, /* 1667 */
128'h00000000000000000000000000000000, /* 1668 */
128'h00000000000000000000000000000000, /* 1669 */
128'h00000000000000000000000000000000, /* 1670 */
128'h00000000000000000000000000000000, /* 1671 */
128'h00000000000000000000000000000000, /* 1672 */
128'h00000000000000000000000000000000, /* 1673 */
128'h00000000000000000000000000000000, /* 1674 */
128'h00000000000000000000000000000000, /* 1675 */
128'h00000000000000000000000000000000, /* 1676 */
128'h00000000000000000000000000000000, /* 1677 */
128'h00000000000000000000000000000000, /* 1678 */
128'h00000000000000000000000000000000, /* 1679 */
128'h00000000000000000000000000000000, /* 1680 */
128'h00000000000000000000000000000000, /* 1681 */
128'h00000000000000000000000000000000, /* 1682 */
128'h00000000000000000000000000000000, /* 1683 */
128'h00000000000000000000000000000000, /* 1684 */
128'h00000000000000000000000000000000, /* 1685 */
128'h00000000000000000000000000000000, /* 1686 */
128'h00000000000000000000000000000000, /* 1687 */
128'h00000000000000000000000000000000, /* 1688 */
128'h00000000000000000000000000000000, /* 1689 */
128'h00000000000000000000000000000000, /* 1690 */
128'h00000000000000000000000000000000, /* 1691 */
128'h00000000000000000000000000000000, /* 1692 */
128'h00000000000000000000000000000000, /* 1693 */
128'h00000000000000000000000000000000, /* 1694 */
128'h00000000000000000000000000000000, /* 1695 */
128'h00000000000000000000000000000000, /* 1696 */
128'h00000000000000000000000000000000, /* 1697 */
128'h00000000000000000000000000000000, /* 1698 */
128'h00000000000000000000000000000000, /* 1699 */
128'h00000000000000000000000000000000, /* 1700 */
128'h00000000000000000000000000000000, /* 1701 */
128'h00000000000000000000000000000000, /* 1702 */
128'h00000000000000000000000000000000, /* 1703 */
128'h00000000000000000000000000000000, /* 1704 */
128'h00000000000000000000000000000000, /* 1705 */
128'h00000000000000000000000000000000, /* 1706 */
128'h00000000000000000000000000000000, /* 1707 */
128'h00000000000000000000000000000000, /* 1708 */
128'h00000000000000000000000000000000, /* 1709 */
128'h00000000000000000000000000000000, /* 1710 */
128'h00000000000000000000000000000000, /* 1711 */
128'h00000000000000000000000000000000, /* 1712 */
128'h00000000000000000000000000000000, /* 1713 */
128'h00000000000000000000000000000000, /* 1714 */
128'h00000000000000000000000000000000, /* 1715 */
128'h00000000000000000000000000000000, /* 1716 */
128'h00000000000000000000000000000000, /* 1717 */
128'h00000000000000000000000000000000, /* 1718 */
128'h00000000000000000000000000000000, /* 1719 */
128'h00000000000000000000000000000000, /* 1720 */
128'h00000000000000000000000000000000, /* 1721 */
128'h00000000000000000000000000000000, /* 1722 */
128'h00000000000000000000000000000000, /* 1723 */
128'h00000000000000000000000000000000, /* 1724 */
128'h00000000000000000000000000000000, /* 1725 */
128'h00000000000000000000000000000000, /* 1726 */
128'h00000000000000000000000000000000, /* 1727 */
128'h00000000000000000000000000000000, /* 1728 */
128'h00000000000000000000000000000000, /* 1729 */
128'h00000000000000000000000000000000, /* 1730 */
128'h00000000000000000000000000000000, /* 1731 */
128'h00000000000000000000000000000000, /* 1732 */
128'h00000000000000000000000000000000, /* 1733 */
128'h00000000000000000000000000000000, /* 1734 */
128'h00000000000000000000000000000000, /* 1735 */
128'h00000000000000000000000000000000, /* 1736 */
128'h00000000000000000000000000000000, /* 1737 */
128'h00000000000000000000000000000000, /* 1738 */
128'h00000000000000000000000000000000, /* 1739 */
128'h00000000000000000000000000000000, /* 1740 */
128'h00000000000000000000000000000000, /* 1741 */
128'h00000000000000000000000000000000, /* 1742 */
128'h00000000000000000000000000000000, /* 1743 */
128'h00000000000000000000000000000000, /* 1744 */
128'h00000000000000000000000000000000, /* 1745 */
128'h00000000000000000000000000000000, /* 1746 */
128'h00000000000000000000000000000000, /* 1747 */
128'h00000000000000000000000000000000, /* 1748 */
128'h00000000000000000000000000000000, /* 1749 */
128'h00000000000000000000000000000000, /* 1750 */
128'h00000000000000000000000000000000, /* 1751 */
128'h00000000000000000000000000000000, /* 1752 */
128'h00000000000000000000000000000000, /* 1753 */
128'h00000000000000000000000000000000, /* 1754 */
128'h00000000000000000000000000000000, /* 1755 */
128'h00000000000000000000000000000000, /* 1756 */
128'h00000000000000000000000000000000, /* 1757 */
128'h00000000000000000000000000000000, /* 1758 */
128'h00000000000000000000000000000000, /* 1759 */
128'h00000000000000000000000000000000, /* 1760 */
128'h00000000000000000000000000000000, /* 1761 */
128'h00000000000000000000000000000000, /* 1762 */
128'h00000000000000000000000000000000, /* 1763 */
128'h00000000000000000000000000000000, /* 1764 */
128'h00000000000000000000000000000000, /* 1765 */
128'h00000000000000000000000000000000, /* 1766 */
128'h00000000000000000000000000000000, /* 1767 */
128'h00000000000000000000000000000000, /* 1768 */
128'h00000000000000000000000000000000, /* 1769 */
128'h00000000000000000000000000000000, /* 1770 */
128'h00000000000000000000000000000000, /* 1771 */
128'h00000000000000000000000000000000, /* 1772 */
128'h00000000000000000000000000000000, /* 1773 */
128'h00000000000000000000000000000000, /* 1774 */
128'h00000000000000000000000000000000, /* 1775 */
128'h00000000000000000000000000000000, /* 1776 */
128'h00000000000000000000000000000000, /* 1777 */
128'h00000000000000000000000000000000, /* 1778 */
128'h00000000000000000000000000000000, /* 1779 */
128'h00000000000000000000000000000000, /* 1780 */
128'h00000000000000000000000000000000, /* 1781 */
128'h00000000000000000000000000000000, /* 1782 */
128'h00000000000000000000000000000000, /* 1783 */
128'h00000000000000000000000000000000, /* 1784 */
128'h00000000000000000000000000000000, /* 1785 */
128'h00000000000000000000000000000000, /* 1786 */
128'h00000000000000000000000000000000, /* 1787 */
128'h00000000000000000000000000000000, /* 1788 */
128'h00000000000000000000000000000000, /* 1789 */
128'h00000000000000000000000000000000, /* 1790 */
128'h00000000000000000000000000000000, /* 1791 */
128'h00000000000000000000000000000000, /* 1792 */
128'h00000000000000000000000000000000, /* 1793 */
128'h00000000000000000000000000000000, /* 1794 */
128'h00000000000000000000000000000000, /* 1795 */
128'h00000000000000000000000000000000, /* 1796 */
128'h00000000000000000000000000000000, /* 1797 */
128'h00000000000000000000000000000000, /* 1798 */
128'h00000000000000000000000000000000, /* 1799 */
128'h00000000000000000000000000000000, /* 1800 */
128'h00000000000000000000000000000000, /* 1801 */
128'h00000000000000000000000000000000, /* 1802 */
128'h00000000000000000000000000000000, /* 1803 */
128'h00000000000000000000000000000000, /* 1804 */
128'h00000000000000000000000000000000, /* 1805 */
128'h00000000000000000000000000000000, /* 1806 */
128'h00000000000000000000000000000000, /* 1807 */
128'h00000000000000000000000000000000, /* 1808 */
128'h00000000000000000000000000000000, /* 1809 */
128'h00000000000000000000000000000000, /* 1810 */
128'h00000000000000000000000000000000, /* 1811 */
128'h00000000000000000000000000000000, /* 1812 */
128'h00000000000000000000000000000000, /* 1813 */
128'h00000000000000000000000000000000, /* 1814 */
128'h00000000000000000000000000000000, /* 1815 */
128'h00000000000000000000000000000000, /* 1816 */
128'h00000000000000000000000000000000, /* 1817 */
128'h00000000000000000000000000000000, /* 1818 */
128'h00000000000000000000000000000000, /* 1819 */
128'h00000000000000000000000000000000, /* 1820 */
128'h00000000000000000000000000000000, /* 1821 */
128'h00000000000000000000000000000000, /* 1822 */
128'h00000000000000000000000000000000, /* 1823 */
128'h00000000000000000000000000000000, /* 1824 */
128'h00000000000000000000000000000000, /* 1825 */
128'h00000000000000000000000000000000, /* 1826 */
128'h00000000000000000000000000000000, /* 1827 */
128'h00000000000000000000000000000000, /* 1828 */
128'h00000000000000000000000000000000, /* 1829 */
128'h00000000000000000000000000000000, /* 1830 */
128'h00000000000000000000000000000000, /* 1831 */
128'h00000000000000000000000000000000, /* 1832 */
128'h00000000000000000000000000000000, /* 1833 */
128'h00000000000000000000000000000000, /* 1834 */
128'h00000000000000000000000000000000, /* 1835 */
128'h00000000000000000000000000000000, /* 1836 */
128'h00000000000000000000000000000000, /* 1837 */
128'h00000000000000000000000000000000, /* 1838 */
128'h00000000000000000000000000000000, /* 1839 */
128'h00000000000000000000000000000000, /* 1840 */
128'h00000000000000000000000000000000, /* 1841 */
128'h00000000000000000000000000000000, /* 1842 */
128'h00000000000000000000000000000000, /* 1843 */
128'h00000000000000000000000000000000, /* 1844 */
128'h00000000000000000000000000000000, /* 1845 */
128'h00000000000000000000000000000000, /* 1846 */
128'h00000000000000000000000000000000, /* 1847 */
128'h00000000000000000000000000000000, /* 1848 */
128'h00000000000000000000000000000000, /* 1849 */
128'h00000000000000000000000000000000, /* 1850 */
128'h00000000000000000000000000000000, /* 1851 */
128'h00000000000000000000000000000000, /* 1852 */
128'h00000000000000000000000000000000, /* 1853 */
128'h00000000000000000000000000000000, /* 1854 */
128'h00000000000000000000000000000000, /* 1855 */
128'h00000000000000000000000000000000, /* 1856 */
128'h00000000000000000000000000000000, /* 1857 */
128'h00000000000000000000000000000000, /* 1858 */
128'h00000000000000000000000000000000, /* 1859 */
128'h00000000000000000000000000000000, /* 1860 */
128'h00000000000000000000000000000000, /* 1861 */
128'h00000000000000000000000000000000, /* 1862 */
128'h00000000000000000000000000000000, /* 1863 */
128'h00000000000000000000000000000000, /* 1864 */
128'h00000000000000000000000000000000, /* 1865 */
128'h00000000000000000000000000000000, /* 1866 */
128'h00000000000000000000000000000000, /* 1867 */
128'h00000000000000000000000000000000, /* 1868 */
128'h00000000000000000000000000000000, /* 1869 */
128'h00000000000000000000000000000000, /* 1870 */
128'h00000000000000000000000000000000, /* 1871 */
128'h00000000000000000000000000000000, /* 1872 */
128'h00000000000000000000000000000000, /* 1873 */
128'h00000000000000000000000000000000, /* 1874 */
128'h00000000000000000000000000000000, /* 1875 */
128'h00000000000000000000000000000000, /* 1876 */
128'h00000000000000000000000000000000, /* 1877 */
128'h00000000000000000000000000000000, /* 1878 */
128'h00000000000000000000000000000000, /* 1879 */
128'h00000000000000000000000000000000, /* 1880 */
128'h00000000000000000000000000000000, /* 1881 */
128'h00000000000000000000000000000000, /* 1882 */
128'h00000000000000000000000000000000, /* 1883 */
128'h00000000000000000000000000000000, /* 1884 */
128'h00000000000000000000000000000000, /* 1885 */
128'h00000000000000000000000000000000, /* 1886 */
128'h00000000000000000000000000000000, /* 1887 */
128'h00000000000000000000000000000000, /* 1888 */
128'h00000000000000000000000000000000, /* 1889 */
128'h00000000000000000000000000000000, /* 1890 */
128'h00000000000000000000000000000000, /* 1891 */
128'h00000000000000000000000000000000, /* 1892 */
128'h00000000000000000000000000000000, /* 1893 */
128'h00000000000000000000000000000000, /* 1894 */
128'h00000000000000000000000000000000, /* 1895 */
128'h00000000000000000000000000000000, /* 1896 */
128'h00000000000000000000000000000000, /* 1897 */
128'h00000000000000000000000000000000, /* 1898 */
128'h00000000000000000000000000000000, /* 1899 */
128'h00000000000000000000000000000000, /* 1900 */
128'h00000000000000000000000000000000, /* 1901 */
128'h00000000000000000000000000000000, /* 1902 */
128'h00000000000000000000000000000000, /* 1903 */
128'h00000000000000000000000000000000, /* 1904 */
128'h00000000000000000000000000000000, /* 1905 */
128'h00000000000000000000000000000000, /* 1906 */
128'h00000000000000000000000000000000, /* 1907 */
128'h00000000000000000000000000000000, /* 1908 */
128'h00000000000000000000000000000000, /* 1909 */
128'h00000000000000000000000000000000, /* 1910 */
128'h00000000000000000000000000000000, /* 1911 */
128'h00000000000000000000000000000000, /* 1912 */
128'h00000000000000000000000000000000, /* 1913 */
128'h00000000000000000000000000000000, /* 1914 */
128'h00000000000000000000000000000000, /* 1915 */
128'h00000000000000000000000000000000, /* 1916 */
128'h00000000000000000000000000000000, /* 1917 */
128'h00000000000000000000000000000000, /* 1918 */
128'h00000000000000000000000000000000, /* 1919 */
128'h00000000000000000000000000000000, /* 1920 */
128'h00000000000000000000000000000000, /* 1921 */
128'h00000000000000000000000000000000, /* 1922 */
128'h00000000000000000000000000000000, /* 1923 */
128'h00000000000000000000000000000000, /* 1924 */
128'h00000000000000000000000000000000, /* 1925 */
128'h00000000000000000000000000000000, /* 1926 */
128'h00000000000000000000000000000000, /* 1927 */
128'h00000000000000000000000000000000, /* 1928 */
128'h00000000000000000000000000000000, /* 1929 */
128'h00000000000000000000000000000000, /* 1930 */
128'h00000000000000000000000000000000, /* 1931 */
128'h00000000000000000000000000000000, /* 1932 */
128'h00000000000000000000000000000000, /* 1933 */
128'h00000000000000000000000000000000, /* 1934 */
128'h00000000000000000000000000000000, /* 1935 */
128'h00000000000000000000000000000000, /* 1936 */
128'h00000000000000000000000000000000, /* 1937 */
128'h00000000000000000000000000000000, /* 1938 */
128'h00000000000000000000000000000000, /* 1939 */
128'h00000000000000000000000000000000, /* 1940 */
128'h00000000000000000000000000000000, /* 1941 */
128'h00000000000000000000000000000000, /* 1942 */
128'h00000000000000000000000000000000, /* 1943 */
128'h00000000000000000000000000000000, /* 1944 */
128'h00000000000000000000000000000000, /* 1945 */
128'h00000000000000000000000000000000, /* 1946 */
128'h00000000000000000000000000000000, /* 1947 */
128'h00000000000000000000000000000000, /* 1948 */
128'h00000000000000000000000000000000, /* 1949 */
128'h00000000000000000000000000000000, /* 1950 */
128'h00000000000000000000000000000000, /* 1951 */
128'h00000000000000000000000000000000, /* 1952 */
128'h00000000000000000000000000000000, /* 1953 */
128'h00000000000000000000000000000000, /* 1954 */
128'h00000000000000000000000000000000, /* 1955 */
128'h00000000000000000000000000000000, /* 1956 */
128'h00000000000000000000000000000000, /* 1957 */
128'h00000000000000000000000000000000, /* 1958 */
128'h00000000000000000000000000000000, /* 1959 */
128'h00000000000000000000000000000000, /* 1960 */
128'h00000000000000000000000000000000, /* 1961 */
128'h00000000000000000000000000000000, /* 1962 */
128'h00000000000000000000000000000000, /* 1963 */
128'h00000000000000000000000000000000, /* 1964 */
128'h00000000000000000000000000000000, /* 1965 */
128'h00000000000000000000000000000000, /* 1966 */
128'h00000000000000000000000000000000, /* 1967 */
128'h00000000000000000000000000000000, /* 1968 */
128'h00000000000000000000000000000000, /* 1969 */
128'h00000000000000000000000000000000, /* 1970 */
128'h00000000000000000000000000000000, /* 1971 */
128'h00000000000000000000000000000000, /* 1972 */
128'h00000000000000000000000000000000, /* 1973 */
128'h00000000000000000000000000000000, /* 1974 */
128'h00000000000000000000000000000000, /* 1975 */
128'h00000000000000000000000000000000, /* 1976 */
128'h00000000000000000000000000000000, /* 1977 */
128'h00000000000000000000000000000000, /* 1978 */
128'h00000000000000000000000000000000, /* 1979 */
128'h00000000000000000000000000000000, /* 1980 */
128'h00000000000000000000000000000000, /* 1981 */
128'h00000000000000000000000000000000, /* 1982 */
128'h00000000000000000000000000000000, /* 1983 */
128'h00000000000000000000000000000000, /* 1984 */
128'h00000000000000000000000000000000, /* 1985 */
128'h00000000000000000000000000000000, /* 1986 */
128'h00000000000000000000000000000000, /* 1987 */
128'h00000000000000000000000000000000, /* 1988 */
128'h00000000000000000000000000000000, /* 1989 */
128'h00000000000000000000000000000000, /* 1990 */
128'h00000000000000000000000000000000, /* 1991 */
128'h00000000000000000000000000000000, /* 1992 */
128'h00000000000000000000000000000000, /* 1993 */
128'h00000000000000000000000000000000, /* 1994 */
128'h00000000000000000000000000000000, /* 1995 */
128'h00000000000000000000000000000000, /* 1996 */
128'h00000000000000000000000000000000, /* 1997 */
128'h00000000000000000000000000000000, /* 1998 */
128'h00000000000000000000000000000000, /* 1999 */
128'h00000000000000000000000000000000, /* 2000 */
128'h00000000000000000000000000000000, /* 2001 */
128'h00000000000000000000000000000000, /* 2002 */
128'h00000000000000000000000000000000, /* 2003 */
128'h00000000000000000000000000000000, /* 2004 */
128'h00000000000000000000000000000000, /* 2005 */
128'h00000000000000000000000000000000, /* 2006 */
128'h00000000000000000000000000000000, /* 2007 */
128'h00000000000000000000000000000000, /* 2008 */
128'h00000000000000000000000000000000, /* 2009 */
128'h00000000000000000000000000000000, /* 2010 */
128'h00000000000000000000000000000000, /* 2011 */
128'h00000000000000000000000000000000, /* 2012 */
128'h00000000000000000000000000000000, /* 2013 */
128'h00000000000000000000000000000000, /* 2014 */
128'h00000000000000000000000000000000, /* 2015 */
128'h00000000000000000000000000000000, /* 2016 */
128'h00000000000000000000000000000000, /* 2017 */
128'h00000000000000000000000000000000, /* 2018 */
128'h00000000000000000000000000000000, /* 2019 */
128'h00000000000000000000000000000000, /* 2020 */
128'h00000000000000000000000000000000, /* 2021 */
128'h00000000000000000000000000000000, /* 2022 */
128'h00000000000000000000000000000000, /* 2023 */
128'h00000000000000000000000000000000, /* 2024 */
128'h00000000000000000000000000000000, /* 2025 */
128'h00000000000000000000000000000000, /* 2026 */
128'h00000000000000000000000000000000, /* 2027 */
128'h00000000000000000000000000000000, /* 2028 */
128'h00000000000000000000000000000000, /* 2029 */
128'h00000000000000000000000000000000, /* 2030 */
128'h00000000000000000000000000000000, /* 2031 */
128'h00000000000000000000000000000000, /* 2032 */
128'h00000000000000000000000000000000, /* 2033 */
128'h00000000000000000000000000000000, /* 2034 */
128'h00000000000000000000000000000000, /* 2035 */
128'h00000000000000000000000000000000, /* 2036 */
128'h00000000000000000000000000000000, /* 2037 */
128'h00000000000000000000000000000000, /* 2038 */
128'h00000000000000000000000000000000, /* 2039 */
128'h00000000000000000000000000000000, /* 2040 */
128'h00000000000000000000000000000000, /* 2041 */
128'h00000000000000000000000000000000, /* 2042 */
128'h00000000000000000000000000000000, /* 2043 */
128'h00000000000000000000000000000000, /* 2044 */
128'h00000000000000000000000000000000, /* 2045 */
128'h00000000000000000000000000000000, /* 2046 */
128'h00000000000000000000000000000000, /* 2047 */
128'h00000000000000000000000000000000, /* 2048 */
128'h00000000000000000000000000000000, /* 2049 */
128'h00000000000000000000000000000000, /* 2050 */
128'h00000000000000000000000000000000, /* 2051 */
128'h00000000000000000000000000000000, /* 2052 */
128'h00000000000000000000000000000000, /* 2053 */
128'h00000000000000000000000000000000, /* 2054 */
128'h00000000000000000000000000000000, /* 2055 */
128'h00000000000000000000000000000000, /* 2056 */
128'h00000000000000000000000000000000, /* 2057 */
128'h00000000000000000000000000000000, /* 2058 */
128'h00000000000000000000000000000000, /* 2059 */
128'h00000000000000000000000000000000, /* 2060 */
128'h00000000000000000000000000000000, /* 2061 */
128'h00000000000000000000000000000000, /* 2062 */
128'h00000000000000000000000000000000, /* 2063 */
128'h00000000000000000000000000000000, /* 2064 */
128'h00000000000000000000000000000000, /* 2065 */
128'h00000000000000000000000000000000, /* 2066 */
128'h00000000000000000000000000000000, /* 2067 */
128'h00000000000000000000000000000000, /* 2068 */
128'h00000000000000000000000000000000, /* 2069 */
128'h00000000000000000000000000000000, /* 2070 */
128'h00000000000000000000000000000000, /* 2071 */
128'h00000000000000000000000000000000, /* 2072 */
128'h00000000000000000000000000000000, /* 2073 */
128'h00000000000000000000000000000000, /* 2074 */
128'h00000000000000000000000000000000, /* 2075 */
128'h00000000000000000000000000000000, /* 2076 */
128'h00000000000000000000000000000000, /* 2077 */
128'h00000000000000000000000000000000, /* 2078 */
128'h00000000000000000000000000000000, /* 2079 */
128'h00000000000000000000000000000000, /* 2080 */
128'h00000000000000000000000000000000, /* 2081 */
128'h00000000000000000000000000000000, /* 2082 */
128'h00000000000000000000000000000000, /* 2083 */
128'h00000000000000000000000000000000, /* 2084 */
128'h00000000000000000000000000000000, /* 2085 */
128'h00000000000000000000000000000000, /* 2086 */
128'h00000000000000000000000000000000, /* 2087 */
128'h00000000000000000000000000000000, /* 2088 */
128'h00000000000000000000000000000000, /* 2089 */
128'h00000000000000000000000000000000, /* 2090 */
128'h00000000000000000000000000000000, /* 2091 */
128'h00000000000000000000000000000000, /* 2092 */
128'h00000000000000000000000000000000, /* 2093 */
128'h00000000000000000000000000000000, /* 2094 */
128'h00000000000000000000000000000000, /* 2095 */
128'h00000000000000000000000000000000, /* 2096 */
128'h00000000000000000000000000000000, /* 2097 */
128'h00000000000000000000000000000000, /* 2098 */
128'h00000000000000000000000000000000, /* 2099 */
128'h00000000000000000000000000000000, /* 2100 */
128'h00000000000000000000000000000000, /* 2101 */
128'h00000000000000000000000000000000, /* 2102 */
128'h00000000000000000000000000000000, /* 2103 */
128'h00000000000000000000000000000000, /* 2104 */
128'h00000000000000000000000000000000, /* 2105 */
128'h00000000000000000000000000000000, /* 2106 */
128'h00000000000000000000000000000000, /* 2107 */
128'h00000000000000000000000000000000, /* 2108 */
128'h00000000000000000000000000000000, /* 2109 */
128'h00000000000000000000000000000000, /* 2110 */
128'h00000000000000000000000000000000, /* 2111 */
128'h00000000000000000000000000000000, /* 2112 */
128'h00000000000000000000000000000000, /* 2113 */
128'h00000000000000000000000000000000, /* 2114 */
128'h00000000000000000000000000000000, /* 2115 */
128'h00000000000000000000000000000000, /* 2116 */
128'h00000000000000000000000000000000, /* 2117 */
128'h00000000000000000000000000000000, /* 2118 */
128'h00000000000000000000000000000000, /* 2119 */
128'h00000000000000000000000000000000, /* 2120 */
128'h00000000000000000000000000000000, /* 2121 */
128'h00000000000000000000000000000000, /* 2122 */
128'h00000000000000000000000000000000, /* 2123 */
128'h00000000000000000000000000000000, /* 2124 */
128'h00000000000000000000000000000000, /* 2125 */
128'h00000000000000000000000000000000, /* 2126 */
128'h00000000000000000000000000000000, /* 2127 */
128'h00000000000000000000000000000000, /* 2128 */
128'h00000000000000000000000000000000, /* 2129 */
128'h00000000000000000000000000000000, /* 2130 */
128'h00000000000000000000000000000000, /* 2131 */
128'h00000000000000000000000000000000, /* 2132 */
128'h00000000000000000000000000000000, /* 2133 */
128'h00000000000000000000000000000000, /* 2134 */
128'h00000000000000000000000000000000, /* 2135 */
128'h00000000000000000000000000000000, /* 2136 */
128'h00000000000000000000000000000000, /* 2137 */
128'h00000000000000000000000000000000, /* 2138 */
128'h00000000000000000000000000000000, /* 2139 */
128'h00000000000000000000000000000000, /* 2140 */
128'h00000000000000000000000000000000, /* 2141 */
128'h00000000000000000000000000000000, /* 2142 */
128'h00000000000000000000000000000000, /* 2143 */
128'h00000000000000000000000000000000, /* 2144 */
128'h00000000000000000000000000000000, /* 2145 */
128'h00000000000000000000000000000000, /* 2146 */
128'h00000000000000000000000000000000, /* 2147 */
128'h00000000000000000000000000000000, /* 2148 */
128'h00000000000000000000000000000000, /* 2149 */
128'h00000000000000000000000000000000, /* 2150 */
128'h00000000000000000000000000000000, /* 2151 */
128'h00000000000000000000000000000000, /* 2152 */
128'h00000000000000000000000000000000, /* 2153 */
128'h00000000000000000000000000000000, /* 2154 */
128'h00000000000000000000000000000000, /* 2155 */
128'h00000000000000000000000000000000, /* 2156 */
128'h00000000000000000000000000000000, /* 2157 */
128'h00000000000000000000000000000000, /* 2158 */
128'h00000000000000000000000000000000, /* 2159 */
128'h00000000000000000000000000000000, /* 2160 */
128'h00000000000000000000000000000000, /* 2161 */
128'h00000000000000000000000000000000, /* 2162 */
128'h00000000000000000000000000000000, /* 2163 */
128'h00000000000000000000000000000000, /* 2164 */
128'h00000000000000000000000000000000, /* 2165 */
128'h00000000000000000000000000000000, /* 2166 */
128'h00000000000000000000000000000000, /* 2167 */
128'h00000000000000000000000000000000, /* 2168 */
128'h00000000000000000000000000000000, /* 2169 */
128'h00000000000000000000000000000000, /* 2170 */
128'h00000000000000000000000000000000, /* 2171 */
128'h00000000000000000000000000000000, /* 2172 */
128'h00000000000000000000000000000000, /* 2173 */
128'h00000000000000000000000000000000, /* 2174 */
128'h00000000000000000000000000000000, /* 2175 */
128'h00000000000000000000000000000000, /* 2176 */
128'h00000000000000000000000000000000, /* 2177 */
128'h00000000000000000000000000000000, /* 2178 */
128'h00000000000000000000000000000000, /* 2179 */
128'h00000000000000000000000000000000, /* 2180 */
128'h00000000000000000000000000000000, /* 2181 */
128'h00000000000000000000000000000000, /* 2182 */
128'h00000000000000000000000000000000, /* 2183 */
128'h00000000000000000000000000000000, /* 2184 */
128'h00000000000000000000000000000000, /* 2185 */
128'h00000000000000000000000000000000, /* 2186 */
128'h00000000000000000000000000000000, /* 2187 */
128'h00000000000000000000000000000000, /* 2188 */
128'h00000000000000000000000000000000, /* 2189 */
128'h00000000000000000000000000000000, /* 2190 */
128'h00000000000000000000000000000000, /* 2191 */
128'h00000000000000000000000000000000, /* 2192 */
128'h00000000000000000000000000000000, /* 2193 */
128'h00000000000000000000000000000000, /* 2194 */
128'h00000000000000000000000000000000, /* 2195 */
128'h00000000000000000000000000000000, /* 2196 */
128'h00000000000000000000000000000000, /* 2197 */
128'h00000000000000000000000000000000, /* 2198 */
128'h00000000000000000000000000000000, /* 2199 */
128'h00000000000000000000000000000000, /* 2200 */
128'h00000000000000000000000000000000, /* 2201 */
128'h00000000000000000000000000000000, /* 2202 */
128'h00000000000000000000000000000000, /* 2203 */
128'h00000000000000000000000000000000, /* 2204 */
128'h00000000000000000000000000000000, /* 2205 */
128'h00000000000000000000000000000000, /* 2206 */
128'h00000000000000000000000000000000, /* 2207 */
128'h00000000000000000000000000000000, /* 2208 */
128'h00000000000000000000000000000000, /* 2209 */
128'h00000000000000000000000000000000, /* 2210 */
128'h00000000000000000000000000000000, /* 2211 */
128'h00000000000000000000000000000000, /* 2212 */
128'h00000000000000000000000000000000, /* 2213 */
128'h00000000000000000000000000000000, /* 2214 */
128'h00000000000000000000000000000000, /* 2215 */
128'h00000000000000000000000000000000, /* 2216 */
128'h00000000000000000000000000000000, /* 2217 */
128'h00000000000000000000000000000000, /* 2218 */
128'h00000000000000000000000000000000, /* 2219 */
128'h00000000000000000000000000000000, /* 2220 */
128'h00000000000000000000000000000000, /* 2221 */
128'h00000000000000000000000000000000, /* 2222 */
128'h00000000000000000000000000000000, /* 2223 */
128'h00000000000000000000000000000000, /* 2224 */
128'h00000000000000000000000000000000, /* 2225 */
128'h00000000000000000000000000000000, /* 2226 */
128'h00000000000000000000000000000000, /* 2227 */
128'h00000000000000000000000000000000, /* 2228 */
128'h00000000000000000000000000000000, /* 2229 */
128'h00000000000000000000000000000000, /* 2230 */
128'h00000000000000000000000000000000, /* 2231 */
128'h00000000000000000000000000000000, /* 2232 */
128'h00000000000000000000000000000000, /* 2233 */
128'h00000000000000000000000000000000, /* 2234 */
128'h00000000000000000000000000000000, /* 2235 */
128'h00000000000000000000000000000000, /* 2236 */
128'h00000000000000000000000000000000, /* 2237 */
128'h00000000000000000000000000000000, /* 2238 */
128'h00000000000000000000000000000000, /* 2239 */
128'h00000000000000000000000000000000, /* 2240 */
128'h00000000000000000000000000000000, /* 2241 */
128'h00000000000000000000000000000000, /* 2242 */
128'h00000000000000000000000000000000, /* 2243 */
128'h00000000000000000000000000000000, /* 2244 */
128'h00000000000000000000000000000000, /* 2245 */
128'h00000000000000000000000000000000, /* 2246 */
128'h00000000000000000000000000000000, /* 2247 */
128'h00000000000000000000000000000000, /* 2248 */
128'h00000000000000000000000000000000, /* 2249 */
128'h00000000000000000000000000000000, /* 2250 */
128'h00000000000000000000000000000000, /* 2251 */
128'h00000000000000000000000000000000, /* 2252 */
128'h00000000000000000000000000000000, /* 2253 */
128'h00000000000000000000000000000000, /* 2254 */
128'h00000000000000000000000000000000, /* 2255 */
128'h00000000000000000000000000000000, /* 2256 */
128'h00000000000000000000000000000000, /* 2257 */
128'h00000000000000000000000000000000, /* 2258 */
128'h00000000000000000000000000000000, /* 2259 */
128'h00000000000000000000000000000000, /* 2260 */
128'h00000000000000000000000000000000, /* 2261 */
128'h00000000000000000000000000000000, /* 2262 */
128'h00000000000000000000000000000000, /* 2263 */
128'h00000000000000000000000000000000, /* 2264 */
128'h00000000000000000000000000000000, /* 2265 */
128'h00000000000000000000000000000000, /* 2266 */
128'h00000000000000000000000000000000, /* 2267 */
128'h00000000000000000000000000000000, /* 2268 */
128'h00000000000000000000000000000000, /* 2269 */
128'h00000000000000000000000000000000, /* 2270 */
128'h00000000000000000000000000000000, /* 2271 */
128'h00000000000000000000000000000000, /* 2272 */
128'h00000000000000000000000000000000, /* 2273 */
128'h00000000000000000000000000000000, /* 2274 */
128'h00000000000000000000000000000000, /* 2275 */
128'h00000000000000000000000000000000, /* 2276 */
128'h00000000000000000000000000000000, /* 2277 */
128'h00000000000000000000000000000000, /* 2278 */
128'h00000000000000000000000000000000, /* 2279 */
128'h00000000000000000000000000000000, /* 2280 */
128'h00000000000000000000000000000000, /* 2281 */
128'h00000000000000000000000000000000, /* 2282 */
128'h00000000000000000000000000000000, /* 2283 */
128'h00000000000000000000000000000000, /* 2284 */
128'h00000000000000000000000000000000, /* 2285 */
128'h00000000000000000000000000000000, /* 2286 */
128'h00000000000000000000000000000000, /* 2287 */
128'h00000000000000000000000000000000, /* 2288 */
128'h00000000000000000000000000000000, /* 2289 */
128'h00000000000000000000000000000000, /* 2290 */
128'h00000000000000000000000000000000, /* 2291 */
128'h00000000000000000000000000000000, /* 2292 */
128'h00000000000000000000000000000000, /* 2293 */
128'h00000000000000000000000000000000, /* 2294 */
128'h00000000000000000000000000000000, /* 2295 */
128'h00000000000000000000000000000000, /* 2296 */
128'h00000000000000000000000000000000, /* 2297 */
128'h00000000000000000000000000000000, /* 2298 */
128'h00000000000000000000000000000000, /* 2299 */
128'h00000000000000000000000000000000, /* 2300 */
128'h00000000000000000000000000000000, /* 2301 */
128'h00000000000000000000000000000000, /* 2302 */
128'h00000000000000000000000000000000, /* 2303 */
128'h00000000000000000000000000000000, /* 2304 */
128'h00000000000000000000000000000000, /* 2305 */
128'h00000000000000000000000000000000, /* 2306 */
128'h00000000000000000000000000000000, /* 2307 */
128'h00000000000000000000000000000000, /* 2308 */
128'h00000000000000000000000000000000, /* 2309 */
128'h00000000000000000000000000000000, /* 2310 */
128'h00000000000000000000000000000000, /* 2311 */
128'h00000000000000000000000000000000, /* 2312 */
128'h00000000000000000000000000000000, /* 2313 */
128'h00000000000000000000000000000000, /* 2314 */
128'h00000000000000000000000000000000, /* 2315 */
128'h00000000000000000000000000000000, /* 2316 */
128'h00000000000000000000000000000000, /* 2317 */
128'h00000000000000000000000000000000, /* 2318 */
128'h00000000000000000000000000000000, /* 2319 */
128'h00000000000000000000000000000000, /* 2320 */
128'h00000000000000000000000000000000, /* 2321 */
128'h00000000000000000000000000000000, /* 2322 */
128'h00000000000000000000000000000000, /* 2323 */
128'h00000000000000000000000000000000, /* 2324 */
128'h00000000000000000000000000000000, /* 2325 */
128'h00000000000000000000000000000000, /* 2326 */
128'h00000000000000000000000000000000, /* 2327 */
128'h00000000000000000000000000000000, /* 2328 */
128'h00000000000000000000000000000000, /* 2329 */
128'h00000000000000000000000000000000, /* 2330 */
128'h00000000000000000000000000000000, /* 2331 */
128'h00000000000000000000000000000000, /* 2332 */
128'h00000000000000000000000000000000, /* 2333 */
128'h00000000000000000000000000000000, /* 2334 */
128'h00000000000000000000000000000000, /* 2335 */
128'h00000000000000000000000000000000, /* 2336 */
128'h00000000000000000000000000000000, /* 2337 */
128'h00000000000000000000000000000000, /* 2338 */
128'h00000000000000000000000000000000, /* 2339 */
128'h00000000000000000000000000000000, /* 2340 */
128'h00000000000000000000000000000000, /* 2341 */
128'h00000000000000000000000000000000, /* 2342 */
128'h00000000000000000000000000000000, /* 2343 */
128'h00000000000000000000000000000000, /* 2344 */
128'h00000000000000000000000000000000, /* 2345 */
128'h00000000000000000000000000000000, /* 2346 */
128'h00000000000000000000000000000000, /* 2347 */
128'h00000000000000000000000000000000, /* 2348 */
128'h00000000000000000000000000000000, /* 2349 */
128'h00000000000000000000000000000000, /* 2350 */
128'h00000000000000000000000000000000, /* 2351 */
128'h00000000000000000000000000000000, /* 2352 */
128'h00000000000000000000000000000000, /* 2353 */
128'h00000000000000000000000000000000, /* 2354 */
128'h00000000000000000000000000000000, /* 2355 */
128'h00000000000000000000000000000000, /* 2356 */
128'h00000000000000000000000000000000, /* 2357 */
128'h00000000000000000000000000000000, /* 2358 */
128'h00000000000000000000000000000000, /* 2359 */
128'h00000000000000000000000000000000, /* 2360 */
128'h00000000000000000000000000000000, /* 2361 */
128'h00000000000000000000000000000000, /* 2362 */
128'h00000000000000000000000000000000, /* 2363 */
128'h00000000000000000000000000000000, /* 2364 */
128'h00000000000000000000000000000000, /* 2365 */
128'h00000000000000000000000000000000, /* 2366 */
128'h00000000000000000000000000000000, /* 2367 */
128'h00000000000000000000000000000000, /* 2368 */
128'h00000000000000000000000000000000, /* 2369 */
128'h00000000000000000000000000000000, /* 2370 */
128'h00000000000000000000000000000000, /* 2371 */
128'h00000000000000000000000000000000, /* 2372 */
128'h00000000000000000000000000000000, /* 2373 */
128'h00000000000000000000000000000000, /* 2374 */
128'h00000000000000000000000000000000, /* 2375 */
128'h00000000000000000000000000000000, /* 2376 */
128'h00000000000000000000000000000000, /* 2377 */
128'h00000000000000000000000000000000, /* 2378 */
128'h00000000000000000000000000000000, /* 2379 */
128'h00000000000000000000000000000000, /* 2380 */
128'h00000000000000000000000000000000, /* 2381 */
128'h00000000000000000000000000000000, /* 2382 */
128'h00000000000000000000000000000000, /* 2383 */
128'h00000000000000000000000000000000, /* 2384 */
128'h00000000000000000000000000000000, /* 2385 */
128'h00000000000000000000000000000000, /* 2386 */
128'h00000000000000000000000000000000, /* 2387 */
128'h00000000000000000000000000000000, /* 2388 */
128'h00000000000000000000000000000000, /* 2389 */
128'h00000000000000000000000000000000, /* 2390 */
128'h00000000000000000000000000000000, /* 2391 */
128'h00000000000000000000000000000000, /* 2392 */
128'h00000000000000000000000000000000, /* 2393 */
128'h00000000000000000000000000000000, /* 2394 */
128'h00000000000000000000000000000000, /* 2395 */
128'h00000000000000000000000000000000, /* 2396 */
128'h00000000000000000000000000000000, /* 2397 */
128'h00000000000000000000000000000000, /* 2398 */
128'h00000000000000000000000000000000, /* 2399 */
128'h00000000000000000000000000000000, /* 2400 */
128'h00000000000000000000000000000000, /* 2401 */
128'h00000000000000000000000000000000, /* 2402 */
128'h00000000000000000000000000000000, /* 2403 */
128'h00000000000000000000000000000000, /* 2404 */
128'h00000000000000000000000000000000, /* 2405 */
128'h00000000000000000000000000000000, /* 2406 */
128'h00000000000000000000000000000000, /* 2407 */
128'h00000000000000000000000000000000, /* 2408 */
128'h00000000000000000000000000000000, /* 2409 */
128'h00000000000000000000000000000000, /* 2410 */
128'h00000000000000000000000000000000, /* 2411 */
128'h00000000000000000000000000000000, /* 2412 */
128'h00000000000000000000000000000000, /* 2413 */
128'h00000000000000000000000000000000, /* 2414 */
128'h00000000000000000000000000000000, /* 2415 */
128'h00000000000000000000000000000000, /* 2416 */
128'h00000000000000000000000000000000, /* 2417 */
128'h00000000000000000000000000000000, /* 2418 */
128'h00000000000000000000000000000000, /* 2419 */
128'h00000000000000000000000000000000, /* 2420 */
128'h00000000000000000000000000000000, /* 2421 */
128'h00000000000000000000000000000000, /* 2422 */
128'h00000000000000000000000000000000, /* 2423 */
128'h00000000000000000000000000000000, /* 2424 */
128'h00000000000000000000000000000000, /* 2425 */
128'h00000000000000000000000000000000, /* 2426 */
128'h00000000000000000000000000000000, /* 2427 */
128'h00000000000000000000000000000000, /* 2428 */
128'h00000000000000000000000000000000, /* 2429 */
128'h00000000000000000000000000000000, /* 2430 */
128'h00000000000000000000000000000000, /* 2431 */
128'h00000000000000000000000000000000, /* 2432 */
128'h00000000000000000000000000000000, /* 2433 */
128'h00000000000000000000000000000000, /* 2434 */
128'h00000000000000000000000000000000, /* 2435 */
128'h00000000000000000000000000000000, /* 2436 */
128'h00000000000000000000000000000000, /* 2437 */
128'h00000000000000000000000000000000, /* 2438 */
128'h00000000000000000000000000000000, /* 2439 */
128'h00000000000000000000000000000000, /* 2440 */
128'h00000000000000000000000000000000, /* 2441 */
128'h00000000000000000000000000000000, /* 2442 */
128'h00000000000000000000000000000000, /* 2443 */
128'h00000000000000000000000000000000, /* 2444 */
128'h00000000000000000000000000000000, /* 2445 */
128'h00000000000000000000000000000000, /* 2446 */
128'h00000000000000000000000000000000, /* 2447 */
128'h00000000000000000000000000000000, /* 2448 */
128'h00000000000000000000000000000000, /* 2449 */
128'h00000000000000000000000000000000, /* 2450 */
128'h00000000000000000000000000000000, /* 2451 */
128'h00000000000000000000000000000000, /* 2452 */
128'h00000000000000000000000000000000, /* 2453 */
128'h00000000000000000000000000000000, /* 2454 */
128'h00000000000000000000000000000000, /* 2455 */
128'h00000000000000000000000000000000, /* 2456 */
128'h00000000000000000000000000000000, /* 2457 */
128'h00000000000000000000000000000000, /* 2458 */
128'h00000000000000000000000000000000, /* 2459 */
128'h00000000000000000000000000000000, /* 2460 */
128'h00000000000000000000000000000000, /* 2461 */
128'h00000000000000000000000000000000, /* 2462 */
128'h00000000000000000000000000000000, /* 2463 */
128'h00000000000000000000000000000000, /* 2464 */
128'h00000000000000000000000000000000, /* 2465 */
128'h00000000000000000000000000000000, /* 2466 */
128'h00000000000000000000000000000000, /* 2467 */
128'h00000000000000000000000000000000, /* 2468 */
128'h00000000000000000000000000000000, /* 2469 */
128'h00000000000000000000000000000000, /* 2470 */
128'h00000000000000000000000000000000, /* 2471 */
128'h00000000000000000000000000000000, /* 2472 */
128'h00000000000000000000000000000000, /* 2473 */
128'h00000000000000000000000000000000, /* 2474 */
128'h00000000000000000000000000000000, /* 2475 */
128'h00000000000000000000000000000000, /* 2476 */
128'h00000000000000000000000000000000, /* 2477 */
128'h00000000000000000000000000000000, /* 2478 */
128'h00000000000000000000000000000000, /* 2479 */
128'h00000000000000000000000000000000, /* 2480 */
128'h00000000000000000000000000000000, /* 2481 */
128'h00000000000000000000000000000000, /* 2482 */
128'h00000000000000000000000000000000, /* 2483 */
128'h00000000000000000000000000000000, /* 2484 */
128'h00000000000000000000000000000000, /* 2485 */
128'h00000000000000000000000000000000, /* 2486 */
128'h00000000000000000000000000000000, /* 2487 */
128'h00000000000000000000000000000000, /* 2488 */
128'h00000000000000000000000000000000, /* 2489 */
128'h00000000000000000000000000000000, /* 2490 */
128'h00000000000000000000000000000000, /* 2491 */
128'h00000000000000000000000000000000, /* 2492 */
128'h00000000000000000000000000000000, /* 2493 */
128'h00000000000000000000000000000000, /* 2494 */
128'h00000000000000000000000000000000, /* 2495 */
128'h00000000000000000000000000000000, /* 2496 */
128'h00000000000000000000000000000000, /* 2497 */
128'h00000000000000000000000000000000, /* 2498 */
128'h00000000000000000000000000000000, /* 2499 */
128'h00000000000000000000000000000000, /* 2500 */
128'h00000000000000000000000000000000, /* 2501 */
128'h00000000000000000000000000000000, /* 2502 */
128'h00000000000000000000000000000000, /* 2503 */
128'h00000000000000000000000000000000, /* 2504 */
128'h00000000000000000000000000000000, /* 2505 */
128'h00000000000000000000000000000000, /* 2506 */
128'h00000000000000000000000000000000, /* 2507 */
128'h00000000000000000000000000000000, /* 2508 */
128'h00000000000000000000000000000000, /* 2509 */
128'h00000000000000000000000000000000, /* 2510 */
128'h00000000000000000000000000000000, /* 2511 */
128'h00000000000000000000000000000000, /* 2512 */
128'h00000000000000000000000000000000, /* 2513 */
128'h00000000000000000000000000000000, /* 2514 */
128'h00000000000000000000000000000000, /* 2515 */
128'h00000000000000000000000000000000, /* 2516 */
128'h00000000000000000000000000000000, /* 2517 */
128'h00000000000000000000000000000000, /* 2518 */
128'h00000000000000000000000000000000, /* 2519 */
128'h00000000000000000000000000000000, /* 2520 */
128'h00000000000000000000000000000000, /* 2521 */
128'h00000000000000000000000000000000, /* 2522 */
128'h00000000000000000000000000000000, /* 2523 */
128'h00000000000000000000000000000000, /* 2524 */
128'h00000000000000000000000000000000, /* 2525 */
128'h00000000000000000000000000000000, /* 2526 */
128'h00000000000000000000000000000000, /* 2527 */
128'h00000000000000000000000000000000, /* 2528 */
128'h00000000000000000000000000000000, /* 2529 */
128'h00000000000000000000000000000000, /* 2530 */
128'h00000000000000000000000000000000, /* 2531 */
128'h00000000000000000000000000000000, /* 2532 */
128'h00000000000000000000000000000000, /* 2533 */
128'h00000000000000000000000000000000, /* 2534 */
128'h00000000000000000000000000000000, /* 2535 */
128'h00000000000000000000000000000000, /* 2536 */
128'h00000000000000000000000000000000, /* 2537 */
128'h00000000000000000000000000000000, /* 2538 */
128'h00000000000000000000000000000000, /* 2539 */
128'h00000000000000000000000000000000, /* 2540 */
128'h00000000000000000000000000000000, /* 2541 */
128'h00000000000000000000000000000000, /* 2542 */
128'h00000000000000000000000000000000, /* 2543 */
128'h00000000000000000000000000000000, /* 2544 */
128'h00000000000000000000000000000000, /* 2545 */
128'h00000000000000000000000000000000, /* 2546 */
128'h00000000000000000000000000000000, /* 2547 */
128'h00000000000000000000000000000000, /* 2548 */
128'h00000000000000000000000000000000, /* 2549 */
128'h00000000000000000000000000000000, /* 2550 */
128'h00000000000000000000000000000000, /* 2551 */
128'h00000000000000000000000000000000, /* 2552 */
128'h00000000000000000000000000000000, /* 2553 */
128'h00000000000000000000000000000000, /* 2554 */
128'h00000000000000000000000000000000, /* 2555 */
128'h00000000000000000000000000000000, /* 2556 */
128'h00000000000000000000000000000000, /* 2557 */
128'h00000000000000000000000000000000, /* 2558 */
128'h00000000000000000000000000000000, /* 2559 */
128'h00000000000000000000000000000000, /* 2560 */
128'h00000000000000000000000000000000, /* 2561 */
128'h00000000000000000000000000000000, /* 2562 */
128'h00000000000000000000000000000000, /* 2563 */
128'h00000000000000000000000000000000, /* 2564 */
128'h00000000000000000000000000000000, /* 2565 */
128'h00000000000000000000000000000000, /* 2566 */
128'h00000000000000000000000000000000, /* 2567 */
128'h00000000000000000000000000000000, /* 2568 */
128'h00000000000000000000000000000000, /* 2569 */
128'h00000000000000000000000000000000, /* 2570 */
128'h00000000000000000000000000000000, /* 2571 */
128'h00000000000000000000000000000000, /* 2572 */
128'h00000000000000000000000000000000, /* 2573 */
128'h00000000000000000000000000000000, /* 2574 */
128'h00000000000000000000000000000000, /* 2575 */
128'h00000000000000000000000000000000, /* 2576 */
128'h00000000000000000000000000000000, /* 2577 */
128'h00000000000000000000000000000000, /* 2578 */
128'h00000000000000000000000000000000, /* 2579 */
128'h00000000000000000000000000000000, /* 2580 */
128'h00000000000000000000000000000000, /* 2581 */
128'h00000000000000000000000000000000, /* 2582 */
128'h00000000000000000000000000000000, /* 2583 */
128'h00000000000000000000000000000000, /* 2584 */
128'h00000000000000000000000000000000, /* 2585 */
128'h00000000000000000000000000000000, /* 2586 */
128'h00000000000000000000000000000000, /* 2587 */
128'h00000000000000000000000000000000, /* 2588 */
128'h00000000000000000000000000000000, /* 2589 */
128'h00000000000000000000000000000000, /* 2590 */
128'h00000000000000000000000000000000, /* 2591 */
128'h00000000000000000000000000000000, /* 2592 */
128'h00000000000000000000000000000000, /* 2593 */
128'h00000000000000000000000000000000, /* 2594 */
128'h00000000000000000000000000000000, /* 2595 */
128'h00000000000000000000000000000000, /* 2596 */
128'h00000000000000000000000000000000, /* 2597 */
128'h00000000000000000000000000000000, /* 2598 */
128'h00000000000000000000000000000000, /* 2599 */
128'h00000000000000000000000000000000, /* 2600 */
128'h00000000000000000000000000000000, /* 2601 */
128'h00000000000000000000000000000000, /* 2602 */
128'h00000000000000000000000000000000, /* 2603 */
128'h00000000000000000000000000000000, /* 2604 */
128'h00000000000000000000000000000000, /* 2605 */
128'h00000000000000000000000000000000, /* 2606 */
128'h00000000000000000000000000000000, /* 2607 */
128'h00000000000000000000000000000000, /* 2608 */
128'h00000000000000000000000000000000, /* 2609 */
128'h00000000000000000000000000000000, /* 2610 */
128'h00000000000000000000000000000000, /* 2611 */
128'h00000000000000000000000000000000, /* 2612 */
128'h00000000000000000000000000000000, /* 2613 */
128'h00000000000000000000000000000000, /* 2614 */
128'h00000000000000000000000000000000, /* 2615 */
128'h00000000000000000000000000000000, /* 2616 */
128'h00000000000000000000000000000000, /* 2617 */
128'h00000000000000000000000000000000, /* 2618 */
128'h00000000000000000000000000000000, /* 2619 */
128'h00000000000000000000000000000000, /* 2620 */
128'h00000000000000000000000000000000, /* 2621 */
128'h00000000000000000000000000000000, /* 2622 */
128'h00000000000000000000000000000000, /* 2623 */
128'h00000000000000000000000000000000, /* 2624 */
128'h00000000000000000000000000000000, /* 2625 */
128'h00000000000000000000000000000000, /* 2626 */
128'h00000000000000000000000000000000, /* 2627 */
128'h00000000000000000000000000000000, /* 2628 */
128'h00000000000000000000000000000000, /* 2629 */
128'h00000000000000000000000000000000, /* 2630 */
128'h00000000000000000000000000000000, /* 2631 */
128'h00000000000000000000000000000000, /* 2632 */
128'h00000000000000000000000000000000, /* 2633 */
128'h00000000000000000000000000000000, /* 2634 */
128'h00000000000000000000000000000000, /* 2635 */
128'h00000000000000000000000000000000, /* 2636 */
128'h00000000000000000000000000000000, /* 2637 */
128'h00000000000000000000000000000000, /* 2638 */
128'h00000000000000000000000000000000, /* 2639 */
128'h00000000000000000000000000000000, /* 2640 */
128'h00000000000000000000000000000000, /* 2641 */
128'h00000000000000000000000000000000, /* 2642 */
128'h00000000000000000000000000000000, /* 2643 */
128'h00000000000000000000000000000000, /* 2644 */
128'h00000000000000000000000000000000, /* 2645 */
128'h00000000000000000000000000000000, /* 2646 */
128'h00000000000000000000000000000000, /* 2647 */
128'h00000000000000000000000000000000, /* 2648 */
128'h00000000000000000000000000000000, /* 2649 */
128'h00000000000000000000000000000000, /* 2650 */
128'h00000000000000000000000000000000, /* 2651 */
128'h00000000000000000000000000000000, /* 2652 */
128'h00000000000000000000000000000000, /* 2653 */
128'h00000000000000000000000000000000, /* 2654 */
128'h00000000000000000000000000000000, /* 2655 */
128'h00000000000000000000000000000000, /* 2656 */
128'h00000000000000000000000000000000, /* 2657 */
128'h00000000000000000000000000000000, /* 2658 */
128'h00000000000000000000000000000000, /* 2659 */
128'h00000000000000000000000000000000, /* 2660 */
128'h00000000000000000000000000000000, /* 2661 */
128'h00000000000000000000000000000000, /* 2662 */
128'h00000000000000000000000000000000, /* 2663 */
128'h00000000000000000000000000000000, /* 2664 */
128'h00000000000000000000000000000000, /* 2665 */
128'h00000000000000000000000000000000, /* 2666 */
128'h00000000000000000000000000000000, /* 2667 */
128'h00000000000000000000000000000000, /* 2668 */
128'h00000000000000000000000000000000, /* 2669 */
128'h00000000000000000000000000000000, /* 2670 */
128'h00000000000000000000000000000000, /* 2671 */
128'h00000000000000000000000000000000, /* 2672 */
128'h00000000000000000000000000000000, /* 2673 */
128'h00000000000000000000000000000000, /* 2674 */
128'h00000000000000000000000000000000, /* 2675 */
128'h00000000000000000000000000000000, /* 2676 */
128'h00000000000000000000000000000000, /* 2677 */
128'h00000000000000000000000000000000, /* 2678 */
128'h00000000000000000000000000000000, /* 2679 */
128'h00000000000000000000000000000000, /* 2680 */
128'h00000000000000000000000000000000, /* 2681 */
128'h00000000000000000000000000000000, /* 2682 */
128'h00000000000000000000000000000000, /* 2683 */
128'h00000000000000000000000000000000, /* 2684 */
128'h00000000000000000000000000000000, /* 2685 */
128'h00000000000000000000000000000000, /* 2686 */
128'h00000000000000000000000000000000, /* 2687 */
128'h00000000000000000000000000000000, /* 2688 */
128'h00000000000000000000000000000000, /* 2689 */
128'h00000000000000000000000000000000, /* 2690 */
128'h00000000000000000000000000000000, /* 2691 */
128'h00000000000000000000000000000000, /* 2692 */
128'h00000000000000000000000000000000, /* 2693 */
128'h00000000000000000000000000000000, /* 2694 */
128'h00000000000000000000000000000000, /* 2695 */
128'h00000000000000000000000000000000, /* 2696 */
128'h00000000000000000000000000000000, /* 2697 */
128'h00000000000000000000000000000000, /* 2698 */
128'h00000000000000000000000000000000, /* 2699 */
128'h00000000000000000000000000000000, /* 2700 */
128'h00000000000000000000000000000000, /* 2701 */
128'h00000000000000000000000000000000, /* 2702 */
128'h00000000000000000000000000000000, /* 2703 */
128'h00000000000000000000000000000000, /* 2704 */
128'h00000000000000000000000000000000, /* 2705 */
128'h00000000000000000000000000000000, /* 2706 */
128'h00000000000000000000000000000000, /* 2707 */
128'h00000000000000000000000000000000, /* 2708 */
128'h00000000000000000000000000000000, /* 2709 */
128'h00000000000000000000000000000000, /* 2710 */
128'h00000000000000000000000000000000, /* 2711 */
128'h00000000000000000000000000000000, /* 2712 */
128'h00000000000000000000000000000000, /* 2713 */
128'h00000000000000000000000000000000, /* 2714 */
128'h00000000000000000000000000000000, /* 2715 */
128'h00000000000000000000000000000000, /* 2716 */
128'h00000000000000000000000000000000, /* 2717 */
128'h00000000000000000000000000000000, /* 2718 */
128'h00000000000000000000000000000000, /* 2719 */
128'h00000000000000000000000000000000, /* 2720 */
128'h00000000000000000000000000000000, /* 2721 */
128'h00000000000000000000000000000000, /* 2722 */
128'h00000000000000000000000000000000, /* 2723 */
128'h00000000000000000000000000000000, /* 2724 */
128'h00000000000000000000000000000000, /* 2725 */
128'h00000000000000000000000000000000, /* 2726 */
128'h00000000000000000000000000000000, /* 2727 */
128'h00000000000000000000000000000000, /* 2728 */
128'h00000000000000000000000000000000, /* 2729 */
128'h00000000000000000000000000000000, /* 2730 */
128'h00000000000000000000000000000000, /* 2731 */
128'h00000000000000000000000000000000, /* 2732 */
128'h00000000000000000000000000000000, /* 2733 */
128'h00000000000000000000000000000000, /* 2734 */
128'h00000000000000000000000000000000, /* 2735 */
128'h00000000000000000000000000000000, /* 2736 */
128'h00000000000000000000000000000000, /* 2737 */
128'h00000000000000000000000000000000, /* 2738 */
128'h00000000000000000000000000000000, /* 2739 */
128'h00000000000000000000000000000000, /* 2740 */
128'h00000000000000000000000000000000, /* 2741 */
128'h00000000000000000000000000000000, /* 2742 */
128'h00000000000000000000000000000000, /* 2743 */
128'h00000000000000000000000000000000, /* 2744 */
128'h00000000000000000000000000000000, /* 2745 */
128'h00000000000000000000000000000000, /* 2746 */
128'h00000000000000000000000000000000, /* 2747 */
128'h00000000000000000000000000000000, /* 2748 */
128'h00000000000000000000000000000000, /* 2749 */
128'h00000000000000000000000000000000, /* 2750 */
128'h00000000000000000000000000000000, /* 2751 */
128'h00000000000000000000000000000000, /* 2752 */
128'h00000000000000000000000000000000, /* 2753 */
128'h00000000000000000000000000000000, /* 2754 */
128'h00000000000000000000000000000000, /* 2755 */
128'h00000000000000000000000000000000, /* 2756 */
128'h00000000000000000000000000000000, /* 2757 */
128'h00000000000000000000000000000000, /* 2758 */
128'h00000000000000000000000000000000, /* 2759 */
128'h00000000000000000000000000000000, /* 2760 */
128'h00000000000000000000000000000000, /* 2761 */
128'h00000000000000000000000000000000, /* 2762 */
128'h00000000000000000000000000000000, /* 2763 */
128'h00000000000000000000000000000000, /* 2764 */
128'h00000000000000000000000000000000, /* 2765 */
128'h00000000000000000000000000000000, /* 2766 */
128'h00000000000000000000000000000000, /* 2767 */
128'h00000000000000000000000000000000, /* 2768 */
128'h00000000000000000000000000000000, /* 2769 */
128'h00000000000000000000000000000000, /* 2770 */
128'h00000000000000000000000000000000, /* 2771 */
128'h00000000000000000000000000000000, /* 2772 */
128'h00000000000000000000000000000000, /* 2773 */
128'h00000000000000000000000000000000, /* 2774 */
128'h00000000000000000000000000000000, /* 2775 */
128'h00000000000000000000000000000000, /* 2776 */
128'h00000000000000000000000000000000, /* 2777 */
128'h00000000000000000000000000000000, /* 2778 */
128'h00000000000000000000000000000000, /* 2779 */
128'h00000000000000000000000000000000, /* 2780 */
128'h00000000000000000000000000000000, /* 2781 */
128'h00000000000000000000000000000000, /* 2782 */
128'h00000000000000000000000000000000, /* 2783 */
128'h00000000000000000000000000000000, /* 2784 */
128'h00000000000000000000000000000000, /* 2785 */
128'h00000000000000000000000000000000, /* 2786 */
128'h00000000000000000000000000000000, /* 2787 */
128'h00000000000000000000000000000000, /* 2788 */
128'h00000000000000000000000000000000, /* 2789 */
128'h00000000000000000000000000000000, /* 2790 */
128'h00000000000000000000000000000000, /* 2791 */
128'h00000000000000000000000000000000, /* 2792 */
128'h00000000000000000000000000000000, /* 2793 */
128'h00000000000000000000000000000000, /* 2794 */
128'h00000000000000000000000000000000, /* 2795 */
128'h00000000000000000000000000000000, /* 2796 */
128'h00000000000000000000000000000000, /* 2797 */
128'h00000000000000000000000000000000, /* 2798 */
128'h00000000000000000000000000000000, /* 2799 */
128'h00000000000000000000000000000000, /* 2800 */
128'h00000000000000000000000000000000, /* 2801 */
128'h00000000000000000000000000000000, /* 2802 */
128'h00000000000000000000000000000000, /* 2803 */
128'h00000000000000000000000000000000, /* 2804 */
128'h00000000000000000000000000000000, /* 2805 */
128'h00000000000000000000000000000000, /* 2806 */
128'h00000000000000000000000000000000, /* 2807 */
128'h00000000000000000000000000000000, /* 2808 */
128'h00000000000000000000000000000000, /* 2809 */
128'h00000000000000000000000000000000, /* 2810 */
128'h00000000000000000000000000000000, /* 2811 */
128'h00000000000000000000000000000000, /* 2812 */
128'h00000000000000000000000000000000, /* 2813 */
128'h00000000000000000000000000000000, /* 2814 */
128'h00000000000000000000000000000000, /* 2815 */
128'h00000000000000000000000000000000, /* 2816 */
128'h00000000000000000000000000000000, /* 2817 */
128'h00000000000000000000000000000000, /* 2818 */
128'h00000000000000000000000000000000, /* 2819 */
128'h00000000000000000000000000000000, /* 2820 */
128'h00000000000000000000000000000000, /* 2821 */
128'h00000000000000000000000000000000, /* 2822 */
128'h00000000000000000000000000000000, /* 2823 */
128'h00000000000000000000000000000000, /* 2824 */
128'h00000000000000000000000000000000, /* 2825 */
128'h00000000000000000000000000000000, /* 2826 */
128'h00000000000000000000000000000000, /* 2827 */
128'h00000000000000000000000000000000, /* 2828 */
128'h00000000000000000000000000000000, /* 2829 */
128'h00000000000000000000000000000000, /* 2830 */
128'h00000000000000000000000000000000, /* 2831 */
128'h00000000000000000000000000000000, /* 2832 */
128'h00000000000000000000000000000000, /* 2833 */
128'h00000000000000000000000000000000, /* 2834 */
128'h00000000000000000000000000000000, /* 2835 */
128'h00000000000000000000000000000000, /* 2836 */
128'h00000000000000000000000000000000, /* 2837 */
128'h00000000000000000000000000000000, /* 2838 */
128'h00000000000000000000000000000000, /* 2839 */
128'h00000000000000000000000000000000, /* 2840 */
128'h00000000000000000000000000000000, /* 2841 */
128'h00000000000000000000000000000000, /* 2842 */
128'h00000000000000000000000000000000, /* 2843 */
128'h00000000000000000000000000000000, /* 2844 */
128'h00000000000000000000000000000000, /* 2845 */
128'h00000000000000000000000000000000, /* 2846 */
128'h00000000000000000000000000000000, /* 2847 */
128'h00000000000000000000000000000000, /* 2848 */
128'h00000000000000000000000000000000, /* 2849 */
128'h00000000000000000000000000000000, /* 2850 */
128'h00000000000000000000000000000000, /* 2851 */
128'h00000000000000000000000000000000, /* 2852 */
128'h00000000000000000000000000000000, /* 2853 */
128'h00000000000000000000000000000000, /* 2854 */
128'h00000000000000000000000000000000, /* 2855 */
128'h00000000000000000000000000000000, /* 2856 */
128'h00000000000000000000000000000000, /* 2857 */
128'h00000000000000000000000000000000, /* 2858 */
128'h00000000000000000000000000000000, /* 2859 */
128'h00000000000000000000000000000000, /* 2860 */
128'h00000000000000000000000000000000, /* 2861 */
128'h00000000000000000000000000000000, /* 2862 */
128'h00000000000000000000000000000000, /* 2863 */
128'h00000000000000000000000000000000, /* 2864 */
128'h00000000000000000000000000000000, /* 2865 */
128'h00000000000000000000000000000000, /* 2866 */
128'h00000000000000000000000000000000, /* 2867 */
128'h00000000000000000000000000000000, /* 2868 */
128'h00000000000000000000000000000000, /* 2869 */
128'h00000000000000000000000000000000, /* 2870 */
128'h00000000000000000000000000000000, /* 2871 */
128'h00000000000000000000000000000000, /* 2872 */
128'h00000000000000000000000000000000, /* 2873 */
128'h00000000000000000000000000000000, /* 2874 */
128'h00000000000000000000000000000000, /* 2875 */
128'h00000000000000000000000000000000, /* 2876 */
128'h00000000000000000000000000000000, /* 2877 */
128'h00000000000000000000000000000000, /* 2878 */
128'h00000000000000000000000000000000, /* 2879 */
128'h00000000000000000000000000000000, /* 2880 */
128'h00000000000000000000000000000000, /* 2881 */
128'h00000000000000000000000000000000, /* 2882 */
128'h00000000000000000000000000000000, /* 2883 */
128'h00000000000000000000000000000000, /* 2884 */
128'h00000000000000000000000000000000, /* 2885 */
128'h00000000000000000000000000000000, /* 2886 */
128'h00000000000000000000000000000000, /* 2887 */
128'h00000000000000000000000000000000, /* 2888 */
128'h00000000000000000000000000000000, /* 2889 */
128'h00000000000000000000000000000000, /* 2890 */
128'h00000000000000000000000000000000, /* 2891 */
128'h00000000000000000000000000000000, /* 2892 */
128'h00000000000000000000000000000000, /* 2893 */
128'h00000000000000000000000000000000, /* 2894 */
128'h00000000000000000000000000000000, /* 2895 */
128'h00000000000000000000000000000000, /* 2896 */
128'h00000000000000000000000000000000, /* 2897 */
128'h00000000000000000000000000000000, /* 2898 */
128'h00000000000000000000000000000000, /* 2899 */
128'h00000000000000000000000000000000, /* 2900 */
128'h00000000000000000000000000000000, /* 2901 */
128'h00000000000000000000000000000000, /* 2902 */
128'h00000000000000000000000000000000, /* 2903 */
128'h00000000000000000000000000000000, /* 2904 */
128'h00000000000000000000000000000000, /* 2905 */
128'h00000000000000000000000000000000, /* 2906 */
128'h00000000000000000000000000000000, /* 2907 */
128'h00000000000000000000000000000000, /* 2908 */
128'h00000000000000000000000000000000, /* 2909 */
128'h00000000000000000000000000000000, /* 2910 */
128'h00000000000000000000000000000000, /* 2911 */
128'h00000000000000000000000000000000, /* 2912 */
128'h00000000000000000000000000000000, /* 2913 */
128'h00000000000000000000000000000000, /* 2914 */
128'h00000000000000000000000000000000, /* 2915 */
128'h00000000000000000000000000000000, /* 2916 */
128'h00000000000000000000000000000000, /* 2917 */
128'h00000000000000000000000000000000, /* 2918 */
128'h00000000000000000000000000000000, /* 2919 */
128'h00000000000000000000000000000000, /* 2920 */
128'h00000000000000000000000000000000, /* 2921 */
128'h00000000000000000000000000000000, /* 2922 */
128'h00000000000000000000000000000000, /* 2923 */
128'h00000000000000000000000000000000, /* 2924 */
128'h00000000000000000000000000000000, /* 2925 */
128'h00000000000000000000000000000000, /* 2926 */
128'h00000000000000000000000000000000, /* 2927 */
128'h00000000000000000000000000000000, /* 2928 */
128'h00000000000000000000000000000000, /* 2929 */
128'h00000000000000000000000000000000, /* 2930 */
128'h00000000000000000000000000000000, /* 2931 */
128'h00000000000000000000000000000000, /* 2932 */
128'h00000000000000000000000000000000, /* 2933 */
128'h00000000000000000000000000000000, /* 2934 */
128'h00000000000000000000000000000000, /* 2935 */
128'h00000000000000000000000000000000, /* 2936 */
128'h00000000000000000000000000000000, /* 2937 */
128'h00000000000000000000000000000000, /* 2938 */
128'h00000000000000000000000000000000, /* 2939 */
128'h00000000000000000000000000000000, /* 2940 */
128'h00000000000000000000000000000000, /* 2941 */
128'h00000000000000000000000000000000, /* 2942 */
128'h00000000000000000000000000000000, /* 2943 */
128'h00000000000000000000000000000000, /* 2944 */
128'h00000000000000000000000000000000, /* 2945 */
128'h00000000000000000000000000000000, /* 2946 */
128'h00000000000000000000000000000000, /* 2947 */
128'h00000000000000000000000000000000, /* 2948 */
128'h00000000000000000000000000000000, /* 2949 */
128'h00000000000000000000000000000000, /* 2950 */
128'h00000000000000000000000000000000, /* 2951 */
128'h00000000000000000000000000000000, /* 2952 */
128'h00000000000000000000000000000000, /* 2953 */
128'h00000000000000000000000000000000, /* 2954 */
128'h00000000000000000000000000000000, /* 2955 */
128'h00000000000000000000000000000000, /* 2956 */
128'h00000000000000000000000000000000, /* 2957 */
128'h00000000000000000000000000000000, /* 2958 */
128'h00000000000000000000000000000000, /* 2959 */
128'h00000000000000000000000000000000, /* 2960 */
128'h00000000000000000000000000000000, /* 2961 */
128'h00000000000000000000000000000000, /* 2962 */
128'h00000000000000000000000000000000, /* 2963 */
128'h00000000000000000000000000000000, /* 2964 */
128'h00000000000000000000000000000000, /* 2965 */
128'h00000000000000000000000000000000, /* 2966 */
128'h00000000000000000000000000000000, /* 2967 */
128'h00000000000000000000000000000000, /* 2968 */
128'h00000000000000000000000000000000, /* 2969 */
128'h00000000000000000000000000000000, /* 2970 */
128'h00000000000000000000000000000000, /* 2971 */
128'h00000000000000000000000000000000, /* 2972 */
128'h00000000000000000000000000000000, /* 2973 */
128'h00000000000000000000000000000000, /* 2974 */
128'h00000000000000000000000000000000, /* 2975 */
128'h00000000000000000000000000000000, /* 2976 */
128'h00000000000000000000000000000000, /* 2977 */
128'h00000000000000000000000000000000, /* 2978 */
128'h00000000000000000000000000000000, /* 2979 */
128'h00000000000000000000000000000000, /* 2980 */
128'h00000000000000000000000000000000, /* 2981 */
128'h00000000000000000000000000000000, /* 2982 */
128'h00000000000000000000000000000000, /* 2983 */
128'h00000000000000000000000000000000, /* 2984 */
128'h00000000000000000000000000000000, /* 2985 */
128'h00000000000000000000000000000000, /* 2986 */
128'h00000000000000000000000000000000, /* 2987 */
128'h00000000000000000000000000000000, /* 2988 */
128'h00000000000000000000000000000000, /* 2989 */
128'h00000000000000000000000000000000, /* 2990 */
128'h00000000000000000000000000000000, /* 2991 */
128'h00000000000000000000000000000000, /* 2992 */
128'h00000000000000000000000000000000, /* 2993 */
128'h00000000000000000000000000000000, /* 2994 */
128'h00000000000000000000000000000000, /* 2995 */
128'h00000000000000000000000000000000, /* 2996 */
128'h00000000000000000000000000000000, /* 2997 */
128'h00000000000000000000000000000000, /* 2998 */
128'h00000000000000000000000000000000, /* 2999 */
128'h00000000000000000000000000000000, /* 3000 */
128'h00000000000000000000000000000000, /* 3001 */
128'h00000000000000000000000000000000, /* 3002 */
128'h00000000000000000000000000000000, /* 3003 */
128'h00000000000000000000000000000000, /* 3004 */
128'h00000000000000000000000000000000, /* 3005 */
128'h00000000000000000000000000000000, /* 3006 */
128'h00000000000000000000000000000000, /* 3007 */
128'h00000000000000000000000000000000, /* 3008 */
128'h00000000000000000000000000000000, /* 3009 */
128'h00000000000000000000000000000000, /* 3010 */
128'h00000000000000000000000000000000, /* 3011 */
128'h00000000000000000000000000000000, /* 3012 */
128'h00000000000000000000000000000000, /* 3013 */
128'h00000000000000000000000000000000, /* 3014 */
128'h00000000000000000000000000000000, /* 3015 */
128'h00000000000000000000000000000000, /* 3016 */
128'h00000000000000000000000000000000, /* 3017 */
128'h00000000000000000000000000000000, /* 3018 */
128'h00000000000000000000000000000000, /* 3019 */
128'h00000000000000000000000000000000, /* 3020 */
128'h00000000000000000000000000000000, /* 3021 */
128'h00000000000000000000000000000000, /* 3022 */
128'h00000000000000000000000000000000, /* 3023 */
128'h00000000000000000000000000000000, /* 3024 */
128'h00000000000000000000000000000000, /* 3025 */
128'h00000000000000000000000000000000, /* 3026 */
128'h00000000000000000000000000000000, /* 3027 */
128'h00000000000000000000000000000000, /* 3028 */
128'h00000000000000000000000000000000, /* 3029 */
128'h00000000000000000000000000000000, /* 3030 */
128'h00000000000000000000000000000000, /* 3031 */
128'h00000000000000000000000000000000, /* 3032 */
128'h00000000000000000000000000000000, /* 3033 */
128'h00000000000000000000000000000000, /* 3034 */
128'h00000000000000000000000000000000, /* 3035 */
128'h00000000000000000000000000000000, /* 3036 */
128'h00000000000000000000000000000000, /* 3037 */
128'h00000000000000000000000000000000, /* 3038 */
128'h00000000000000000000000000000000, /* 3039 */
128'h00000000000000000000000000000000, /* 3040 */
128'h00000000000000000000000000000000, /* 3041 */
128'h00000000000000000000000000000000, /* 3042 */
128'h00000000000000000000000000000000, /* 3043 */
128'h00000000000000000000000000000000, /* 3044 */
128'h00000000000000000000000000000000, /* 3045 */
128'h00000000000000000000000000000000, /* 3046 */
128'h00000000000000000000000000000000, /* 3047 */
128'h00000000000000000000000000000000, /* 3048 */
128'h00000000000000000000000000000000, /* 3049 */
128'h00000000000000000000000000000000, /* 3050 */
128'h00000000000000000000000000000000, /* 3051 */
128'h00000000000000000000000000000000, /* 3052 */
128'h00000000000000000000000000000000, /* 3053 */
128'h00000000000000000000000000000000, /* 3054 */
128'h00000000000000000000000000000000, /* 3055 */
128'h00000000000000000000000000000000, /* 3056 */
128'h00000000000000000000000000000000, /* 3057 */
128'h00000000000000000000000000000000, /* 3058 */
128'h00000000000000000000000000000000, /* 3059 */
128'h00000000000000000000000000000000, /* 3060 */
128'h00000000000000000000000000000000, /* 3061 */
128'h00000000000000000000000000000000, /* 3062 */
128'h00000000000000000000000000000000, /* 3063 */
128'h00000000000000000000000000000000, /* 3064 */
128'h00000000000000000000000000000000, /* 3065 */
128'h00000000000000000000000000000000, /* 3066 */
128'h00000000000000000000000000000000, /* 3067 */
128'h00000000000000000000000000000000, /* 3068 */
128'h00000000000000000000000000000000, /* 3069 */
128'h00000000000000000000000000000000, /* 3070 */
128'h00000000000000000000000000000000, /* 3071 */
128'h00000000000000000000000000000000, /* 3072 */
128'h00000000000000000000000000000000, /* 3073 */
128'h00000000000000000000000000000000, /* 3074 */
128'h00000000000000000000000000000000, /* 3075 */
128'h00000000000000000000000000000000, /* 3076 */
128'h00000000000000000000000000000000, /* 3077 */
128'h00000000000000000000000000000000, /* 3078 */
128'h00000000000000000000000000000000, /* 3079 */
128'h00000000000000000000000000000000, /* 3080 */
128'h00000000000000000000000000000000, /* 3081 */
128'h00000000000000000000000000000000, /* 3082 */
128'h00000000000000000000000000000000, /* 3083 */
128'h00000000000000000000000000000000, /* 3084 */
128'h00000000000000000000000000000000, /* 3085 */
128'h00000000000000000000000000000000, /* 3086 */
128'h00000000000000000000000000000000, /* 3087 */
128'h00000000000000000000000000000000, /* 3088 */
128'h00000000000000000000000000000000, /* 3089 */
128'h00000000000000000000000000000000, /* 3090 */
128'h00000000000000000000000000000000, /* 3091 */
128'h00000000000000000000000000000000, /* 3092 */
128'h00000000000000000000000000000000, /* 3093 */
128'h00000000000000000000000000000000, /* 3094 */
128'h00000000000000000000000000000000, /* 3095 */
128'h00000000000000000000000000000000, /* 3096 */
128'h00000000000000000000000000000000, /* 3097 */
128'h00000000000000000000000000000000, /* 3098 */
128'h00000000000000000000000000000000, /* 3099 */
128'h00000000000000000000000000000000, /* 3100 */
128'h00000000000000000000000000000000, /* 3101 */
128'h00000000000000000000000000000000, /* 3102 */
128'h00000000000000000000000000000000, /* 3103 */
128'h00000000000000000000000000000000, /* 3104 */
128'h00000000000000000000000000000000, /* 3105 */
128'h00000000000000000000000000000000, /* 3106 */
128'h00000000000000000000000000000000, /* 3107 */
128'h00000000000000000000000000000000, /* 3108 */
128'h00000000000000000000000000000000, /* 3109 */
128'h00000000000000000000000000000000, /* 3110 */
128'h00000000000000000000000000000000, /* 3111 */
128'h00000000000000000000000000000000, /* 3112 */
128'h00000000000000000000000000000000, /* 3113 */
128'h00000000000000000000000000000000, /* 3114 */
128'h00000000000000000000000000000000, /* 3115 */
128'h00000000000000000000000000000000, /* 3116 */
128'h00000000000000000000000000000000, /* 3117 */
128'h00000000000000000000000000000000, /* 3118 */
128'h00000000000000000000000000000000, /* 3119 */
128'h00000000000000000000000000000000, /* 3120 */
128'h00000000000000000000000000000000, /* 3121 */
128'h00000000000000000000000000000000, /* 3122 */
128'h00000000000000000000000000000000, /* 3123 */
128'h00000000000000000000000000000000, /* 3124 */
128'h00000000000000000000000000000000, /* 3125 */
128'h00000000000000000000000000000000, /* 3126 */
128'h00000000000000000000000000000000, /* 3127 */
128'h00000000000000000000000000000000, /* 3128 */
128'h00000000000000000000000000000000, /* 3129 */
128'h00000000000000000000000000000000, /* 3130 */
128'h00000000000000000000000000000000, /* 3131 */
128'h00000000000000000000000000000000, /* 3132 */
128'h00000000000000000000000000000000, /* 3133 */
128'h00000000000000000000000000000000, /* 3134 */
128'h00000000000000000000000000000000, /* 3135 */
128'h00000000000000000000000000000000, /* 3136 */
128'h00000000000000000000000000000000, /* 3137 */
128'h00000000000000000000000000000000, /* 3138 */
128'h00000000000000000000000000000000, /* 3139 */
128'h00000000000000000000000000000000, /* 3140 */
128'h00000000000000000000000000000000, /* 3141 */
128'h00000000000000000000000000000000, /* 3142 */
128'h00000000000000000000000000000000, /* 3143 */
128'h00000000000000000000000000000000, /* 3144 */
128'h00000000000000000000000000000000, /* 3145 */
128'h00000000000000000000000000000000, /* 3146 */
128'h00000000000000000000000000000000, /* 3147 */
128'h00000000000000000000000000000000, /* 3148 */
128'h00000000000000000000000000000000, /* 3149 */
128'h00000000000000000000000000000000, /* 3150 */
128'h00000000000000000000000000000000, /* 3151 */
128'h00000000000000000000000000000000, /* 3152 */
128'h00000000000000000000000000000000, /* 3153 */
128'h00000000000000000000000000000000, /* 3154 */
128'h00000000000000000000000000000000, /* 3155 */
128'h00000000000000000000000000000000, /* 3156 */
128'h00000000000000000000000000000000, /* 3157 */
128'h00000000000000000000000000000000, /* 3158 */
128'h00000000000000000000000000000000, /* 3159 */
128'h00000000000000000000000000000000, /* 3160 */
128'h00000000000000000000000000000000, /* 3161 */
128'h00000000000000000000000000000000, /* 3162 */
128'h00000000000000000000000000000000, /* 3163 */
128'h00000000000000000000000000000000, /* 3164 */
128'h00000000000000000000000000000000, /* 3165 */
128'h00000000000000000000000000000000, /* 3166 */
128'h00000000000000000000000000000000, /* 3167 */
128'h00000000000000000000000000000000, /* 3168 */
128'h00000000000000000000000000000000, /* 3169 */
128'h00000000000000000000000000000000, /* 3170 */
128'h00000000000000000000000000000000, /* 3171 */
128'h00000000000000000000000000000000, /* 3172 */
128'h00000000000000000000000000000000, /* 3173 */
128'h00000000000000000000000000000000, /* 3174 */
128'h00000000000000000000000000000000, /* 3175 */
128'h00000000000000000000000000000000, /* 3176 */
128'h00000000000000000000000000000000, /* 3177 */
128'h00000000000000000000000000000000, /* 3178 */
128'h00000000000000000000000000000000, /* 3179 */
128'h00000000000000000000000000000000, /* 3180 */
128'h00000000000000000000000000000000, /* 3181 */
128'h00000000000000000000000000000000, /* 3182 */
128'h00000000000000000000000000000000, /* 3183 */
128'h00000000000000000000000000000000, /* 3184 */
128'h00000000000000000000000000000000, /* 3185 */
128'h00000000000000000000000000000000, /* 3186 */
128'h00000000000000000000000000000000, /* 3187 */
128'h00000000000000000000000000000000, /* 3188 */
128'h00000000000000000000000000000000, /* 3189 */
128'h00000000000000000000000000000000, /* 3190 */
128'h00000000000000000000000000000000, /* 3191 */
128'h00000000000000000000000000000000, /* 3192 */
128'h00000000000000000000000000000000, /* 3193 */
128'h00000000000000000000000000000000, /* 3194 */
128'h00000000000000000000000000000000, /* 3195 */
128'h00000000000000000000000000000000, /* 3196 */
128'h00000000000000000000000000000000, /* 3197 */
128'h00000000000000000000000000000000, /* 3198 */
128'h00000000000000000000000000000000, /* 3199 */
128'h00000000000000000000000000000000, /* 3200 */
128'h00000000000000000000000000000000, /* 3201 */
128'h00000000000000000000000000000000, /* 3202 */
128'h00000000000000000000000000000000, /* 3203 */
128'h00000000000000000000000000000000, /* 3204 */
128'h00000000000000000000000000000000, /* 3205 */
128'h00000000000000000000000000000000, /* 3206 */
128'h00000000000000000000000000000000, /* 3207 */
128'h00000000000000000000000000000000, /* 3208 */
128'h00000000000000000000000000000000, /* 3209 */
128'h00000000000000000000000000000000, /* 3210 */
128'h00000000000000000000000000000000, /* 3211 */
128'h00000000000000000000000000000000, /* 3212 */
128'h00000000000000000000000000000000, /* 3213 */
128'h00000000000000000000000000000000, /* 3214 */
128'h00000000000000000000000000000000, /* 3215 */
128'h00000000000000000000000000000000, /* 3216 */
128'h00000000000000000000000000000000, /* 3217 */
128'h00000000000000000000000000000000, /* 3218 */
128'h00000000000000000000000000000000, /* 3219 */
128'h00000000000000000000000000000000, /* 3220 */
128'h00000000000000000000000000000000, /* 3221 */
128'h00000000000000000000000000000000, /* 3222 */
128'h00000000000000000000000000000000, /* 3223 */
128'h00000000000000000000000000000000, /* 3224 */
128'h00000000000000000000000000000000, /* 3225 */
128'h00000000000000000000000000000000, /* 3226 */
128'h00000000000000000000000000000000, /* 3227 */
128'h00000000000000000000000000000000, /* 3228 */
128'h00000000000000000000000000000000, /* 3229 */
128'h00000000000000000000000000000000, /* 3230 */
128'h00000000000000000000000000000000, /* 3231 */
128'h00000000000000000000000000000000, /* 3232 */
128'h00000000000000000000000000000000, /* 3233 */
128'h00000000000000000000000000000000, /* 3234 */
128'h00000000000000000000000000000000, /* 3235 */
128'h00000000000000000000000000000000, /* 3236 */
128'h00000000000000000000000000000000, /* 3237 */
128'h00000000000000000000000000000000, /* 3238 */
128'h00000000000000000000000000000000, /* 3239 */
128'h00000000000000000000000000000000, /* 3240 */
128'h00000000000000000000000000000000, /* 3241 */
128'h00000000000000000000000000000000, /* 3242 */
128'h00000000000000000000000000000000, /* 3243 */
128'h00000000000000000000000000000000, /* 3244 */
128'h00000000000000000000000000000000, /* 3245 */
128'h00000000000000000000000000000000, /* 3246 */
128'h00000000000000000000000000000000, /* 3247 */
128'h00000000000000000000000000000000, /* 3248 */
128'h00000000000000000000000000000000, /* 3249 */
128'h00000000000000000000000000000000, /* 3250 */
128'h00000000000000000000000000000000, /* 3251 */
128'h00000000000000000000000000000000, /* 3252 */
128'h00000000000000000000000000000000, /* 3253 */
128'h00000000000000000000000000000000, /* 3254 */
128'h00000000000000000000000000000000, /* 3255 */
128'h00000000000000000000000000000000, /* 3256 */
128'h00000000000000000000000000000000, /* 3257 */
128'h00000000000000000000000000000000, /* 3258 */
128'h00000000000000000000000000000000, /* 3259 */
128'h00000000000000000000000000000000, /* 3260 */
128'h00000000000000000000000000000000, /* 3261 */
128'h00000000000000000000000000000000, /* 3262 */
128'h00000000000000000000000000000000, /* 3263 */
128'h00000000000000000000000000000000, /* 3264 */
128'h00000000000000000000000000000000, /* 3265 */
128'h00000000000000000000000000000000, /* 3266 */
128'h00000000000000000000000000000000, /* 3267 */
128'h00000000000000000000000000000000, /* 3268 */
128'h00000000000000000000000000000000, /* 3269 */
128'h00000000000000000000000000000000, /* 3270 */
128'h00000000000000000000000000000000, /* 3271 */
128'h00000000000000000000000000000000, /* 3272 */
128'h00000000000000000000000000000000, /* 3273 */
128'h00000000000000000000000000000000, /* 3274 */
128'h00000000000000000000000000000000, /* 3275 */
128'h00000000000000000000000000000000, /* 3276 */
128'h00000000000000000000000000000000, /* 3277 */
128'h00000000000000000000000000000000, /* 3278 */
128'h00000000000000000000000000000000, /* 3279 */
128'h00000000000000000000000000000000, /* 3280 */
128'h00000000000000000000000000000000, /* 3281 */
128'h00000000000000000000000000000000, /* 3282 */
128'h00000000000000000000000000000000, /* 3283 */
128'h00000000000000000000000000000000, /* 3284 */
128'h00000000000000000000000000000000, /* 3285 */
128'h00000000000000000000000000000000, /* 3286 */
128'h00000000000000000000000000000000, /* 3287 */
128'h00000000000000000000000000000000, /* 3288 */
128'h00000000000000000000000000000000, /* 3289 */
128'h00000000000000000000000000000000, /* 3290 */
128'h00000000000000000000000000000000, /* 3291 */
128'h00000000000000000000000000000000, /* 3292 */
128'h00000000000000000000000000000000, /* 3293 */
128'h00000000000000000000000000000000, /* 3294 */
128'h00000000000000000000000000000000, /* 3295 */
128'h00000000000000000000000000000000, /* 3296 */
128'h00000000000000000000000000000000, /* 3297 */
128'h00000000000000000000000000000000, /* 3298 */
128'h00000000000000000000000000000000, /* 3299 */
128'h00000000000000000000000000000000, /* 3300 */
128'h00000000000000000000000000000000, /* 3301 */
128'h00000000000000000000000000000000, /* 3302 */
128'h00000000000000000000000000000000, /* 3303 */
128'h00000000000000000000000000000000, /* 3304 */
128'h00000000000000000000000000000000, /* 3305 */
128'h00000000000000000000000000000000, /* 3306 */
128'h00000000000000000000000000000000, /* 3307 */
128'h00000000000000000000000000000000, /* 3308 */
128'h00000000000000000000000000000000, /* 3309 */
128'h00000000000000000000000000000000, /* 3310 */
128'h00000000000000000000000000000000, /* 3311 */
128'h00000000000000000000000000000000, /* 3312 */
128'h00000000000000000000000000000000, /* 3313 */
128'h00000000000000000000000000000000, /* 3314 */
128'h00000000000000000000000000000000, /* 3315 */
128'h00000000000000000000000000000000, /* 3316 */
128'h00000000000000000000000000000000, /* 3317 */
128'h00000000000000000000000000000000, /* 3318 */
128'h00000000000000000000000000000000, /* 3319 */
128'h00000000000000000000000000000000, /* 3320 */
128'h00000000000000000000000000000000, /* 3321 */
128'h00000000000000000000000000000000, /* 3322 */
128'h00000000000000000000000000000000, /* 3323 */
128'h00000000000000000000000000000000, /* 3324 */
128'h00000000000000000000000000000000, /* 3325 */
128'h00000000000000000000000000000000, /* 3326 */
128'h00000000000000000000000000000000, /* 3327 */
128'h00000000000000000000000000000000, /* 3328 */
128'h00000000000000000000000000000000, /* 3329 */
128'h00000000000000000000000000000000, /* 3330 */
128'h00000000000000000000000000000000, /* 3331 */
128'h00000000000000000000000000000000, /* 3332 */
128'h00000000000000000000000000000000, /* 3333 */
128'h00000000000000000000000000000000, /* 3334 */
128'h00000000000000000000000000000000, /* 3335 */
128'h00000000000000000000000000000000, /* 3336 */
128'h00000000000000000000000000000000, /* 3337 */
128'h00000000000000000000000000000000, /* 3338 */
128'h00000000000000000000000000000000, /* 3339 */
128'h00000000000000000000000000000000, /* 3340 */
128'h00000000000000000000000000000000, /* 3341 */
128'h00000000000000000000000000000000, /* 3342 */
128'h00000000000000000000000000000000, /* 3343 */
128'h00000000000000000000000000000000, /* 3344 */
128'h00000000000000000000000000000000, /* 3345 */
128'h00000000000000000000000000000000, /* 3346 */
128'h00000000000000000000000000000000, /* 3347 */
128'h00000000000000000000000000000000, /* 3348 */
128'h00000000000000000000000000000000, /* 3349 */
128'h00000000000000000000000000000000, /* 3350 */
128'h00000000000000000000000000000000, /* 3351 */
128'h00000000000000000000000000000000, /* 3352 */
128'h00000000000000000000000000000000, /* 3353 */
128'h00000000000000000000000000000000, /* 3354 */
128'h00000000000000000000000000000000, /* 3355 */
128'h00000000000000000000000000000000, /* 3356 */
128'h00000000000000000000000000000000, /* 3357 */
128'h00000000000000000000000000000000, /* 3358 */
128'h00000000000000000000000000000000, /* 3359 */
128'h00000000000000000000000000000000, /* 3360 */
128'h00000000000000000000000000000000, /* 3361 */
128'h00000000000000000000000000000000, /* 3362 */
128'h00000000000000000000000000000000, /* 3363 */
128'h00000000000000000000000000000000, /* 3364 */
128'h00000000000000000000000000000000, /* 3365 */
128'h00000000000000000000000000000000, /* 3366 */
128'h00000000000000000000000000000000, /* 3367 */
128'h00000000000000000000000000000000, /* 3368 */
128'h00000000000000000000000000000000, /* 3369 */
128'h00000000000000000000000000000000, /* 3370 */
128'h00000000000000000000000000000000, /* 3371 */
128'h00000000000000000000000000000000, /* 3372 */
128'h00000000000000000000000000000000, /* 3373 */
128'h00000000000000000000000000000000, /* 3374 */
128'h00000000000000000000000000000000, /* 3375 */
128'h00000000000000000000000000000000, /* 3376 */
128'h00000000000000000000000000000000, /* 3377 */
128'h00000000000000000000000000000000, /* 3378 */
128'h00000000000000000000000000000000, /* 3379 */
128'h00000000000000000000000000000000, /* 3380 */
128'h00000000000000000000000000000000, /* 3381 */
128'h00000000000000000000000000000000, /* 3382 */
128'h00000000000000000000000000000000, /* 3383 */
128'h00000000000000000000000000000000, /* 3384 */
128'h00000000000000000000000000000000, /* 3385 */
128'h00000000000000000000000000000000, /* 3386 */
128'h00000000000000000000000000000000, /* 3387 */
128'h00000000000000000000000000000000, /* 3388 */
128'h00000000000000000000000000000000, /* 3389 */
128'h00000000000000000000000000000000, /* 3390 */
128'h00000000000000000000000000000000, /* 3391 */
128'h00000000000000000000000000000000, /* 3392 */
128'h00000000000000000000000000000000, /* 3393 */
128'h00000000000000000000000000000000, /* 3394 */
128'h00000000000000000000000000000000, /* 3395 */
128'h00000000000000000000000000000000, /* 3396 */
128'h00000000000000000000000000000000, /* 3397 */
128'h00000000000000000000000000000000, /* 3398 */
128'h00000000000000000000000000000000, /* 3399 */
128'h00000000000000000000000000000000, /* 3400 */
128'h00000000000000000000000000000000, /* 3401 */
128'h00000000000000000000000000000000, /* 3402 */
128'h00000000000000000000000000000000, /* 3403 */
128'h00000000000000000000000000000000, /* 3404 */
128'h00000000000000000000000000000000, /* 3405 */
128'h00000000000000000000000000000000, /* 3406 */
128'h00000000000000000000000000000000, /* 3407 */
128'h00000000000000000000000000000000, /* 3408 */
128'h00000000000000000000000000000000, /* 3409 */
128'h00000000000000000000000000000000, /* 3410 */
128'h00000000000000000000000000000000, /* 3411 */
128'h00000000000000000000000000000000, /* 3412 */
128'h00000000000000000000000000000000, /* 3413 */
128'h00000000000000000000000000000000, /* 3414 */
128'h00000000000000000000000000000000, /* 3415 */
128'h00000000000000000000000000000000, /* 3416 */
128'h00000000000000000000000000000000, /* 3417 */
128'h00000000000000000000000000000000, /* 3418 */
128'h00000000000000000000000000000000, /* 3419 */
128'h00000000000000000000000000000000, /* 3420 */
128'h00000000000000000000000000000000, /* 3421 */
128'h00000000000000000000000000000000, /* 3422 */
128'h00000000000000000000000000000000, /* 3423 */
128'h00000000000000000000000000000000, /* 3424 */
128'h00000000000000000000000000000000, /* 3425 */
128'h00000000000000000000000000000000, /* 3426 */
128'h00000000000000000000000000000000, /* 3427 */
128'h00000000000000000000000000000000, /* 3428 */
128'h00000000000000000000000000000000, /* 3429 */
128'h00000000000000000000000000000000, /* 3430 */
128'h00000000000000000000000000000000, /* 3431 */
128'h00000000000000000000000000000000, /* 3432 */
128'h00000000000000000000000000000000, /* 3433 */
128'h00000000000000000000000000000000, /* 3434 */
128'h00000000000000000000000000000000, /* 3435 */
128'h00000000000000000000000000000000, /* 3436 */
128'h00000000000000000000000000000000, /* 3437 */
128'h00000000000000000000000000000000, /* 3438 */
128'h00000000000000000000000000000000, /* 3439 */
128'h00000000000000000000000000000000, /* 3440 */
128'h00000000000000000000000000000000, /* 3441 */
128'h00000000000000000000000000000000, /* 3442 */
128'h00000000000000000000000000000000, /* 3443 */
128'h00000000000000000000000000000000, /* 3444 */
128'h00000000000000000000000000000000, /* 3445 */
128'h00000000000000000000000000000000, /* 3446 */
128'h00000000000000000000000000000000, /* 3447 */
128'h00000000000000000000000000000000, /* 3448 */
128'h00000000000000000000000000000000, /* 3449 */
128'h00000000000000000000000000000000, /* 3450 */
128'h00000000000000000000000000000000, /* 3451 */
128'h00000000000000000000000000000000, /* 3452 */
128'h00000000000000000000000000000000, /* 3453 */
128'h00000000000000000000000000000000, /* 3454 */
128'h00000000000000000000000000000000, /* 3455 */
128'h00000000000000000000000000000000, /* 3456 */
128'h00000000000000000000000000000000, /* 3457 */
128'h00000000000000000000000000000000, /* 3458 */
128'h00000000000000000000000000000000, /* 3459 */
128'h00000000000000000000000000000000, /* 3460 */
128'h00000000000000000000000000000000, /* 3461 */
128'h00000000000000000000000000000000, /* 3462 */
128'h00000000000000000000000000000000, /* 3463 */
128'h00000000000000000000000000000000, /* 3464 */
128'h00000000000000000000000000000000, /* 3465 */
128'h00000000000000000000000000000000, /* 3466 */
128'h00000000000000000000000000000000, /* 3467 */
128'h00000000000000000000000000000000, /* 3468 */
128'h00000000000000000000000000000000, /* 3469 */
128'h00000000000000000000000000000000, /* 3470 */
128'h00000000000000000000000000000000, /* 3471 */
128'h00000000000000000000000000000000, /* 3472 */
128'h00000000000000000000000000000000, /* 3473 */
128'h00000000000000000000000000000000, /* 3474 */
128'h00000000000000000000000000000000, /* 3475 */
128'h00000000000000000000000000000000, /* 3476 */
128'h00000000000000000000000000000000, /* 3477 */
128'h00000000000000000000000000000000, /* 3478 */
128'h00000000000000000000000000000000, /* 3479 */
128'h00000000000000000000000000000000, /* 3480 */
128'h00000000000000000000000000000000, /* 3481 */
128'h00000000000000000000000000000000, /* 3482 */
128'h00000000000000000000000000000000, /* 3483 */
128'h00000000000000000000000000000000, /* 3484 */
128'h00000000000000000000000000000000, /* 3485 */
128'h00000000000000000000000000000000, /* 3486 */
128'h00000000000000000000000000000000, /* 3487 */
128'h00000000000000000000000000000000, /* 3488 */
128'h00000000000000000000000000000000, /* 3489 */
128'h00000000000000000000000000000000, /* 3490 */
128'h00000000000000000000000000000000, /* 3491 */
128'h00000000000000000000000000000000, /* 3492 */
128'h00000000000000000000000000000000, /* 3493 */
128'h00000000000000000000000000000000, /* 3494 */
128'h00000000000000000000000000000000, /* 3495 */
128'h00000000000000000000000000000000, /* 3496 */
128'h00000000000000000000000000000000, /* 3497 */
128'h00000000000000000000000000000000, /* 3498 */
128'h00000000000000000000000000000000, /* 3499 */
128'h00000000000000000000000000000000, /* 3500 */
128'h00000000000000000000000000000000, /* 3501 */
128'h00000000000000000000000000000000, /* 3502 */
128'h00000000000000000000000000000000, /* 3503 */
128'h00000000000000000000000000000000, /* 3504 */
128'h00000000000000000000000000000000, /* 3505 */
128'h00000000000000000000000000000000, /* 3506 */
128'h00000000000000000000000000000000, /* 3507 */
128'h00000000000000000000000000000000, /* 3508 */
128'h00000000000000000000000000000000, /* 3509 */
128'h00000000000000000000000000000000, /* 3510 */
128'h00000000000000000000000000000000, /* 3511 */
128'h00000000000000000000000000000000, /* 3512 */
128'h00000000000000000000000000000000, /* 3513 */
128'h00000000000000000000000000000000, /* 3514 */
128'h00000000000000000000000000000000, /* 3515 */
128'h00000000000000000000000000000000, /* 3516 */
128'h00000000000000000000000000000000, /* 3517 */
128'h00000000000000000000000000000000, /* 3518 */
128'h00000000000000000000000000000000, /* 3519 */
128'h00000000000000000000000000000000, /* 3520 */
128'h00000000000000000000000000000000, /* 3521 */
128'h00000000000000000000000000000000, /* 3522 */
128'h00000000000000000000000000000000, /* 3523 */
128'h00000000000000000000000000000000, /* 3524 */
128'h00000000000000000000000000000000, /* 3525 */
128'h00000000000000000000000000000000, /* 3526 */
128'h00000000000000000000000000000000, /* 3527 */
128'h00000000000000000000000000000000, /* 3528 */
128'h00000000000000000000000000000000, /* 3529 */
128'h00000000000000000000000000000000, /* 3530 */
128'h00000000000000000000000000000000, /* 3531 */
128'h00000000000000000000000000000000, /* 3532 */
128'h00000000000000000000000000000000, /* 3533 */
128'h00000000000000000000000000000000, /* 3534 */
128'h00000000000000000000000000000000, /* 3535 */
128'h00000000000000000000000000000000, /* 3536 */
128'h00000000000000000000000000000000, /* 3537 */
128'h00000000000000000000000000000000, /* 3538 */
128'h00000000000000000000000000000000, /* 3539 */
128'h00000000000000000000000000000000, /* 3540 */
128'h00000000000000000000000000000000, /* 3541 */
128'h00000000000000000000000000000000, /* 3542 */
128'h00000000000000000000000000000000, /* 3543 */
128'h00000000000000000000000000000000, /* 3544 */
128'h00000000000000000000000000000000, /* 3545 */
128'h00000000000000000000000000000000, /* 3546 */
128'h00000000000000000000000000000000, /* 3547 */
128'h00000000000000000000000000000000, /* 3548 */
128'h00000000000000000000000000000000, /* 3549 */
128'h00000000000000000000000000000000, /* 3550 */
128'h00000000000000000000000000000000, /* 3551 */
128'h00000000000000000000000000000000, /* 3552 */
128'h00000000000000000000000000000000, /* 3553 */
128'h00000000000000000000000000000000, /* 3554 */
128'h00000000000000000000000000000000, /* 3555 */
128'h00000000000000000000000000000000, /* 3556 */
128'h00000000000000000000000000000000, /* 3557 */
128'h00000000000000000000000000000000, /* 3558 */
128'h00000000000000000000000000000000, /* 3559 */
128'h00000000000000000000000000000000, /* 3560 */
128'h00000000000000000000000000000000, /* 3561 */
128'h00000000000000000000000000000000, /* 3562 */
128'h00000000000000000000000000000000, /* 3563 */
128'h00000000000000000000000000000000, /* 3564 */
128'h00000000000000000000000000000000, /* 3565 */
128'h00000000000000000000000000000000, /* 3566 */
128'h00000000000000000000000000000000, /* 3567 */
128'h00000000000000000000000000000000, /* 3568 */
128'h00000000000000000000000000000000, /* 3569 */
128'h00000000000000000000000000000000, /* 3570 */
128'h00000000000000000000000000000000, /* 3571 */
128'h00000000000000000000000000000000, /* 3572 */
128'h00000000000000000000000000000000, /* 3573 */
128'h00000000000000000000000000000000, /* 3574 */
128'h00000000000000000000000000000000, /* 3575 */
128'h00000000000000000000000000000000, /* 3576 */
128'h00000000000000000000000000000000, /* 3577 */
128'h00000000000000000000000000000000, /* 3578 */
128'h00000000000000000000000000000000, /* 3579 */
128'h00000000000000000000000000000000, /* 3580 */
128'h00000000000000000000000000000000, /* 3581 */
128'h00000000000000000000000000000000, /* 3582 */
128'h00000000000000000000000000000000, /* 3583 */
128'h00000000000000000000000000000000, /* 3584 */
128'h00000000000000000000000000000000, /* 3585 */
128'h00000000000000000000000000000000, /* 3586 */
128'h00000000000000000000000000000000, /* 3587 */
128'h00000000000000000000000000000000, /* 3588 */
128'h00000000000000000000000000000000, /* 3589 */
128'h00000000000000000000000000000000, /* 3590 */
128'h00000000000000000000000000000000, /* 3591 */
128'h00000000000000000000000000000000, /* 3592 */
128'h00000000000000000000000000000000, /* 3593 */
128'h00000000000000000000000000000000, /* 3594 */
128'h00000000000000000000000000000000, /* 3595 */
128'h00000000000000000000000000000000, /* 3596 */
128'h00000000000000000000000000000000, /* 3597 */
128'h00000000000000000000000000000000, /* 3598 */
128'h00000000000000000000000000000000, /* 3599 */
128'h00000000000000000000000000000000, /* 3600 */
128'h00000000000000000000000000000000, /* 3601 */
128'h00000000000000000000000000000000, /* 3602 */
128'h00000000000000000000000000000000, /* 3603 */
128'h00000000000000000000000000000000, /* 3604 */
128'h00000000000000000000000000000000, /* 3605 */
128'h00000000000000000000000000000000, /* 3606 */
128'h00000000000000000000000000000000, /* 3607 */
128'h00000000000000000000000000000000, /* 3608 */
128'h00000000000000000000000000000000, /* 3609 */
128'h00000000000000000000000000000000, /* 3610 */
128'h00000000000000000000000000000000, /* 3611 */
128'h00000000000000000000000000000000, /* 3612 */
128'h00000000000000000000000000000000, /* 3613 */
128'h00000000000000000000000000000000, /* 3614 */
128'h00000000000000000000000000000000, /* 3615 */
128'h00000000000000000000000000000000, /* 3616 */
128'h00000000000000000000000000000000, /* 3617 */
128'h00000000000000000000000000000000, /* 3618 */
128'h00000000000000000000000000000000, /* 3619 */
128'h00000000000000000000000000000000, /* 3620 */
128'h00000000000000000000000000000000, /* 3621 */
128'h00000000000000000000000000000000, /* 3622 */
128'h00000000000000000000000000000000, /* 3623 */
128'h00000000000000000000000000000000, /* 3624 */
128'h00000000000000000000000000000000, /* 3625 */
128'h00000000000000000000000000000000, /* 3626 */
128'h00000000000000000000000000000000, /* 3627 */
128'h00000000000000000000000000000000, /* 3628 */
128'h00000000000000000000000000000000, /* 3629 */
128'h00000000000000000000000000000000, /* 3630 */
128'h00000000000000000000000000000000, /* 3631 */
128'h00000000000000000000000000000000, /* 3632 */
128'h00000000000000000000000000000000, /* 3633 */
128'h00000000000000000000000000000000, /* 3634 */
128'h00000000000000000000000000000000, /* 3635 */
128'h00000000000000000000000000000000, /* 3636 */
128'h00000000000000000000000000000000, /* 3637 */
128'h00000000000000000000000000000000, /* 3638 */
128'h00000000000000000000000000000000, /* 3639 */
128'h00000000000000000000000000000000, /* 3640 */
128'h00000000000000000000000000000000, /* 3641 */
128'h00000000000000000000000000000000, /* 3642 */
128'h00000000000000000000000000000000, /* 3643 */
128'h00000000000000000000000000000000, /* 3644 */
128'h00000000000000000000000000000000, /* 3645 */
128'h00000000000000000000000000000000, /* 3646 */
128'h00000000000000000000000000000000, /* 3647 */
128'h00000000000000000000000000000000, /* 3648 */
128'h00000000000000000000000000000000, /* 3649 */
128'h00000000000000000000000000000000, /* 3650 */
128'h00000000000000000000000000000000, /* 3651 */
128'h00000000000000000000000000000000, /* 3652 */
128'h00000000000000000000000000000000, /* 3653 */
128'h00000000000000000000000000000000, /* 3654 */
128'h00000000000000000000000000000000, /* 3655 */
128'h00000000000000000000000000000000, /* 3656 */
128'h00000000000000000000000000000000, /* 3657 */
128'h00000000000000000000000000000000, /* 3658 */
128'h00000000000000000000000000000000, /* 3659 */
128'h00000000000000000000000000000000, /* 3660 */
128'h00000000000000000000000000000000, /* 3661 */
128'h00000000000000000000000000000000, /* 3662 */
128'h00000000000000000000000000000000, /* 3663 */
128'h00000000000000000000000000000000, /* 3664 */
128'h00000000000000000000000000000000, /* 3665 */
128'h00000000000000000000000000000000, /* 3666 */
128'h00000000000000000000000000000000, /* 3667 */
128'h00000000000000000000000000000000, /* 3668 */
128'h00000000000000000000000000000000, /* 3669 */
128'h00000000000000000000000000000000, /* 3670 */
128'h00000000000000000000000000000000, /* 3671 */
128'h00000000000000000000000000000000, /* 3672 */
128'h00000000000000000000000000000000, /* 3673 */
128'h00000000000000000000000000000000, /* 3674 */
128'h00000000000000000000000000000000, /* 3675 */
128'h00000000000000000000000000000000, /* 3676 */
128'h00000000000000000000000000000000, /* 3677 */
128'h00000000000000000000000000000000, /* 3678 */
128'h00000000000000000000000000000000, /* 3679 */
128'h00000000000000000000000000000000, /* 3680 */
128'h00000000000000000000000000000000, /* 3681 */
128'h00000000000000000000000000000000, /* 3682 */
128'h00000000000000000000000000000000, /* 3683 */
128'h00000000000000000000000000000000, /* 3684 */
128'h00000000000000000000000000000000, /* 3685 */
128'h00000000000000000000000000000000, /* 3686 */
128'h00000000000000000000000000000000, /* 3687 */
128'h00000000000000000000000000000000, /* 3688 */
128'h00000000000000000000000000000000, /* 3689 */
128'h00000000000000000000000000000000, /* 3690 */
128'h00000000000000000000000000000000, /* 3691 */
128'h00000000000000000000000000000000, /* 3692 */
128'h00000000000000000000000000000000, /* 3693 */
128'h00000000000000000000000000000000, /* 3694 */
128'h00000000000000000000000000000000, /* 3695 */
128'h00000000000000000000000000000000, /* 3696 */
128'h00000000000000000000000000000000, /* 3697 */
128'h00000000000000000000000000000000, /* 3698 */
128'h00000000000000000000000000000000, /* 3699 */
128'h00000000000000000000000000000000, /* 3700 */
128'h00000000000000000000000000000000, /* 3701 */
128'h00000000000000000000000000000000, /* 3702 */
128'h00000000000000000000000000000000, /* 3703 */
128'h00000000000000000000000000000000, /* 3704 */
128'h00000000000000000000000000000000, /* 3705 */
128'h00000000000000000000000000000000, /* 3706 */
128'h00000000000000000000000000000000, /* 3707 */
128'h00000000000000000000000000000000, /* 3708 */
128'h00000000000000000000000000000000, /* 3709 */
128'h00000000000000000000000000000000, /* 3710 */
128'h00000000000000000000000000000000, /* 3711 */
128'h00000000000000000000000000000000, /* 3712 */
128'h00000000000000000000000000000000, /* 3713 */
128'h00000000000000000000000000000000, /* 3714 */
128'h00000000000000000000000000000000, /* 3715 */
128'h00000000000000000000000000000000, /* 3716 */
128'h00000000000000000000000000000000, /* 3717 */
128'h00000000000000000000000000000000, /* 3718 */
128'h00000000000000000000000000000000, /* 3719 */
128'h00000000000000000000000000000000, /* 3720 */
128'h00000000000000000000000000000000, /* 3721 */
128'h00000000000000000000000000000000, /* 3722 */
128'h00000000000000000000000000000000, /* 3723 */
128'h00000000000000000000000000000000, /* 3724 */
128'h00000000000000000000000000000000, /* 3725 */
128'h00000000000000000000000000000000, /* 3726 */
128'h00000000000000000000000000000000, /* 3727 */
128'h00000000000000000000000000000000, /* 3728 */
128'h00000000000000000000000000000000, /* 3729 */
128'h00000000000000000000000000000000, /* 3730 */
128'h00000000000000000000000000000000, /* 3731 */
128'h00000000000000000000000000000000, /* 3732 */
128'h00000000000000000000000000000000, /* 3733 */
128'h00000000000000000000000000000000, /* 3734 */
128'h00000000000000000000000000000000, /* 3735 */
128'h00000000000000000000000000000000, /* 3736 */
128'h00000000000000000000000000000000, /* 3737 */
128'h00000000000000000000000000000000, /* 3738 */
128'h00000000000000000000000000000000, /* 3739 */
128'h00000000000000000000000000000000, /* 3740 */
128'h00000000000000000000000000000000, /* 3741 */
128'h00000000000000000000000000000000, /* 3742 */
128'h00000000000000000000000000000000, /* 3743 */
128'h00000000000000000000000000000000, /* 3744 */
128'h00000000000000000000000000000000, /* 3745 */
128'h00000000000000000000000000000000, /* 3746 */
128'h00000000000000000000000000000000, /* 3747 */
128'h00000000000000000000000000000000, /* 3748 */
128'h00000000000000000000000000000000, /* 3749 */
128'h00000000000000000000000000000000, /* 3750 */
128'h00000000000000000000000000000000, /* 3751 */
128'h00000000000000000000000000000000, /* 3752 */
128'h00000000000000000000000000000000, /* 3753 */
128'h00000000000000000000000000000000, /* 3754 */
128'h00000000000000000000000000000000, /* 3755 */
128'h00000000000000000000000000000000, /* 3756 */
128'h00000000000000000000000000000000, /* 3757 */
128'h00000000000000000000000000000000, /* 3758 */
128'h00000000000000000000000000000000, /* 3759 */
128'h00000000000000000000000000000000, /* 3760 */
128'h00000000000000000000000000000000, /* 3761 */
128'h00000000000000000000000000000000, /* 3762 */
128'h00000000000000000000000000000000, /* 3763 */
128'h00000000000000000000000000000000, /* 3764 */
128'h00000000000000000000000000000000, /* 3765 */
128'h00000000000000000000000000000000, /* 3766 */
128'h00000000000000000000000000000000, /* 3767 */
128'h00000000000000000000000000000000, /* 3768 */
128'h00000000000000000000000000000000, /* 3769 */
128'h00000000000000000000000000000000, /* 3770 */
128'h00000000000000000000000000000000, /* 3771 */
128'h00000000000000000000000000000000, /* 3772 */
128'h00000000000000000000000000000000, /* 3773 */
128'h00000000000000000000000000000000, /* 3774 */
128'h00000000000000000000000000000000, /* 3775 */
128'h00000000000000000000000000000000, /* 3776 */
128'h00000000000000000000000000000000, /* 3777 */
128'h00000000000000000000000000000000, /* 3778 */
128'h00000000000000000000000000000000, /* 3779 */
128'h00000000000000000000000000000000, /* 3780 */
128'h00000000000000000000000000000000, /* 3781 */
128'h00000000000000000000000000000000, /* 3782 */
128'h00000000000000000000000000000000, /* 3783 */
128'h00000000000000000000000000000000, /* 3784 */
128'h00000000000000000000000000000000, /* 3785 */
128'h00000000000000000000000000000000, /* 3786 */
128'h00000000000000000000000000000000, /* 3787 */
128'h00000000000000000000000000000000, /* 3788 */
128'h00000000000000000000000000000000, /* 3789 */
128'h00000000000000000000000000000000, /* 3790 */
128'h00000000000000000000000000000000, /* 3791 */
128'h00000000000000000000000000000000, /* 3792 */
128'h00000000000000000000000000000000, /* 3793 */
128'h00000000000000000000000000000000, /* 3794 */
128'h00000000000000000000000000000000, /* 3795 */
128'h00000000000000000000000000000000, /* 3796 */
128'h00000000000000000000000000000000, /* 3797 */
128'h00000000000000000000000000000000, /* 3798 */
128'h00000000000000000000000000000000, /* 3799 */
128'h00000000000000000000000000000000, /* 3800 */
128'h00000000000000000000000000000000, /* 3801 */
128'h00000000000000000000000000000000, /* 3802 */
128'h00000000000000000000000000000000, /* 3803 */
128'h00000000000000000000000000000000, /* 3804 */
128'h00000000000000000000000000000000, /* 3805 */
128'h00000000000000000000000000000000, /* 3806 */
128'h00000000000000000000000000000000, /* 3807 */
128'h00000000000000000000000000000000, /* 3808 */
128'h00000000000000000000000000000000, /* 3809 */
128'h00000000000000000000000000000000, /* 3810 */
128'h00000000000000000000000000000000, /* 3811 */
128'h00000000000000000000000000000000, /* 3812 */
128'h00000000000000000000000000000000, /* 3813 */
128'h00000000000000000000000000000000, /* 3814 */
128'h00000000000000000000000000000000, /* 3815 */
128'h00000000000000000000000000000000, /* 3816 */
128'h00000000000000000000000000000000, /* 3817 */
128'h00000000000000000000000000000000, /* 3818 */
128'h00000000000000000000000000000000, /* 3819 */
128'h00000000000000000000000000000000, /* 3820 */
128'h00000000000000000000000000000000, /* 3821 */
128'h00000000000000000000000000000000, /* 3822 */
128'h00000000000000000000000000000000, /* 3823 */
128'h00000000000000000000000000000000, /* 3824 */
128'h00000000000000000000000000000000, /* 3825 */
128'h00000000000000000000000000000000, /* 3826 */
128'h00000000000000000000000000000000, /* 3827 */
128'h00000000000000000000000000000000, /* 3828 */
128'h00000000000000000000000000000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00000000000000000000000000000000, /* 3840 */
128'h00000000000000000000000000000000, /* 3841 */
128'h00000000000000000000000000000000, /* 3842 */
128'h00000000000000000000000000000000, /* 3843 */
128'h00000000000000000000000000000000, /* 3844 */
128'h00000000000000000000000000000000, /* 3845 */
128'h00000000000000000000000000000000, /* 3846 */
128'h00000000000000000000000000000000, /* 3847 */
128'h00000000000000000000000000000000, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule

