/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 1195;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h0a646c25_2e646c25,
        64'h203d2049_5043202c,
        64'h73656c63_79632064,
        64'h6c25202c_736e6f69,
        64'h74637572_74736e69,
        64'h20646c25_202c424b,
        64'h6425203d_20746573,
        64'h5f676e69_6b726f77,
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h00000000_0000000a,
        64'h0d6b636f_6c622044,
        64'h53206461_65722074,
        64'h6f6e2064_6c756f63,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00322d74_6c756166,
        64'h65642d69_72742c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_6972742c,
        64'h786e6c78_006c6175,
        64'h642d7369_2c786e6c,
        64'h7800746e_65736572,
        64'h702d7470_75727265,
        64'h746e692c_786e6c78,
        64'h00687464_69772d32,
        64'h6f697067_2c786e6c,
        64'h78006874_6469772d,
        64'h6f697067_2c786e6c,
        64'h7800322d_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800746c,
        64'h75616665_642d7475,
        64'h6f642c78_6e6c7800,
        64'h322d7374_75706e69,
        64'h2d6c6c61_2c786e6c,
        64'h78007374_75706e69,
        64'h2d6c6c61_2c786e6c,
        64'h78007265_6c6c6f72,
        64'h746e6f63_2d6f6970,
        64'h6700736c_6c65632d,
        64'h6f697067_23007373,
        64'h65726464_612d6361,
        64'h6d2d6c61_636f6c00,
        64'h70772d65_6c626173,
        64'h69640073_65676e61,
        64'h722d6567_61746c6f,
        64'h76007963_6e657571,
        64'h6572662d_78616d2d,
        64'h69707300_6f697461,
        64'h722d6b63_732c786e,
        64'h6c780073_7469622d,
        64'h72656673_6e617274,
        64'h2d6d756e_2c786e6c,
        64'h78007374_69622d73,
        64'h732d6d75_6e2c786e,
        64'h6c780074_73697865,
        64'h2d6f6669_662c786e,
        64'h6c780079_6c696d61,
        64'h662c786e_6c780068,
        64'h74646977_2d6f692d,
        64'h67657200_74666968,
        64'h732d6765_72007374,
        64'h70757272_65746e69,
        64'h00746e65_7261702d,
        64'h74707572_7265746e,
        64'h69006465_6570732d,
        64'h746e6572_72756300,
        64'h7665646e_2c766373,
        64'h69720079_7469726f,
        64'h6972702d_78616d2c,
        64'h76637369_72007365,
        64'h6d616e2d_67657200,
        64'h6465646e_65747865,
        64'h2d737470_75727265,
        64'h746e6900_7365676e,
        64'h61720064_65646e65,
        64'h70737573_2d657461,
        64'h74732d6e_69617465,
        64'h72007265_67676972,
        64'h742d746c_75616665,
        64'h642c7875_6e696c00,
        64'h736f6970_6700656c,
        64'h646e6168_702c7875,
        64'h6e696c00_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_bb000000,
        64'h04000000_03000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_c5020000,
        64'h04000000_03000000,
        64'hffffffff_b4020000,
        64'h04000000_03000000,
        64'h01000000_a7020000,
        64'h04000000_03000000,
        64'h00000000_90020000,
        64'h04000000_03000000,
        64'h08000000_7f020000,
        64'h04000000_03000000,
        64'h08000000_6f020000,
        64'h04000000_03000000,
        64'h00000000_5b020000,
        64'h04000000_03000000,
        64'h00000000_49020000,
        64'h04000000_03000000,
        64'h00000000_37020000,
        64'h04000000_03000000,
        64'h00000000_27020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_17020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h0b020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf9010000_06000000,
        64'h03000000_00000000,
        64'h03000000_58010000,
        64'h08000000_03000000,
        64'h03000000_47010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'hee010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_df010000,
        64'h08000000_03000000,
        64'h20bcbe00_cd010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_be010000,
        64'h04000000_03000000,
        64'h08000000_a7010000,
        64'h04000000_03000000,
        64'h01000000_96010000,
        64'h04000000_03000000,
        64'h01000000_86010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h7a010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h58010000_08000000,
        64'h03000000_03000000,
        64'h47010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_04000000,
        64'h6d010000_04000000,
        64'h03000000_02000000,
        64'h63010000_04000000,
        64'h03000000_01000000,
        64'h58010000_04000000,
        64'h03000000_03000000,
        64'h47010000_04000000,
        64'h03000000_00c20100,
        64'h39010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_11010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_fd000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_bb000000,
        64'h04000000_03000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_2e010000,
        64'h04000000_03000000,
        64'h07000000_1b010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_fd000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_11010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_fd000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf6000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hdf000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc9000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hc3000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_bb000000,
        64'h04000000_03000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00007573_63616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00090000_d8020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h38090000_38000000,
        64'h100c0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha0018402_2ec58593,
        64'h00000597_01f41413,
        64'h0010041b_e911cacf,
        64'hf0ef057e_65a14505,
        64'hfecff0ef_e6bfe0ef,
        64'hf2050513_00001517,
        64'he45fe0ef_e4061141,
        64'hb7f1377d_87aabfa5,
        64'hfef51be3_0785f8b7,
        64'h12e30007_c70300d8,
        64'h0a630087_85130007,
        64'hb803bfcd_367d0785,
        64'hf8b71fe3_0007c703,
        64'hd24d8a1d_eb1187aa,
        64'h27018edd_00365713,
        64'h02079693_8fd90107,
        64'h179300b7_e7330085,
        64'h97938e1d_953e9381,
        64'h02071793_faf50785,
        64'h36fdfcb8_1ce30007,
        64'hc80387aa_0007069b,
        64'h40e7873b_47a1c31d,
        64'h00757713_b7f5367d,
        64'h0785feb7_1ce30007,
        64'hc7038082_853e4781,
        64'he60187aa_260100c7,
        64'hef630ff5_f59347c1,
        64'hb7ed853e_feb70be3,
        64'h00150793_00054703,
        64'h80824501_00c51463,
        64'h0ff5f593_962abfe9,
        64'h0405d175_f8bff0ef,
        64'h397d8522_85ce8626,
        64'h80826145_69a26942,
        64'h64e27402_70a28522,
        64'h44010099_5b630005,
        64'h091bd15f_f0ef8522,
        64'hc8890005_049bd21f,
        64'hf0ef89ae_e84af406,
        64'he44eec26_852e842a,
        64'hf0227179_bfc50505,
        64'hfeb78de3_00054783,
        64'h808200c5_1363962a,
        64'hb7dd0585_0505fbed,
        64'h9f990005_c7030005,
        64'h47838082_853e4781,
        64'h00c51563_962ab7fd,
        64'h00f68023_16fd0005,
        64'hc78315fd_d7e500e5,
        64'h87b340b6_073300c5,
        64'h06b395b2_80820141,
        64'h640260a2_8522f57f,
        64'hf0ef00a5_e963842a,
        64'he406e022_11418082,
        64'h614564e2_69428526,
        64'h740270a2_00040023,
        64'hf79ff0ef_944a864a,
        64'h8522fff6_091300c5,
        64'h64636582_892ace11,
        64'h84aa6622_dcfff0ef,
        64'he02ee84a_f406e432,
        64'hec26852e_842af022,
        64'h7179bf65_fee78fa3,
        64'h0785fff5_c7030585,
        64'hbfe1469d_00c508b3,
        64'h87aa872e_bfc100e5,
        64'h07b3963e_95ba070e,
        64'h02f707b3_57e10036,
        64'h5713ff06_e8e340f8,
        64'h8833ff07_bc2307a1,
        64'hff873803_07218082,
        64'h02c79e63_963e87aa,
        64'hcb9d8b9d_00a5e7b3,
        64'h00b50a63_bf6dfeb7,
        64'h8fa30785_bfe1fef7,
        64'h3c230721_bfd10ff5,
        64'hf6934725_bfc1963a,
        64'h97aa078e_02e78733,
        64'h57610036_57930106,
        64'hef6340e8_8833469d,
        64'h00c508b3_872aff6d,
        64'h377d8fd5_07a28082,
        64'h04c79063_963e87aa,
        64'hcb9d0075_77938082,
        64'h4501b7e5_078900d7,
        64'h80a300e7_80238082,
        64'he3110017_c703ce81,
        64'h0007c683_87aacf99,
        64'h00054783_c11d8082,
        64'h610564a2_85266442,
        64'h60e2e008_05050005,
        64'h0023c501_f75ff0ef,
        64'h8526842a_c891e822,
        64'hec066104_e4261101,
        64'hbfd94ca7_bd230000,
        64'h07970505_00050023,
        64'hc7810005_4783c519,
        64'hfa1ff0ef_852285a6,
        64'h80826105_64a26442,
        64'h60e28522_44015007,
        64'hb3230000_0797ef81,
        64'h00044783_942af9ff,
        64'hf0ef85a6_8522cc11,
        64'h5207b403_00000797,
        64'he511842a_84aeec06,
        64'he426e822_1101bfd5,
        64'h87aeb7e5_0505fafd,
        64'h0007c683_0785fee6,
        64'h8fe38082_4501eb19,
        64'h00054703_bff90785,
        64'hbfd5872e_8082fe08,
        64'h1be30007_48030705,
        64'h00c80a63_8082ea11,
        64'h40d78533_0007c603,
        64'h87aa86aa_bfcd872e,
        64'hb7d50785_fe081be3,
        64'h00074803_0705fed8,
        64'h0fe38082_ea9940c7,
        64'h85330007_c68387aa,
        64'h862ab7fd_07858082,
        64'h40a78533_e7010007,
        64'hc70300b7_856387aa,
        64'h95aa8082_61056442,
        64'h60e24501_fe857be3,
        64'h157d00b7_86630005,
        64'h47830ff5_f5939522,
        64'h65a2fe5f_f0efec06,
        64'h842ae42e_e8221101,
        64'hbfcd0785_808240a7,
        64'h8533e701_0007c703,
        64'h87aabfcd_0505dffd,
        64'h808200b7_93630005,
        64'h47830ff5_f5938082,
        64'h4501bfcd_0505c399,
        64'h808200b7_93630005,
        64'h47830ff5_f5938082,
        64'h853eff79_0505e399,
        64'h4187d79b_0187979b,
        64'h40f707bb_fff5c783,
        64'h00054703_0585a839,
        64'h478100c5_9463962e,
        64'h8082853e_f37d0505,
        64'he3994187_d79b0187,
        64'h979b40f7_07bbfff5,
        64'hc7830005_47030585,
        64'hb7cd87ba_80820007,
        64'h80a300c7_15638082,
        64'he291fed7_0fa30017,
        64'h8713fff5_c6830585,
        64'h963efb7d_00178693,
        64'h0007c703_87b68082,
        64'he21987aa_b7d587b6,
        64'h8082fb75_fee78fa3,
        64'h0785fff5_c7030585,
        64'heb090017_86930007,
        64'hc70387aa_8082fb65,
        64'hfee78fa3_0785fff5,
        64'hc7030585_00c78963,
        64'h87aa962a_8082fb75,
        64'hfee78fa3_0785fff5,
        64'hc7030585_87aa8082,
        64'h61356452_60f28522,
        64'hb56ff0ef_0808842a,
        64'he3fff0ef_e436eec6,
        64'heac2e6be_e2baea22,
        64'hee060808_10000593,
        64'h1234862a_fe36fa32,
        64'hf62e710d_80826161,
        64'h60e2e69f_f0efe436,
        64'he4c6e0c2_fc3ef83a,
        64'hec061000_05931014,
        64'h862ef436_f032715d,
        64'h80826161_60e2e8df,
        64'hf0efe436_e4c6e0c2,
        64'hfc3ef83a_ec061034,
        64'hf436715d_b7f18522,
        64'h02010393_0005059b,
        64'h17a000ef_85220124,
        64'h74336000_00840b13,
        64'hb5fd845a_d93ff0ef,
        64'h00840b13_02010393,
        64'h00044503_a809ddbf,
        64'hf0ef0028_02010393,
        64'h0005059b_e37ff0ef,
        64'h400845a9_46010016,
        64'hb6930038_00840b13,
        64'hf8b50693_a81145c1,
        64'h00163613_46850038,
        64'h00840b13_fa850613,
        64'hf6e510e3_07800713,
        64'h02e50063_07500713,
        64'ha00d4601_46850038,
        64'h00840b13_f6e51ee3,
        64'h07000713_00a76c63,
        64'h06e50e63_07300713,
        64'hb74d048d_0024c503,
        64'h80826109_0007051b,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_744670e6,
        64'hf55d08f5_09630630,
        64'h079304d5_0f630580,
        64'h069302a6_eb6306d5,
        64'h0f630640_06930489,
        64'h0014c503_478100f6,
        64'hf36346a5_0ff7f793,
        64'hfd07879b_cb9d0004,
        64'hc7830355_10634781,
        64'h04890545_0f630014,
        64'hc503bfe1_e7bff0ef,
        64'h02010393_04850135,
        64'h086304d7_ff639381,
        64'h17827682_0017079b,
        64'hc52d8f1d_0004c503,
        64'h77a27742_02095913,
        64'h03000a93_06c00a13,
        64'h02500993_f82af02e,
        64'hf42afc3e_843684b2,
        64'he0dafc86_e4d6e8d2,
        64'heccef4a6_f8a2597d,
        64'h011cf0ca_7119b7f1,
        64'h06850117_80230066,
        64'h80232605_0006c883,
        64'h0007c303_97ba9381,
        64'h178240c8_07bbb7d9,
        64'h2585fea6_8fa30685,
        64'hbf5d00a8_053b8082,
        64'h00b61b63_fff5081b,
        64'h86ba2581_00068023,
        64'h0015559b_40e6853b,
        64'h068500f6_802302d0,
        64'h07930008_876302f5,
        64'he9630300_051340e6,
        64'h85bbfe71_8532fea6,
        64'h8fa30685_0ff57513,
        64'h02b6563b_0305051b,
        64'h046e6763_0ff37513,
        64'h02b6733b_0005061b,
        64'h385986ba_4e250ff6,
        64'hf8130410_0693c219,
        64'h06100693_488540a0,
        64'h053be681_00055663,
        64'h4881bfe9_00d70023,
        64'h07850007_c68300d3,
        64'hb8230017_06938082,
        64'h852e0007_002300b6,
        64'he6630103_b70340a7,
        64'h86bb87aa_9d9dfff7,
        64'h059b00c6_f5638e9d,
        64'hfff70693_0003b703,
        64'h8f999201_02059613,
        64'h0103b783_0083b703,
        64'h80824501_80820007,
        64'h80234505_0103b783,
        64'h00a70023_00f3b823,
        64'h00170793_00d7fe63,
        64'h93811782_278540f7,
        64'h07b30003_b6830083,
        64'hb7830103_b703bff1,
        64'hf5dff0ef_4541f63f,
        64'hf0ef4521_f69ff0ef,
        64'h4511f6ff_f0ef4509,
        64'hf75ff0ef_4505f7bf,
        64'hf0ef4501_e4061141,
        64'hbf51c000_28f3c020,
        64'h26f3fac7_10e330e0,
        64'h006fa425_05130000,
        64'h251702a7_473302a7,
        64'h67b302b3_45bb02c7,
        64'h47334000_059302a6,
        64'h87334116_86b33e80,
        64'h0513c000_26f38e15,
        64'hc0202673_02b71d63,
        64'h2705fe08_13e397aa,
        64'h387d0007_802397aa,
        64'h00078023_97aa0007,
        64'h802397aa_00078023,
        64'h40000813_87f245a9,
        64'h01f61e13_46814881,
        64'h470100c5_131b4605,
        64'hbbb5f00f_f0efaa65,
        64'h05130000_2517b3f5,
        64'h80050513_00002517,
        64'hf98ff0ef_8526f1cf,
        64'hf0ef9025_05130000,
        64'h2517f28f_f0ef8f65,
        64'h05130000_2517c50d,
        64'h84aac33f_f0ef8552,
        64'h865a020a_a583f44f,
        64'hf0efad25_05130000,
        64'h2517f579_93e30804,
        64'h8493f58f_f0ef2985,
        64'h85050513_00002517,
        64'hff2c1be3_82fff0ef,
        64'h09050009_4503f74f,
        64'hf0efaf25_05130000,
        64'h2517803f_f0ef7088,
        64'hf86ff0ef_af450513,
        64'h00002517_815ff0ef,
        64'h6c88f98f_f0efaf65,
        64'h05130000_2517827f,
        64'hf0ef0704_8c130284,
        64'h89136888_fb2ff0ef,
        64'hb0050513_00002517,
        64'hff2c1be3_887ff0ef,
        64'h09050009_45030109,
        64'h0c13fd0f_f0efafe5,
        64'h05130000_2517fe99,
        64'h1be38a5f_f0ef0905,
        64'h00094503_ff048913,
        64'hfeeff0ef_afc50513,
        64'h00002517_8bfff0ef,
        64'h0ff9f513_803ff0ef,
        64'haf850513_00002517,
        64'hb5fd9025_05130000,
        64'h251789bf_f0ef854e,
        64'h81fff0ef_a0450513,
        64'h00002517_82bff0ef,
        64'h9f850513_00002517,
        64'hc50d0804_89aa8a8a,
        64'hd39ff0ef_850a4605,
        64'h71010489_258384df,
        64'hf0ef9425_05130000,
        64'h251789bf_f0ef4556,
        64'h85fff0ef_b3450513,
        64'h00002517_8adff0ef,
        64'h4546871f_f0efb265,
        64'h05130000_25178fff,
        64'hf0ef6526_883ff0ef,
        64'hb1850513_00002517,
        64'h911ff0ef_7502895f,
        64'hf0efb1a5_05130000,
        64'h2517923f_f0ef6562,
        64'h8a7ff0ef_b1450513,
        64'h00002517_8f5ff0ef,
        64'h45528b9f_f0efb165,
        64'h05130000_2517907f,
        64'hf0ef4542_8cbff0ef,
        64'hb1850513_00002517,
        64'h919ff0ef_45328ddf,
        64'hf0efb1a5_05130000,
        64'h251792bf_f0ef4522,
        64'h8efff0ef_b1c50513,
        64'h00002517_97dff0ef,
        64'h4b916502_903ff0ef,
        64'hb2050513_00002517,
        64'h90fff0ef_b0c50513,
        64'h00002517_bf6154f9,
        64'h91fff0ef_a1450513,
        64'h00002517_9adff0ef,
        64'h8526931f_f0efb165,
        64'h05130000_251793df,
        64'hf0efb0a5_05130000,
        64'h2517c905_84aa890a,
        64'he49ff0ef_850a4585,
        64'h46057101_95bff0ef,
        64'hb1050513_00002517,
        64'h80826161_6c026ba2,
        64'h6b426ae2_7a0279a2,
        64'h794274e2_64068526,
        64'h60a6fb04_011354fd,
        64'h987ff0ef_b1450513,
        64'h00002517_c51ddf3f,
        64'hf0ef8b2e_8a2a0880,
        64'he062e45e_ec56f44e,
        64'hf84afc26_e486e85a,
        64'hf052e0a2_715db765,
        64'h54798082_61696baa,
        64'h6b4a6aea_7a0a79aa,
        64'h794a74ea_640e60ae,
        64'h8522547d_9d3ff0ef,
        64'hb3850513_00002517,
        64'hc59ff0ef_c5dff0ef,
        64'hc61ff0ef_c65ff0ef,
        64'hc69ff0ef_c6dff0ef,
        64'hc71ff0ef_c75ff0ef,
        64'ha805c7bf_f0efc87f,
        64'hf0ef4531_45814605,
        64'h4401f930_46e319fd,
        64'ha17ff0ef_b9c50513,
        64'h00002517_e7990359,
        64'he7b30724_1a632901,
        64'h90411442_8c49caff,
        64'hf0ef9041_03051413,
        64'h84a20085_151bcbff,
        64'hf0effd64_1ae30404,
        64'h0413ff74_97e3892a,
        64'hf13ff0ef_0485854a,
        64'h0007c583_009407b3,
        64'h04000b93_4481c67f,
        64'hf0ef850a_04000593,
        64'h86224901_84262004,
        64'h8b13ff45_1ee3cfff,
        64'hf0ef3e80_0a930fe0,
        64'h0a13e951_d15ff0ef,
        64'h454985a2_0ff67613,
        64'h00166613_0015161b,
        64'hf49ff0ef_0ff47593,
        64'hf51ff0ef_0ff5f593,
        64'h0084559b_f5dff0ef,
        64'h0ff5f593_0104559b,
        64'hf69ff0ef_45010ff5,
        64'hf5930184_559bfee7,
        64'h9be30785_00c68023,
        64'h00f106b3_08000713,
        64'h567d4781_0209d993,
        64'h842e84aa_e55ee95a,
        64'hed56f152_f94ae586,
        64'hfd26e1a2_02061993,
        64'hf54e7155_80829141,
        64'h15428d3d_8ff90057,
        64'h979b1701_67090107,
        64'hd79b0105_179b4105,
        64'h551b0105_151b8d2d,
        64'h00c59513_8da9893d,
        64'h0045d51b_8da99141,
        64'h15428d5d_05220085,
        64'h579b8082_07f57513,
        64'h8d2d0045_15938d2d,
        64'h8d3d0045_d51b0075,
        64'hd79b8de9_80820141,
        64'h853e6402_60a24781,
        64'hc11157f5_f89ff0ef,
        64'hc51157f9_efbff0ef,
        64'hc91157fd_eb7ff0ef,
        64'hfc6de03f_f0ef347d,
        64'h4429b91f_f0efcde5,
        64'h05130000_2517c89f,
        64'hf0efe022_e4061141,
        64'h80826105_00153513,
        64'h64a26442_60e20004,
        64'h051bfc94_0ce3e37f,
        64'hf0efeb3f_f0efd065,
        64'h05130000_251785aa,
        64'h842ae53f_f0ef0290,
        64'h05134000_05b70770,
        64'h0613fbdf_f0ef4485,
        64'he822ec06_e4261101,
        64'h80820141_00153513,
        64'h157d6402_60a20004,
        64'h051bef3f_f0efd405,
        64'h051385a2_00002517,
        64'he89ff0ef_842ae97f,
        64'hf0efe022_e4060370,
        64'h05134581_06500613,
        64'h11418082_61056902,
        64'h64a26442_60e20015,
        64'h3513f565_05130004,
        64'h051b0124_986388bd,
        64'h00f91b63_45014785,
        64'hec9ff0ef_ecdff0ef,
        64'h842aed3f_f0ef84aa,
        64'hed9ff0ef_eddff0ef,
        64'hee1ff0ef_892aeeff,
        64'hf0efe04a_e426e822,
        64'hec064521_1aa00593,
        64'h08700613_1101bfcd,
        64'h45018082_61056902,
        64'h64a26442_60e24505,
        64'hf89ff0ef_4585dce5,
        64'h05130000_2517fe99,
        64'h15e3c00d_f25ff0ef,
        64'h892a347d_f35ff0ef,
        64'h45014581_09500613,
        64'h44857104_0413e04a,
        64'hec06e426_6409e822,
        64'h1101cd1f_f06f6105,
        64'hdc850513_00002517,
        64'h60e26442_da7ff0ef,
        64'h852e65a2_cebff0ef,
        64'he1050513_00002517,
        64'hcf7ff0ef_8522cfdf,
        64'hf0efe42e_ec06e165,
        64'h05130000_2517842a,
        64'he8221101_80826145,
        64'h64e27402_70a2f47d,
        64'h147d0007_d4634187,
        64'hd79b0185_179bfa7f,
        64'hf0efeb5f_f0ef8532,
        64'h06400413_6622ec1f,
        64'hf0ef0ff4_7513ec9f,
        64'hf0ef0ff5_75130084,
        64'h551bed5f_f0ef0ff5,
        64'h75130104_551bee1f,
        64'hf0ef0ff5_75130184,
        64'h551beedf_f0ef0404,
        64'he513febf_f0ef84aa,
        64'h842eec26_f022e432,
        64'hf4067179_f07ff06f,
        64'h0ff00513_8082557d,
        64'hb7e900d7_00230785,
        64'h00f60733_06c82683,
        64'hff798b05_5178bf4d,
        64'hd6b80785_0007c703,
        64'h80824501_d3b84719,
        64'hdbb8577d_200007b7,
        64'h00b6ef63_0007869b,
        64'h20000837_20000537,
        64'hfff58b85_537c2000,
        64'h0737d3b8_200007b7,
        64'h10600713_fff537fd,
        64'h00010320_079304b7,
        64'h616340a7_873b87aa,
        64'h200006b7_dbb85779,
        64'h200007b7_06b7ec63,
        64'h10000793_80826105,
        64'h64a2d3b8_4719dbb8,
        64'h644260e2_0ff47513,
        64'h577d2000_07b7e25f,
        64'hf0eff1a5_05130000,
        64'h2517eb3f_f0ef9101,
        64'h15024088_e3bff0ef,
        64'hf3850513_00002517,
        64'he3958b85_240153fc,
        64'h57e0ff65_8b050647,
        64'h849353f8_d3b81060,
        64'h07132000_07b7fff5,
        64'h37fd0001_06400793,
        64'hd7a8dbb8_5779e426,
        64'he822ec06_200007b7,
        64'h1101e81f_f06f6105,
        64'hf6850513_00002517,
        64'h64a260e2_6442d03c,
        64'h4799e99f_f0eff8e5,
        64'h05130000_2517f27f,
        64'hf0ef9101_02049513,
        64'h2481eb1f_f0eff865,
        64'h05130000_25175064,
        64'hd03c1660_0793ec5f,
        64'hf0effba5_05130000,
        64'h2517f53f_f0ef9101,
        64'h02049513_2481eddf,
        64'hf0effb25_05130000,
        64'h25175064_d03c1040,
        64'h07932000_0437fff5,
        64'h37fd0001_47a9c3b8,
        64'h47292000_07b7f05f,
        64'hf0efe426_e822ec06,
        64'hfd250513_11010000,
        64'h25178082_41088082,
        64'hc10c8082_610560e2,
        64'hee1ff0ef_00914503,
        64'hee9ff0ef_00814503,
        64'hf55ff0ef_ec06002c,
        64'h11018082_61456942,
        64'h64e27402_70a2fe94,
        64'h10e3f0bf_f0ef0091,
        64'h4503f13f_f0ef3461,
        64'h00814503_f81ff0ef,
        64'h0ff57513_002c0089,
        64'h553354e1_03800413,
        64'h892af406_e84aec26,
        64'hf0227179_80826145,
        64'h694264e2_740270a2,
        64'hfe9410e3_f4dff0ef,
        64'h00914503_f55ff0ef,
        64'h34610081_4503fc3f,
        64'hf0ef0ff5_7513002c,
        64'h0089553b_54e14461,
        64'h892af406_e84aec26,
        64'hf0227179_808200f5,
        64'h80230007_c78300e5,
        64'h80a397aa_81110007,
        64'h4703973e_00f57713,
        64'h28078793_00001797,
        64'hb7f50405_fa5ff0ef,
        64'h80820141_640260a2,
        64'he5090004_4503842a,
        64'he406e022_11418082,
        64'h00e78823_02000713,
        64'h00e78423_fc700713,
        64'h00e78623_470d0007,
        64'h822300e7_8023476d,
        64'h00e78623_f8000713,
        64'h00078223_100007b7,
        64'h808200a7_0023dfe5,
        64'h0207f793_01474783,
        64'h10000737_80820205,
        64'h75130147_c5031000,
        64'h07b78082_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_58458593,
        64'h00001597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h2cc010ef_01a11113,
        64'h0210011b_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
