/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'h0000a617fec58593000005970d249063, /*    1 */
128'h011696933ff6869b000046b773c60613, /*    2 */
128'h0085b70300e6b0230005b70300d007b3, /*    3 */
128'h0185b70300e6b8230105b70300e6b423, /*    4 */
128'hfcc5cce3020686930205859300e6bc23, /*    5 */
128'h40b787b300d787b30147879300000797, /*    6 */
128'h305790730b4787930000079700078067, /*    7 */
128'h778585930000a59701b111130110011b, /*    8 */
128'h0005b4230005b023cb0606130000c617, /*    9 */
128'hfec5c6e3020585930005bc230005b823, /*   10 */
128'h0124a02300100913020004b7372080ef, /*   11 */
128'hff24c6e34009091b0200093700448493, /*   12 */
128'hfe090ae3008979133440297310500073, /*   13 */
128'h0099093300291913f1402973020004b7, /*   14 */
128'h00448493fe091ee30004a90300092023, /*   15 */
128'hf1402573ff24c6e34009091b02000937, /*   16 */
128'h3ff4849b000044b79805859300009597, /*   17 */
128'h34102373342022f30004806701149493, /*   18 */
128'h0000000000000000ffdff06f10500073, /*   19 */
128'h00000000000000000000000000000000, /*   20 */
128'h00000000000000000000000000000000, /*   21 */
128'h00000000000000000000000000000000, /*   22 */
128'h00000000000000000000000000000000, /*   23 */
128'h00000000000000000000000000000000, /*   24 */
128'h00000000000000000000000000000000, /*   25 */
128'h00000000000000000000000000000000, /*   26 */
128'h00000000000000000000000000000000, /*   27 */
128'h00000000000000000000000000000000, /*   28 */
128'h00000000000000000000000000000000, /*   29 */
128'h00000000000000000000000000000000, /*   30 */
128'h00000000000000000000000000000000, /*   31 */
128'hd963454c0005cc635735c28587ae6914, /*   32 */
128'he21c97b6470102a787b30a00051300b7, /*   33 */
128'h853e85b200030563018533038082853a, /*   34 */
128'h3d8686930000a697b7edfda007138302, /*   35 */
128'h87930000a7976294518707130000a717, /*   36 */
128'h87b30280069302d787bb878d8f9950e7, /*   37 */
128'h47148082853a470100e7956397ba02d7, /*   38 */
128'hf0efe4061141b7f502870713fea68de3, /*   39 */
128'hbfe545018082014160a26108c509fbbf, /*   40 */
128'hf0efe852ec4ef04af426f822fc067139, /*   41 */
128'h0000aa17440144814985892acd31f9bf, /*   42 */
128'hc091553500f44d6300c927831fca0a13, /*   43 */
128'h61216a4269e2790274a2744270e24501, /*   44 */
128'h67a2ed19f29ff0ef854a85a200308082, /*   45 */
128'h50ef8552000995632485cb990087c783, /*   46 */
128'h0513bf65240511c080ef498165224a20, /*   47 */
128'hf2dff0efe42ef406f0227179b7c1fda0, /*   48 */
128'h842aee7ff0ef083065a2c105fda00413, /*   49 */
128'h00f7096300c547030ff007936562e911, /*   50 */
128'h547980826145740270a285220e2080ef, /*   51 */
128'hf0efec4ef04af426f822fc067139bfd5, /*   52 */
128'h000099970ff00913440184aacd01eebf, /*   53 */
128'h74a2744270e200f4496344dc34498993, /*   54 */
128'hf0ef852685a200308082612169e27902, /*   55 */
128'h85a20127896300c7c78367a2ed09e83f, /*   56 */
128'hb7d9240507c080ef65223fe050ef854e, /*   57 */
128'he8dff0ef892eec26f406e84af0227179, /*   58 */
128'he45ff0ef84aa85ca0030c11dfda00413, /*   59 */
128'h2e85051300009517864a608ced01842a, /*   60 */
128'h740270a2852203e080ef65223c0050ef, /*   61 */
128'hf406ec26f022717980826145694264e2, /*   62 */
128'h85a6842ac11dfda00413e47ff0ef84ae, /*   63 */
128'hcf63445c388050ef2c05051300009517, /*   64 */
128'h5435004080ef2be505130000951700f4, /*   65 */
128'h003085228082614564e2740270a28522, /*   66 */
128'h7d9070ef6522f565842adcfff0ef85a6, /*   67 */
128'h5479fcf71be30ff0079300c7c70367a2, /*   68 */
128'he50965a2de1ff0eff406e42e7179bfc1, /*   69 */
128'hf96dd97ff0ef08308082614570a24501, /*   70 */
128'he42eec064108842ae8221101bfc56562, /*   71 */
128'h852200030e6302053303c919db9ff0ef, /*   72 */
128'h60e2fda005138302610560e265a26442, /*   73 */
128'h0000a7977139bfdd4501808261056442, /*   74 */
128'h04130000a417f426f822639c16478793, /*   75 */
128'h043b840d8c05296484930000a49729e4, /*   76 */
128'h892afc06e852ec4ef04a0280079302f4, /*   77 */
128'h942602f404331fea0a1300009a1789ae, /*   78 */
128'h69e2790274a2744270e2450100849b63, /*   79 */
128'h284050ef855285ca6090808261216a42, /*   80 */
128'hbfc902848493c501691060ef854a608c, /*   81 */
128'hb7e16522f569cdbff0ef852685ce0030, /*   82 */
128'h84b68432e42efc06f04af426f8227139, /*   83 */
128'hcb5ff0ef083065a2c115cf7ff0ef893a, /*   84 */
128'h70e2978285a2615c862686ca6562e519, /*   85 */
128'hbfc5fda0051380826121790274a27442, /*   86 */
128'h84b68432e42efc06f04af426f8227139, /*   87 */
128'hc75ff0ef083065a2c115cb7ff0ef893a, /*   88 */
128'h70e2978285a2655c862686ca6562e519, /*   89 */
128'hbfc5fda0051380826121790274a27442, /*   90 */
128'hc7dff0ef84b2e42ef822fc06f4267139, /*   91 */
128'h701ce509c39ff0ef842a083065a2c105, /*   92 */
128'h8082612174a2744270e2978285a66562, /*   93 */
128'h2785c3190017f713419cbfcdfda00513, /*   94 */
128'hd71b8e5927a106220086571b419cc19c, /*   95 */
128'h0ff77713c19c0087d7138ed906a20086, /*   96 */
128'h122300d5112300c510238fd90087979b, /*   97 */
128'hf022f4067179419c80820005132300f5, /*   98 */
128'h419c00f510230457879b6785c19c27d1, /*   99 */
128'h0087979b0ff777130087d713c632842a, /*  100 */
128'hc4360509084c57fd460900f11a238fd9, /*  101 */
128'h051301610593460977f060ef00f11b23, /*  102 */
128'h00041323082c462147c1771060ef0044, /*  103 */
128'h00f404a347c575d060efec3e00840513, /*  104 */
128'h747060ef00c4051300041523006c4611, /*  105 */
128'h0144069373b060ef01040513002c4611, /*  106 */
128'hfed79ce39f31ffe7d6030789470187a2, /*  107 */
128'h9fb94107d71b9fb9934117424107579b, /*  108 */
128'h80826145740270a200f41523fff7c793, /*  109 */
128'h97ba46a167856398038787930000a797, /*  110 */
128'hc7bb27850077e793fff6079b8007bc23, /*  111 */
128'h3823973e678500f547636805450102d7, /*  112 */
128'h010686bb0035169b0005b883808280c7, /*  113 */
128'he0221141bff105a125050116b02396ba, /*  114 */
128'hfa5ff0efe406450185aa86220005841b, /*  115 */
128'hec26f022717980820141640260a28522, /*  116 */
128'h687060efe436f4064619051984b2842a, /*  117 */
128'h162347a167b060ef85b64619852266a2, /*  118 */
128'h614564e200e4859b70a27402852200f4, /*  119 */
128'h3a8130236785737dc5010113fadff06f, /*  120 */
128'h3931342338913c233a11342339213823, /*  121 */
128'h377134233761382337513c2339413023, /*  122 */
128'h3507879335a1382335913c2337813023, /*  123 */
128'hce042023d00007b7943e747d978a911a, /*  124 */
128'hd0040023f0040023e0040023ca040b23, /*  125 */
128'h951785aa00e7ea63892a5800073797aa, /*  126 */
128'h00054703a00179b040eff02505130000, /*  127 */
128'h970a3507871374fd678526f711634789, /*  128 */
128'hcb848b13970a350787139abacd848a93, /*  129 */
128'h9c3a9b3a49818a368cb28baed0048c13, /*  130 */
128'hc7830015cd03013907b395ca0f098593, /*  131 */
128'h869b01a989bb058902a0071329890f07, /*  132 */
128'h24e78163471904f76b6326e78d630007, /*  133 */
128'hcc848513470d2ae78963470502f76263, /*  134 */
128'h40efff2505130000951785b622e78963, /*  135 */
128'hfee794e3473d22e785634731b77d7130, /*  136 */
128'h953e866ae0048513978a350787936785, /*  137 */
128'h03600713b759e00d0023541060ef9d22, /*  138 */
128'h22e780630330071300f76e6322e78363, /*  139 */
128'haad94605cb648513fae798e303500713, /*  140 */
128'hf8e79ce30ff0071324e7856303800713, /*  141 */
128'h24e781630007859b747d471500614783, /*  142 */
128'h000ca7833ae79063470936e784634719, /*  143 */
128'h05134985978a350a87936a8516079263, /*  144 */
128'h60ef013ca023953e461101090593ce44, /*  145 */
128'h01490593ce840513978a350a87934c50, /*  146 */
128'hdd850513000095174af060ef953e4611, /*  147 */
128'h978a350a879364b040efde0254e25a52, /*  148 */
128'h435060ef854a55fd4619993ecf840913, /*  149 */
128'h879346f115231350079300f103a3478d, /*  150 */
128'h85a6460594becb740493c2a6978a350a, /*  151 */
128'h06a30320079345d060efc0d246c10513, /*  152 */
128'h4a1195becf040593978a350a879346f1, /*  153 */
128'h0793439060ef4741072346f105134611, /*  154 */
128'hcf440593978a350a879346f109a30360, /*  155 */
128'h417060ef47410a2347510513461195be, /*  156 */
128'h03a346f10ca347b1051385a6460557fd, /*  157 */
128'h0613102007933fd060ef47310d230001, /*  158 */
128'h0793397060efde3e37a1051345810f00, /*  159 */
128'h3961051385de4799464136f11d231010, /*  160 */
128'h13232637879377e13cf060ef36f10e23, /*  161 */
128'h350a879346f1142335378793679946f1, /*  162 */
128'h0440061304300693943ecec40413978a, /*  163 */
128'h85a2460156fdba1ff0ef3721051385a2, /*  164 */
128'h0e8885de86ca5672bd5ff0ef35e10513, /*  165 */
128'h3a0134033a813083911a6305cebff0ef, /*  166 */
128'h38013a03388139833901390339813483, /*  167 */
128'h36013c0336813b8337013b0337813a83, /*  168 */
128'h851380823b01011335013d0335813c83, /*  169 */
128'ha00d953e978a3507879367854611cd04, /*  170 */
128'h953e866af0048513978a350787936785, /*  171 */
128'h85564611b39df00d0023321060ef9d22, /*  172 */
128'h87936785bfdd855a4611bbb1313060ef, /*  173 */
128'h2f7060ef4611953ece048513978a3507, /*  174 */
128'h00f40123ce14478300f401a3ce044783, /*  175 */
128'h00f40023ce34478300f400a3ce244783, /*  176 */
128'h866ab759cc048513bb29cef42023401c, /*  177 */
128'h2783b311d00d00232bf060ef9d228562, /*  178 */
128'h0000951700fa2023478510079d63000a, /*  179 */
128'h0e8801090593461144d040efbec50513, /*  180 */
128'hcb840513978a350487936485293060ef, /*  181 */
128'h3531470327b060ef014905934611953e, /*  182 */
128'h00009517350145833511460335214683, /*  183 */
128'h00a146833501578340d040efbbc50513, /*  184 */
128'h35215783ccf71e230000a71700914603, /*  185 */
128'h0000a717bbc505130000951700814583, /*  186 */
128'h01b147033d9040ef00b14703ccf71323, /*  187 */
128'h00009517018145830191460301a14683, /*  188 */
128'h01214683013147033bd040efbbc50513, /*  189 */
128'hbc050513000095170101458301114603, /*  190 */
128'h05130000951755c2010157833a1040ef, /*  191 */
128'ha71701215783c6f713230000a717bce5, /*  192 */
128'h978a3504879337b040efc4f71e230000, /*  193 */
128'h40efbba505130000951795bee0040593, /*  194 */
128'h951795be978af0040593350487933630, /*  195 */
128'h00009517bd2934b040efbb2505130000, /*  196 */
128'h93e3000a2783b53133d040efbb450513, /*  197 */
128'hba8505130000951700fa20234785e007, /*  198 */
128'h315040efbac5051300009517321040ef, /*  199 */
128'h951795be978ad0040593350787936785, /*  200 */
128'hbb85051300009517bf45bb2505130000, /*  201 */
128'he4a6e8a2ec86711d737db3c12f1040ef, /*  202 */
128'h00009517911a89aaf456f852fc4ee0ca, /*  203 */
128'h8793747d2c9040efca026a85bcc50513, /*  204 */
128'h852655fd461994beff840493978a020a, /*  205 */
128'h0913439ca1c787930000a7970b1060ef, /*  206 */
128'h879312f11d2313500793c83e4a05fef4, /*  207 */
128'h014107a31a68460585ca993e978a020a, /*  208 */
128'h0f23479112f10ea3037007930d3060ef, /*  209 */
128'h461195beff040593978a020a879312f1, /*  210 */
128'h0513460585ca57fd0af060ef13f10513, /*  211 */
128'h60ef000107a31541022314f101a31451, /*  212 */
128'h04a1051345810f0006130fc007930950, /*  213 */
128'h85ce04f115231010079302f060efca3e, /*  214 */
128'h067060ef04f106230661051346414799, /*  215 */
128'h35378793679912f11b232637879377e1, /*  216 */
128'h85a2943e1451978a020a879312f11c23, /*  217 */
128'h83bff0ef044006130430069304210513, /*  218 */
128'h465286fff0ef460156fd02e1051385a2, /*  219 */
128'h60e6911a6305985ff0ef85ce86a61008, /*  220 */
128'h61257aa27a4279e2690664a664464501, /*  221 */
128'h1a50406fabc505130000951785aa8082, /*  222 */
128'h7c913c237e8130237e11342381010113, /*  223 */
128'h05a1051384aa71597d3134237d213823, /*  224 */
128'h60efd602e83eec3ae442893689b2e046, /*  225 */
128'h6762747d97ba81078793101867857c40, /*  226 */
128'h0521051385a2864a86ba943e7fc40413, /*  227 */
128'h863e86c285a267c26822fa4ff0efd64e, /*  228 */
128'h85a6180856326882fd4ff0ef03e10513, /*  229 */
128'h340345017e81308361658e9ff0ef86c6, /*  230 */
128'h01137c8139837d0139037d8134837e01, /*  231 */
128'h480300554883e222e606716d80827f01, /*  232 */
128'h46030015468300254703003547830045, /*  233 */
128'h00009517a0c5859300009597842a0005, /*  234 */
128'h842adedff0ef85220dd040efa0c50513, /*  235 */
128'h000095179ec5859300009597860ac10d, /*  236 */
128'h6151641260b285220bd040efa1450513, /*  237 */
128'hab230000a797a2e50513000095178082, /*  238 */
128'he4ceeca6f0a27159b7cd09f040ef9007, /*  239 */
128'hf486e86aec66f062f45ef85afc56e0d2, /*  240 */
128'h9a974401ff05049389ae8a2ae46ee8ca, /*  241 */
128'h0b93a02b0b1300009b17a2aa8a930000, /*  242 */
128'h8c9300009c97a0ec0c1300009c170600, /*  243 */
128'h64e6740670a603344163fff58d1b9fec, /*  244 */
128'h6ce27c027ba27b427ae26a0669a66946, /*  245 */
128'he7a9c42900f47793808261656da26d42, /*  246 */
128'hc583012487b34dc1490101f040ef855a, /*  247 */
128'h856602fbe2630ff7f793fe05879b0007, /*  248 */
128'h051300009517ffb912e30905001040ef, /*  249 */
128'h8562a0317e8040ef85567ee040ef50e5, /*  250 */
128'h000095170104c583dbe5b7c57e0040ef, /*  251 */
128'hfffd4913028d1d637cc040ef99450513, /*  252 */
128'h2d857b6040ef8556a02900f979134d81, /*  253 */
128'h079bff0479137aa040ef855aff2dcce3, /*  254 */
128'h40ef4b2505130000951700f45b630009, /*  255 */
128'h0007c583012a07b3b781048524057920, /*  256 */
128'h40ef856600fbe7630ff7f793fe05879b, /*  257 */
128'h7179bfdd768040ef8562b7e909057720, /*  258 */
128'h893289ae84b6f022f406e44ee84aec26, /*  259 */
128'h869300009697c5091e06869300009697, /*  260 */
128'h061300009617a16707130000871790e6, /*  261 */
128'h00098f63842a6ea040ef854a85a69066, /*  262 */
128'h06130000961786ce40a485bb00955d63, /*  263 */
128'h4463ffe4879b9c296cc040ef954a8ee6, /*  264 */
128'h85930000959700890533ffd4841b00f4, /*  265 */
128'h694264e2854a740270a2284060ef8be5, /*  266 */
128'hf73ff06f4581862e86b28082614569a2, /*  267 */
128'hfebff0efed8645050c800613002c7115, /*  268 */
128'h60ee6b6040ef8a65051300009517002c, /*  269 */
128'h862e9ff787133b9ad7b78082612d4501, /*  270 */
128'h04a7676323f78713000f47b704a76963, /*  271 */
128'h97173e80079346890ca7f7633e700793, /*  272 */
128'h00074903e04a97361101602707130000, /*  273 */
128'h64a260e2644202091663e426e822ec06, /*  274 */
128'h406f610584c505130000951785aa6902, /*  275 */
128'h240787934685b7d9a007879346816520, /*  276 */
128'h3e800793c02102f555b302f57433bf7d, /*  277 */
128'h0713c70502f4773347a90287e6634729, /*  278 */
128'h743302f457b306400713028774630630, /*  279 */
128'h5433a039943e001444130324341302e4, /*  280 */
128'h051300008517f86102f45433bfc102e4, /*  281 */
128'h0000851785a2c8015ec040ef84b27f65, /*  282 */
128'h85ca862660e264425dc040ef7ec50513, /*  283 */
128'h406f61057dc5051300008517690264a2, /*  284 */
128'h862eb78d7ac505130000851785aa5c20, /*  285 */
128'h55b303c6871b02f886bb481958d94781, /*  286 */
128'h510808130000981793811782cd8500e5, /*  287 */
128'he04ae822ec060007c483e42697c21101, /*  288 */
128'h0000851785aa690264a260e26442e495, /*  289 */
128'hfb079de3278556a0406f610578c50513, /*  290 */
128'h97b357fdb7f5776505130000851785aa, /*  291 */
128'h053347a9c10d44018d7dfff7c79300e7, /*  292 */
128'h942a47a500d41433440503b6869b02f5, /*  293 */
128'h00008517058514590087f46300e45433, /*  294 */
128'h851785a2c80151a040ef893272450513, /*  295 */
128'h864a60e2644250a040ef71a505130000, /*  296 */
128'h6105722505130000851764a2690285a6, /*  297 */
128'hf1a202c7073b8cbaed6671514f00406f, /*  298 */
128'hf95afd56e1d2eda6f586e96ae5cee9ca, /*  299 */
128'h8d3289ae892a04000793e56ef162f55e, /*  300 */
128'h956302ccdcbb04000c9300e7f6638436, /*  301 */
128'h020d1a13001d179b03acdcbb4cc1000c, /*  302 */
128'h8b1703810a93020a5a130017849be03e, /*  303 */
128'h7c1762ab8b9300008b976cab0b130000, /*  304 */
128'h64ee740e70ae4501e00d1f2c0c130000, /*  305 */
128'h6cea7c0a7baa7b4a7aea6a0e69ae694e, /*  306 */
128'h05130000851785ca8082616d6daa6d4a, /*  307 */
128'h8d9b008cf46300040d9b44e040ef6865, /*  308 */
128'h0007061b430948a14811470186ce000c, /*  309 */
128'h99ba034707339301020d971305b66c63, /*  310 */
128'h861b02e00813875603bd06bb0d9de663, /*  311 */
128'h85d6963e011c0ac5ed63415705bb0006, /*  312 */
128'h40effa060c23e4366405051300008517, /*  313 */
128'h60ef99369281168241b4043b66a23f20, /*  314 */
128'h15934290030d1b63b795557dd1357c70, /*  315 */
128'h855a658292011602c190260195d60027, /*  316 */
128'h66a23b6040efe436e83aec42f046f41a, /*  317 */
128'h1863bf8568627882070596d273226742, /*  318 */
128'h1c63bfc1e19095d6003715936290011d, /*  319 */
128'h9241164295d6001715930006d603006d, /*  320 */
128'h761300ea85b30006c603bf6500c59023, /*  321 */
128'h7f3060efe43a855eb75d00c580230ff6, /*  322 */
128'hbfdd4701bf1d3cfdfe976ae327056722, /*  323 */
128'h097575130005450300bc053300074583, /*  324 */
128'h00230005d4634185d59b0185959bc519, /*  325 */
128'hf4634501918187aa1582bf3907050107, /*  326 */
128'h04000793bfd58f8d25058082e21c00b7, /*  327 */
128'h57f70713464c47370005668312b7f463, /*  328 */
128'h10e6976347090045468310e69c634789, /*  329 */
128'hf0a202f7073371590380079303855703, /*  330 */
128'he4cee8caeca6f48602059a93fc567100, /*  331 */
128'hda93e46ee86aec66f062f45ef85ae0d2, /*  332 */
128'h942a84aa892e06eae663478d9722020a, /*  333 */
128'h00008c174f4b8b9300008b974b054a01, /*  334 */
128'h0384d783514c8c9300008c97534c0c13, /*  335 */
128'h741c09679b63401ca835478100fa6463, /*  336 */
128'h8d630204398327a040ef855e85d2cbc1, /*  337 */
128'hfa6395ce00b48db301843d03640c0409, /*  338 */
128'h254040ef4b45051300008517864a02ba, /*  339 */
128'h7ae26a0669a6694664e6740670a6478d, /*  340 */
128'h6165853e6da26d426ce27c027ba27b42, /*  341 */
128'h864e226040ef856686ce85ea866e8082, /*  342 */
128'hf163701c0284398306e060ef856a85ee, /*  343 */
128'h85ea9d3e864e40f989b301843d030337, /*  344 */
128'h7f5050ef856a4581864e1fe040ef8562, /*  345 */
128'h45058082853e4785bf99038404132a05, /*  346 */
128'h0713000097178082400005378082057e, /*  347 */
128'h95360017869300756513157d631c26e7, /*  348 */
128'h8082953e057e450597aa20000537e308, /*  349 */
128'h08a74463862a0ce50763820787136785, /*  350 */
128'h06e60b63454505130000851780878713, /*  351 */
128'h43050513000085178006079b04c74963, /*  352 */
128'h4b0505130000851787f787936785c3ad, /*  353 */
128'h85979e3d11417c07879b77fd04c7c963, /*  354 */
128'he4061d250513000095174a2585930000, /*  355 */
128'h01411c2505130000951760a212c040ef, /*  356 */
128'h0a634025051300008517810787138082, /*  357 */
128'h12e340250513000085178187879300e6, /*  358 */
128'h4205051300008517830787138082faf6, /*  359 */
128'h000085178287879300c74963fee609e3, /*  360 */
128'h05130000851783878713bfe93fc50513, /*  361 */
128'h05130000851784078793fce608e340e5, /*  362 */
128'h717980823c45051300008517bf7540e5, /*  363 */
128'h4463440184ae892af406e84aec26f022, /*  364 */
128'h01045513942a90411442010455130290, /*  365 */
128'h694264e21542fff54513740270a29522, /*  366 */
128'h6e7050ef0068460985ca808261459141, /*  367 */
128'h00d1478300f107a334f9090900c14783, /*  368 */
128'h6785715dbf55943e00e1578300f10723, /*  369 */
128'h842e80678793f44ef84afc26e486e0a2, /*  370 */
128'h079b0af50e636dd7879367a13cf50563, /*  371 */
128'h50ef4611082884b205e944079a638005, /*  372 */
128'h051300009517461985ca006409136950, /*  373 */
128'h896302e0079301744583681050ef0c65, /*  374 */
128'h04b7e5631cf5826347b108b7e76332f5, /*  375 */
128'h10f58463478502b7e3631af583634791, /*  376 */
128'h851702f5836334e50513000085174789, /*  377 */
128'h82634799a41d7eb030ef4ea505130000, /*  378 */
128'hfef591e3354505130000851747a118f5, /*  379 */
128'h00b7ed632cf5826347f5a4317d1030ef, /*  380 */
128'h370505130000851747d916f58a6347c5, /*  381 */
128'h07932af5866302100793bf6dfef580e3, /*  382 */
128'hb7c938a5051300008517faf596e30290, /*  383 */
128'h0330079304b7e2632cf5826306200793, /*  384 */
128'h28f5876302f0079300b7ef632af58263, /*  385 */
128'hf8f58ae338c505130000851703200793, /*  386 */
128'h851705e0079328f5846305c00793b7bd, /*  387 */
128'h08400793bf91f6f58de33a2505130000, /*  388 */
128'h26f58b630670079300b7ef6328f58663, /*  389 */
128'hf4f58ae33b4505130000851706c00793, /*  390 */
128'h89630ff0079326f5886308900793b73d, /*  391 */
128'h051300008517f0f59ce30880079326f5, /*  392 */
128'hfd87d7830000979701e45703b73d3be5, /*  393 */
128'h0204570312f71463fd09899300009997, /*  394 */
128'h85ca461910f71c63fc27d78300009797, /*  395 */
128'hf9058593000095974619521050ef8522, /*  396 */
128'h12230204012301a45783511050ef854a, /*  397 */
128'h0513fde4859b01c4578300f41f230204, /*  398 */
128'hd78300f41d230009d78302f410230224, /*  399 */
128'h812100a10ea3db9ff0ef00f41e230029, /*  400 */
128'h85a202f41223862601c1578300a10e23, /*  401 */
128'h1c05051300008517a06ddbffe0ef4501, /*  402 */
128'h00008517b5591ce5051300008517bd41, /*  403 */
128'h0ea30264470302444783bdb51dc50513, /*  404 */
128'h0ea301c1178300f10e230254478300f1, /*  405 */
128'h0224470300e10e2327810274470300e1, /*  406 */
128'h00e10e230234470300e10ea301c11903, /*  407 */
128'h0000979704e79b6301c1568304500713, /*  408 */
128'he885859300009597461947e2ead79823, /*  409 */
128'he8f7282300009717e905051300009517, /*  410 */
128'h87930000979766a24762431050efe436, /*  411 */
128'h4d6060ef450102a40593ff89061be667, /*  412 */
128'h07138082616179a2794274e2640660a6, /*  413 */
128'he4f728230000971747e204e694630430, /*  414 */
128'h00009797c799439ce547879300009797, /*  415 */
128'he386869300009697f7e9439ce4478793, /*  416 */
128'he385859300009597e346061300009617, /*  417 */
128'h98634d200713b765d61fe0ef02a40513, /*  418 */
128'h85a6557030ef0f6505130000851702e7, /*  419 */
128'h30ef0f25051300008517cb6ff0ef8522, /*  420 */
128'h0713bf95ca0ff0ef02a4051385ca5430, /*  421 */
128'h01e317fd67c101e45703f6e787e35fe0, /*  422 */
128'h000095974611f4f70de302045703f6f7, /*  423 */
128'h00008517b79935d050ef0868df458593, /*  424 */
128'hb30d0d25051300008517b3350cc50513, /*  425 */
128'h051300008517bb210e85051300008517, /*  426 */
128'h8517b31110c5051300008517b3390f65, /*  427 */
128'h1305051300008517b9ed112505130000, /*  428 */
128'h00008517b1dd13e5051300008517b9c5, /*  429 */
128'hb9c917a5051300008517b9f115450513, /*  430 */
128'h97970265d703b1e11885051300008517, /*  431 */
128'h11e3d6a4849300009497d727d7830000, /*  432 */
128'h19e3d5c7d783000097970285d703ecf7, /*  433 */
128'h9a23016589930205891320000793eaf7, /*  434 */
128'h959746192ab050ef854a85ce461900f5, /*  435 */
128'h9597461929b050ef854ed1a585930000, /*  436 */
128'h4619289050ef00640513d0a585930000, /*  437 */
128'h02a0061301c4578327f050ef852285ca, /*  438 */
128'h0004d78302f4142301e4578302f41323, /*  439 */
128'h6080079300f41f230024d78300f41e23, /*  440 */
128'h110505130000851785aab36900f41623, /*  441 */
128'h8307b603300017b7bba546013f1030ef, /*  442 */
128'h171b00f674132601608130239f010113, /*  443 */
128'h05379f2d8406871b0387759366850034, /*  444 */
128'h34235e913c23630c8387b783972a3000, /*  445 */
128'h696335b95f200813ffc5849b25816011, /*  446 */
128'hfff7c79300c5963b101005938a1d08b8, /*  447 */
128'h4390c427879300009797cfb527818ff1, /*  448 */
128'h9ebd8006869b7007f7930084179bea25, /*  449 */
128'h0106969b00d100a3872646d496aa068e, /*  450 */
128'h0001550300d100230086d69b0106d69b, /*  451 */
128'h02d51a63806686936685c6918005069b, /*  452 */
128'h46a1007767139fad377d8005859b6585, /*  453 */
128'h08378f95868a83f502d7473b17822705, /*  454 */
128'haa1ff0ef862602e6446397c285b63000, /*  455 */
128'h3403608130838287b823300017b70405, /*  456 */
128'h88338082610101135f81348385266001, /*  457 */
128'hb7e1ff06bc2306a126050008380300d7, /*  458 */
128'h2401ec06e42643c0e8220c2007b71101, /*  459 */
128'hc163033716938304b703300014b74781, /*  460 */
128'h2b5030effec5051300008517e7990206, /*  461 */
128'h8082610564a2644260e2c3c00c2007b7, /*  462 */
128'h8432ec26f0227179bfc14785eb9ff0ef, /*  463 */
128'hf4060068b6c5859300009597461184ae, /*  464 */
128'h0007a803b2478793000097970d3050ef, /*  465 */
128'h9717b0a888930000989785a6862247b2, /*  466 */
128'h05130000951704500693b0e757030000, /*  467 */
128'h614564e2740270a285228aeff0efb165, /*  468 */
128'h8082914115428d5d05220085579b8082, /*  469 */
128'hf00686938fd966c10185579b0185171b, /*  470 */
128'h00ff07370085151b8fd98f750085571b, /*  471 */
128'h051300008517715d808225018d5d8d79, /*  472 */
128'hec56f052f44ef84afc26e0a2e486f4e5, /*  473 */
128'h47e1aa078523000097971ef030efe85a, /*  474 */
128'h0000971703e00793aaf700a300009717, /*  475 */
128'h578da8f706a3000097174789a8f70b23, /*  476 */
128'h959707f007934611a8f7022300009717, /*  477 */
128'ha6840413000094170028a74585930000, /*  478 */
128'h85a246097ea050efa6f702a300009717, /*  479 */
128'h899300009997448145227e0050ef0068, /*  480 */
128'hf00606130100063746b2f4fff0efa2e9, /*  481 */
128'h15028f558f710ff6f69382a10086971b, /*  482 */
128'hb423934180a7b02317429101300017b7, /*  483 */
128'h0513000085178087b7038007b70380e7, /*  484 */
128'h8087b5838007b60382e7b4234721e9e5, /*  485 */
128'h91c115c29dca0a1300009a1700800737, /*  486 */
128'h47030000971711b030ef80e7b4238f4d, /*  487 */
128'h4803000098179d27c783000097979d97, /*  488 */
128'h4603000096179c06c683000096979cb8, /*  489 */
128'h0513000085179ae5c583000095979b76, /*  490 */
128'h00989b376a89000447830df030efe4e5, /*  491 */
128'h300019370014478398f70c2300009717, /*  492 */
128'h000097170024478398f704a300009717, /*  493 */
128'h96f709a3000097170034478396f70f23, /*  494 */
128'h0054478396f704230000971700444783, /*  495 */
128'h92079a230000979794f70ea300009717, /*  496 */
128'h9207a823000097979207a42300009797, /*  497 */
128'h9007ac23000097979207a22300009797, /*  498 */
128'h0493f4bfe0ef8522e78d0009a783e4a9, /*  499 */
128'h3783020745630337971383093783680b, /*  500 */
128'hbfc5c4fff0effc075de3033797138309, /*  501 */
128'h849378d050ef4501dff154fd000a2783, /*  502 */
128'h17b7b7d914fdb7e9c35ff0efbfc1710a, /*  503 */
128'he40616fd1141ff8006b78087b7033000, /*  504 */
128'h82e7b823f0070713670580e7b4238f75, /*  505 */
128'h7e4030efd8450513000085178307b583, /*  506 */
128'h300027f37d8030efda05051300008517, /*  507 */
128'h07fe4785300790738fd9880707136709, /*  508 */
128'h7b4030efd9c505130000851734179073, /*  509 */
128'h47838082014160a2302000730000100f, /*  510 */
128'h4503002547838f5d07a2000547030015, /*  511 */
128'h57fd808225018d5d05628fd907c20035, /*  512 */
128'h058505050005c703808200f61363367d, /*  513 */
128'h808200f61363367d57fdb7f5fee50fa3, /*  514 */
128'hec06e8221101495cbfcd050500b50023, /*  515 */
128'h478101853903cfa500958413e04ae426, /*  516 */
128'h462d02e0031348a5481586ca02000513, /*  517 */
128'h07130107146300a70e6327850006c703, /*  518 */
128'h00e40023040500640023011795630e50, /*  519 */
128'h01c9051300b94783fcc79ee306850405, /*  520 */
128'h01994783c088f59ff0ef00f5842384ae, /*  521 */
128'h478300f492238fd90087979b01894703, /*  522 */
128'h00f493238fd90087979b016947030179, /*  523 */
128'h80826105690264a2644260e200040023, /*  524 */
128'h468303a0061302000593cf99873e611c, /*  525 */
128'h06630017869300c6986302d5fc630007, /*  526 */
128'h46050007c683b7dd0705a00d577d00d7, /*  527 */
128'h078900b666630ff6f593fd06869b577d, /*  528 */
128'h4703000087178082853ae11c0006871b, /*  529 */
128'hc70d0007c703cb85611cc915bfd576e7, /*  530 */
128'he406114102e69063008557030067d683, /*  531 */
128'hc3914501001577932c8060ef0017c503, /*  532 */
128'h01b5c783808245258082014160a24525, /*  533 */
128'h0007079b8f5d0087979b468d01a5c703, /*  534 */
128'h0087979b0145c6830155c78300d51d63, /*  535 */
128'h71798082853e27818fd90107979b8fd5, /*  536 */
128'h0993e052e84af4065904e44eec26f022, /*  537 */
128'h60ef85ce8626468500154503842a0345, /*  538 */
128'h87bb000402234c58505ce13125012560, /*  539 */
128'h694264e2740270a2450100e7eb6340f4, /*  540 */
128'h74e34a0500344903808261456a0269a2, /*  541 */
128'h85ce86269cbd4685001445034c5cff2a, /*  542 */
128'h00454783b7f94505b7e5397d214060ef, /*  543 */
128'he8221101591c80824501f8dff06fc399, /*  544 */
128'h892e84aa02b787634401e04ae426ec06, /*  545 */
128'h46850014c503ec190005041bfddff0ef, /*  546 */
128'h4405c119250119c060ef03448593864a, /*  547 */
128'h690264a2644260e285220324a823597d, /*  548 */
128'h57fde04ae426ec06e822110180826105, /*  549 */
128'he52d2501fa3ff0ef842ad91c00050223, /*  550 */
128'h8fd90087979b45092324470323344783, /*  551 */
128'h1f63a55707134107d79b776d0107979b, /*  552 */
128'h05370005079bd59ff0ef06a4051302f7, /*  553 */
128'hf7b31465049300544537fff509130100, /*  554 */
128'hd33ff0ef0864051300978c6345010127, /*  555 */
128'h644260e200a035338d05012575332501, /*  556 */
128'hf84a715dbfcd450d80826105690264a2, /*  557 */
128'h3023e85aec56f052fc26e0a2e486f44e, /*  558 */
128'h4e6347addd9ff0ef8932852e89aa0005, /*  559 */
128'h97ba5727879300008797003517130205, /*  560 */
128'h000447830089b023c01547b184aa6380, /*  561 */
128'he38d001577930e6060ef00144503cb85, /*  562 */
128'h74e2640660a647a9c111891100090563, /*  563 */
128'h80826161853e6b426ae27a0279a27942, /*  564 */
128'h7f9050ef00a400a3000400230ff4f513, /*  565 */
128'hf569891100090463fb71478d00157713, /*  566 */
128'h848a04f51a634785ee1ff0ef85224581, /*  567 */
128'h4501ffc9478389a623a40a131fa40913, /*  568 */
128'h094100a9a0232501c5bff0ef854ac789, /*  569 */
128'h45090004aa8301048913ff2a14e30991, /*  570 */
128'h0491c10de9dff0ef852285d6000a8763, /*  571 */
128'h470db7bd00e519634785470dfe9915e3, /*  572 */
128'h4783bfb947b5c1194a81f6e504e34785, /*  573 */
128'h0107979b8fd90087979b03f447030404, /*  574 */
128'h04b44983fef711e3200007134107d79b, /*  575 */
128'h1a09866300f9e9b30089999b04a44783, /*  576 */
128'hfff9079b470501342e23044449032981, /*  577 */
128'h04144b03faf769e30ff7f793012401a3, /*  578 */
128'h00fb77b3fffb079bfa0b03e301640123, /*  579 */
128'h6a33008a1a1b0454478304644a03ffc9, /*  580 */
128'h04844503f3c100fa77930144142300fa, /*  581 */
128'h478314050e638d450085151b04744483, /*  582 */
128'hdfb18fd90087979b2501042447030434, /*  583 */
128'h00d7063b9f3d004a571b2781033906bb, /*  584 */
128'h84ae0364d5bb40c504bbf4c564e38732, /*  585 */
128'h0905165500b93933664119556905dd8d, /*  586 */
128'h015787bb248900ea873b490d00b67363, /*  587 */
128'h10e91263470dd05c03542023cc04d458, /*  588 */
128'h949bd408b17ff0ef06040513f00a15e3, /*  589 */
128'hee99e7e324810094d49b1ff4849b0024, /*  590 */
128'h478d00f402a3f8000793c45cc81c57fd, /*  591 */
128'h0087979b064447030654478308f91963, /*  592 */
128'h06f71b6347054107d79b0107979b8fd9, /*  593 */
128'h4783e13d2501ce5ff0ef8522001a859b, /*  594 */
128'h8fd90087979b000402a3232447032334, /*  595 */
128'h1263a55707134107d79b776d0107979b, /*  596 */
128'h2501416157b7a99ff0ef0344051304f7, /*  597 */
128'ha83ff0ef2184051302f5176325278793, /*  598 */
128'h051300f51c63272787932501614177b7, /*  599 */
128'ha63ff0ef22040513c808a6dff0ef21c4, /*  600 */
128'h93c117c227852f87d78300008797c448, /*  601 */
128'h0124002300f413232ef7152300008717, /*  602 */
128'ha33ff0ef05840513b351478100042a23, /*  603 */
128'hb545a25ff0ef05440513b5b90005099b, /*  604 */
128'h949b00f915634789d41c9fb5e00a05e3, /*  605 */
128'h0017d79b8885029787bb478db7010014, /*  606 */
128'hf0ef842ae426ec06e8221101bdc59cbd, /*  607 */
128'h0cf71063478d00044703ed692501bfff, /*  608 */
128'h0613034404930af71b63478500544703, /*  609 */
128'h092305500793a01ff0ef852645812000, /*  610 */
128'h0a230520079322f409a3faa0079322f4, /*  611 */
128'h0da302f40b230610079302f40aa302f4, /*  612 */
128'h20e40d2302e40ba304100713481c20f4, /*  613 */
128'h20f40e230087571b0107571b0107971b, /*  614 */
128'h20f40fa30187d79b0107d71b20e40ea3, /*  615 */
128'h0107571b0107971b501020e40f23445c, /*  616 */
128'h22f4002307200693001445030087571b, /*  617 */
128'h0c230187d79b0107d71b260522e400a3, /*  618 */
128'hd81022f401a322e4012320d40ca320d4, /*  619 */
128'h00144503000402a3541050ef85a64685, /*  620 */
128'h60e200a035332501535050ef45814601, /*  621 */
128'h37f9ffe5869b4d1c8082610564a26442, /*  622 */
128'h9d2d02d585bb55480025458300f6f963, /*  623 */
128'h71794d180eb7f7634785808245018082, /*  624 */
128'h02e5f963892ae44eec26f022f406e84a, /*  625 */
128'h0e63468d06d70c63842e468900054703, /*  626 */
128'hd59b9cad515c0015d49b00f71e6308d7, /*  627 */
128'h70a257fdc9112501ac7ff0ef9dbd0094, /*  628 */
128'h278380826145853e69a2694264e27402, /*  629 */
128'h94ca1ff4f4930099d59b0014899b0249, /*  630 */
128'hf5792501a93ff0ef0344c483854a9dbd, /*  631 */
128'h0087979b880503494783994e1ff9f993, /*  632 */
128'hbf458fe9157d6505bf658391c0198fc5, /*  633 */
128'hfd592501a63ff0ef9dbd0085d59b515c, /*  634 */
128'h45030359478399221fe474130014141b, /*  635 */
128'h0075d59b515cb7598fc90087979b0349, /*  636 */
128'h75130024151bf9352501a39ff0ef9dbd, /*  637 */
128'h100007b7807ff0ef954a034505131fc5, /*  638 */
128'hf82271398082853e4785b76517fd2501, /*  639 */
128'h1523e456e852ec4ef426fc06f04a4540, /*  640 */
128'h744270e2450900f41c63892a478500b5, /*  641 */
128'h611c808261216aa26a4269e2790274a2, /*  642 */
128'h470d0007c683e02184aefee474e34f98, /*  643 */
128'hfce4f7e30087d703eb15579800e69463, /*  644 */
128'h37839d3d0044d79bd171008928235788, /*  645 */
128'h00a92a2394be03478793049688bd0009, /*  646 */
128'h843a0027c9838722b75d450100993c23, /*  647 */
128'h0134f66385a2000935034a8509925a7d, /*  648 */
128'h0005041be6fff0efbf752501e59ff0ef, /*  649 */
128'h76e34f9c00093783f68afbe301440c63, /*  650 */
128'h00a55583b78d4505bfc1413484bbf6f4, /*  651 */
128'h049bf33ff0ef842aec06e426e8221101, /*  652 */
128'h0005049b933ff0ef6008484ce4950005, /*  653 */
128'h6c1cf3cff0ef4581020006136c08ec99, /*  654 */
128'h60e200e782234705601c00e780235715, /*  655 */
128'hfc06e85271398082610564a285266442, /*  656 */
128'h16ba75634a05e456ec4ef04af426f822, /*  657 */
128'h4709000547830af5f063498984aa4d1c, /*  658 */
128'h94630ee78863470d0ae78f63842e8932, /*  659 */
128'h009a559b00ba0a3b515c0015da1b1547, /*  660 */
128'h8805060996630005099b8b9ff0ef9dbd, /*  661 */
128'h87b3cc191ffa7a130ff97793001a0a9b, /*  662 */
128'h179b00f7f71316c166850347c7830144, /*  663 */
128'h02fa0a239a260ff7f7938fd98ff50049, /*  664 */
128'h9dbd8526009ad59b50dc00f482234785, /*  665 */
128'h1ffafa9300099f630005099b86bff0ef, /*  666 */
128'h032a8a239aa60ff979130049591bc40d, /*  667 */
128'h790274a2854e744270e200f482234785, /*  668 */
128'hc783015487b3808261216aa26a4269e2, /*  669 */
128'h0127e9339bc100f979130089591b0347, /*  670 */
128'h099b811ff0ef9dbd0085d59b515cb7e9, /*  671 */
128'h94261fe474130014141bfc0992e30005, /*  672 */
128'h0089591b0109591b0109191b03240a23, /*  673 */
128'h0075d59b515cbf790144822303240aa3, /*  674 */
128'h141bf80996e30005099bfd8ff0ef9dbd, /*  675 */
128'hf0ef85569aa603440a931fc474130024, /*  676 */
128'h179b012569338d71f00006372501da0f, /*  677 */
128'h0087d79b03240a230107d79b94260109, /*  678 */
128'h00fa81230189591b0109579b00fa80a3, /*  679 */
128'hec4ef4267139bf3d4989b745012a81a3, /*  680 */
128'he19d89ae84aae456e852f04af822fc06, /*  681 */
128'h844a04f977634d1c04090a6300c52903, /*  682 */
128'h052a606304f4636324054c9c5afd4a05, /*  683 */
128'hf86347850005041bc43ff0efa8214401, /*  684 */
128'h744270e28522547d00f41d6357fd0887, /*  685 */
128'h4c9c808261216aa26a4269e2790274a2, /*  686 */
128'h85a24409bf554905b7d5faf47ee3894e, /*  687 */
128'h0863fd5507e3c9012501c05ff0ef8526, /*  688 */
128'h85a2167d10000637b76dfb2411e30545, /*  689 */
128'h489c02099063e9052501de9ff0ef8526, /*  690 */
128'h0054c783c89c37fdfae783e3577dc4c0, /*  691 */
128'h852685ce8622bf4900f482a30017e793, /*  692 */
128'h4405f6f50fe34785dd612501dbbff0ef, /*  693 */
128'h2905f822fc0600a55903f04a7139bfad, /*  694 */
128'heb9993c1e456e852ec4ef42603091793, /*  695 */
128'h6aa26a4269e2790274a2744270e24511, /*  696 */
128'h842a8a2e00f97993d7ed495c80826121, /*  697 */
128'h5783e18dc85c61082785480c00099d63, /*  698 */
128'h15230996601cfcf775e30009071b0085, /*  699 */
128'h4783bf5d4501ec1c97ce034787930124, /*  700 */
128'hfc0a9fe30157fab337fd00495a9b0025, /*  701 */
128'h45090097e46347850005049bb27ff0ef, /*  702 */
128'h4d1c6008b761450500f4946357fdbf49, /*  703 */
128'h049be81ff0ef480cf60a0ee306f4e063, /*  704 */
128'h8de357fdfcf48be34785d4bd451d0005, /*  705 */
128'h06136008f5792501dd8ff0ef6008fcf4, /*  706 */
128'h00043a03beeff0ef0345051345812000, /*  707 */
128'h60084a0502aa2823aa5ff0ef855285a6, /*  708 */
128'hd91c415787bb591c00faed6300254783, /*  709 */
128'h0223b7b9c848a83ff0ef85a6c8046008, /*  710 */
128'h5b1c2a856018f1412501d1cff0ef0145, /*  711 */
128'hf04afc06f426f8227139b7e9db1c2785, /*  712 */
128'h02f007130005c783e05ae456e852ec4e, /*  713 */
128'h0ce7906305c0071300e78663842e84aa, /*  714 */
128'h0ae7fc6347fd000447030004a6230405, /*  715 */
128'h47834b2102e0099305c00a9302f00a13, /*  716 */
128'h462d0204b9030d5780630d4782630004, /*  717 */
128'h926300044783b40ff0ef854a02000593, /*  718 */
128'h07930b37906300144783013900230d37, /*  719 */
128'h470d1b378e630024478300f900a302e0, /*  720 */
128'h458100f905a302000793943a09479763, /*  721 */
128'h608848cc100510632501adbff0ef8526, /*  722 */
128'hc7e5000747836c98e96d2501cdaff0ef, /*  723 */
128'h8d6300b78593709cef918ba100b74783, /*  724 */
128'h08e3fff7c683fff74603078507050cb7, /*  725 */
128'h4bdc611cbf75dfdff0ef85264581fed6, /*  726 */
128'hbc232501a85ff0ef85264581b791c55c, /*  727 */
128'h6aa26a4269e2790274a2744270e20004, /*  728 */
128'h8be3bf954709bf1d0405808261216b02, /*  729 */
128'h02400793943a12f6e06302000693f757, /*  730 */
128'h486502000313478145a147014681b7ad, /*  731 */
128'h9101020695130027e793a8dd0505a0d1, /*  732 */
128'h4503c6ed4711a06d268500e50023954a, /*  733 */
128'h00d90023469500d515630e5006930009, /*  734 */
128'h0037f6930ff7f7930027979b01659663, /*  735 */
128'h946346918bb10107671300b694634585, /*  736 */
128'h00e905a39432920116020087671300d7, /*  737 */
128'hc50500b7c783709c4511bf654701bdfd, /*  738 */
128'hcb890207f7930047f713f4e518e34711, /*  739 */
128'hbf154501e80703e30004bc230004a623, /*  740 */
128'h00b5c7836c8cfbf58b91b73d4515fb0d, /*  741 */
128'hc4c8af2ff0ef0007c503609cdbe58bc1, /*  742 */
128'h46a10ff7f7930027979b05659a63bdb9, /*  743 */
128'h47039722930117020017061b873245ad, /*  744 */
128'h0ae3f95704e3f94706e3f4e374e30007, /*  745 */
128'h4c634185551b0187151b02b6f263fd37, /*  746 */
128'h866300054883ed650513000075170005, /*  747 */
128'h7513fbf7051bbd6d4519f11710e30008, /*  748 */
128'h66e30ff57513f9f7051beea87ae30ff5, /*  749 */
128'h7179bdf90ff777130017e7933701eea8, /*  750 */
128'h451184aef406842ae44ee84aec26f022, /*  751 */
128'h6008a0b1c90de199484c49bd0e500913, /*  752 */
128'hc3210007c7036c1ce1292501afaff0ef, /*  753 */
128'h033780630327026303f7f79300b7c783, /*  754 */
128'h70a2450100979a630017b79317e18bfd, /*  755 */
128'h852245818082614569a2694264e27402, /*  756 */
128'h4511b7cd00042a23d9452501c13ff0ef, /*  757 */
128'hf0ef842ae426ec06e82245811101bfe5, /*  758 */
128'hf0ef6008484c0e500493e50d250188ff, /*  759 */
128'h00978d630007c7836c1ced092501a8cf, /*  760 */
128'h4791dd792501bcdff0ef85224585cb99, /*  761 */
128'h8082610564a2644260e2451d00f51363, /*  762 */
128'h049bfa9ff0ef842aec06e426e8221101, /*  763 */
128'h0005049ba42ff0ef6008484ce49d0005, /*  764 */
128'h700c84cff0ef4581020006136c08e085, /*  765 */
128'h00e782234705601c82aff0ef462d6c08, /*  766 */
128'hed6347858082610564a28526644260e2, /*  767 */
128'h694264e2740270a245098082450900b7, /*  768 */
128'hec26f02271794d1c808261456a0269a2, /*  769 */
128'hfcf5fde384ae842ae052e44ee84af406, /*  770 */
128'hf0ef852285a600f4fa634c1c59fd4a05, /*  771 */
128'h0ce3bf754501000914630005091bec8f, /*  772 */
128'h8afff0ef852285a6460103390763fb49, /*  773 */
128'h4783c81c278501378a63481cf15d2501, /*  774 */
128'hbf5d0009049b00f402a30017e7930054, /*  775 */
128'he432e82efc061028ec2a7139b7594505, /*  776 */
128'h8793000077970405426383eff0eff42e, /*  777 */
128'h0023c3196622631800a78733050e7de7, /*  778 */
128'h4501e39897aa00070023c31967620007, /*  779 */
128'hf0ef0828080c460100f618634785cb11, /*  780 */
128'h7175bfe5452d8082612170e22501a0ef, /*  781 */
128'he8daecd6f0d2f4cefca6e122e506f8ca, /*  782 */
128'h84aa89b20005302314050d634925e42e, /*  783 */
128'h10630005091b9d6ff0ef1028002c8a79, /*  784 */
128'h2501b6dff0efe4be1028083c65a21409, /*  785 */
128'h01f9fa1301c9f7934519e011e1196406, /*  786 */
128'he75ff0ef102800f516634791c54dc3e1, /*  787 */
128'hcfcd008a77936406e949008a6a132501, /*  788 */
128'h0ca300f408a302100713046007937aa2, /*  789 */
128'h0b2300e40823000407a30004072300f4, /*  790 */
128'h0e23000405a300e40c2300040ba30004, /*  791 */
128'hc50300040fa300040f2300040ea30004, /*  792 */
128'h0da300040d234785fc9fe0ef85a2000a, /*  793 */
128'h82230005099b00040aa300040a230004, /*  794 */
128'hf0ef030aab03855685ce04098b6300fa, /*  795 */
128'h0135262385da39fd7522e9112501e3ff, /*  796 */
128'h00b44783a895892ac90d250183aff0ef, /*  797 */
128'ha0854921f60981e30049f993e3d98bc5, /*  798 */
128'h0029f993e72d0107f71300b44783f565, /*  799 */
128'h6a13c399008a7793e3ad8b8500098463, /*  800 */
128'h01448523f4800309a78385a279a2020a, /*  801 */
128'hc8c8f33fe0ef0009c503000485a3d09c, /*  802 */
128'ha623c8880069d783dbbfe0ef01c40513, /*  803 */
128'h60aa00f494230134b0230004ae230004, /*  804 */
128'h6b466ae67a0679a6794674e6854a640a, /*  805 */
128'hf8a27119b7d5491db7e5491180826149, /*  806 */
128'hfc5ee0daf0caf4a6fc86e4d6e8d2ecce, /*  807 */
128'h8a2e842a0006a023ec6ef06af466f862, /*  808 */
128'h000998630005099be91fe0ef8ab6e432, /*  809 */
128'h744670e60007899bc39d662200b44783, /*  810 */
128'h7be26b066aa66a4669e6790674a6854e, /*  811 */
128'h00a44783808261096de27d027ca27c42, /*  812 */
128'h40f907bb445c01042903160789638b85, /*  813 */
128'h0b1320000b930006091b00f67463893e, /*  814 */
128'h90631ff777934458fa090ce35c7d0304, /*  815 */
128'hfcb337fd0025478300975c9b60081207, /*  816 */
128'h47854848eb11020c99630ffcfc930197, /*  817 */
128'h4c0cb741498900f405a3478900a7ec63, /*  818 */
128'h05a3478501851763b7e52501bd6ff0ef, /*  819 */
128'h856e4c0c00043d83cc08b7a5498500f4, /*  820 */
128'h0099579b000c861bd5792501b98ff0ef, /*  821 */
128'h002dc683c4b58d3a0007849b00a6073b, /*  822 */
128'h86a6001dc503419684bb00f6f4639fb1, /*  823 */
128'h00a44783f94d250104e050ef85d2863a, /*  824 */
128'h0097fc6341a507bb4c48c3850407f793, /*  825 */
128'h955285da20000613910115020097951b, /*  826 */
128'h9a3e9381020497930094949bc5ffe0ef, /*  827 */
128'h9fa5000aa783c45c9fa54099093b445c, /*  828 */
128'h00a4478304e601634c50b70500faa023, /*  829 */
128'he43a85da4685001dc503c38d0407f793, /*  830 */
128'hf793672200a44783f1392501014050ef, /*  831 */
128'h0017c503863a4685601c00f40523fbf7, /*  832 */
128'h444c01a42e23f11525017c1040ef85da, /*  833 */
128'h0127f46340bb87bb1ff5f5930009049b, /*  834 */
128'he0ef855295a28626030585930007849b, /*  835 */
128'he4cee8caf0a27159b59d499dbf9dbd1f, /*  836 */
128'hec66f062f45ef85aeca6f486fc56e0d2, /*  837 */
128'h8ab689328a2e842a0006a023e46ee86a, /*  838 */
128'h00b44783000997630005099bcb5fe0ef, /*  839 */
128'h694664e6854e740670a60007899bc39d, /*  840 */
128'h6d426ce27c027ba27b427ae26a0669a6, /*  841 */
128'h18078f638b8900a44783808261656da2, /*  842 */
128'h0b1320000b9304f76c630127873b445c, /*  843 */
128'h93631ff777930409046344585c7d0304, /*  844 */
128'hfcb337fd0025478300975c9b60081407, /*  845 */
128'h4581485cef01040c9a630ffcfc930197, /*  846 */
128'h498900f405a3478902e798634705cb91, /*  847 */
128'h445cf3fd0005079bd86ff0ef4c0cb759, /*  848 */
128'h05230207e79300a4478312f76a634818, /*  849 */
128'h498500f405a3478501879763b79500f4, /*  850 */
128'hf79300a44783c85ce311cc1c4858bf99, /*  851 */
128'h85da0017c50346854c50601cc38d0407, /*  852 */
128'hfbf7f79300a44783f96925016b5040ef, /*  853 */
128'h97cff0ef856e4c0c00043d8300f40523, /*  854 */
128'h00a6863b0099579b000c869bd1592501, /*  855 */
128'h74639fb5002dc703c4b58d320007849b, /*  856 */
128'h40ef85d286a6001dc503419704bb00f7, /*  857 */
128'h0297f26341a587bb4c4cf15125016670, /*  858 */
128'h855a95d220000613918115820097959b, /*  859 */
128'h00f40523fbf7f79300a44783a4ffe0ef, /*  860 */
128'h093b445c9a3e9381020497930094949b, /*  861 */
128'h00faa0239fa5000aa783c45c9fa54099, /*  862 */
128'h00e7fa63445c481800c78e634c5cbdd1, /*  863 */
128'hfd0925015cb040ef85da4685001dc503, /*  864 */
128'h87bb1ff575130009049b444801a42e23, /*  865 */
128'h8626030505130007849b0127f46340ab, /*  866 */
128'h0407e79300a447839dbfe0ef952285d2, /*  867 */
128'h1141bd2d499db5f9c81cbf4100f40523, /*  868 */
128'h4783e1752501acffe0ef842ae406e022, /*  869 */
128'h601cc3950407f793cf690207f71300a4, /*  870 */
128'h589040ef030405930017c50346854c50, /*  871 */
128'h00f40523fbf7f79300a44783ed552501, /*  872 */
128'hc703741ce15d2501b77fe0ef6008500c, /*  873 */
128'h0107169b481800e785a30207671300b7, /*  874 */
128'h00d78ea300e78e230086d69b0106d69b, /*  875 */
128'h00e78fa300d78f230187571b0107569b, /*  876 */
128'h169b00e78d2300078ba300078b234858, /*  877 */
128'h0107171b00e78a2327010107571b0107, /*  878 */
128'h0106d69b00e78aa30087571b0107571b, /*  879 */
128'h046007130086d69b00e78c2302100713, /*  880 */
128'h000789a30007892300e78ca300d78da3, /*  881 */
128'h478500f40523fdf7f793600800a44783, /*  882 */
128'h4505ebbfe06f014160a2640200f50223, /*  883 */
128'h842ae406e022114180820141640260a2, /*  884 */
128'h25019cbfe0ef8522e9012501effff0ef, /*  885 */
128'h110180820141640260a200043023e119, /*  886 */
128'h779700054a6395bfe0efec060028e42a, /*  887 */
128'h452d8082610560e2450110a785230000, /*  888 */
128'hf486f0a21028002c4601e42a7159bfe5, /*  889 */
128'h083c65a2ec190005041bb3bfe0efeca6, /*  890 */
128'h6586e41d0005041bcd2ff0efe4be1028, /*  891 */
128'h64e6740670a68522cbd8575277a2e991, /*  892 */
128'hc50374a2cb998bc100b5c78380826165, /*  893 */
128'hfcf41ee34791b7c5c8c897bfe0ef0004, /*  894 */
128'hf8cae122e506e42afca67175bfd94415, /*  895 */
128'h1828002c460184ae00050023f0d2f4ce, /*  896 */
128'h842677e2ecbe081ce5292501acdfe0ef, /*  897 */
128'h040a12634a16c2be02f009934bdc597d, /*  898 */
128'h071b0527470300007717e50567a24501, /*  899 */
128'h186300e780a303a0071300e780230307, /*  900 */
128'h00078023078d00e7812302f007130e94, /*  901 */
128'h808261497a0679a6794674e6640a60aa, /*  902 */
128'h18284581fd452501f89fe0ef18284585, /*  903 */
128'h0007c50365c677e2f5552501e6eff0ef, /*  904 */
128'h2501f63fe0ef18284581c2aa8cdfe0ef, /*  905 */
128'h77e2e1052501e48ff0ef18284581f949, /*  906 */
128'h01450e6325018a7fe0ef0007c50365c6, /*  907 */
128'h67a24711dd612501a9eff0ef18284581, /*  908 */
128'hf5cfe0ef1828100cb7594509f8e516e3, /*  909 */
128'hfc974703973610949301020797134781, /*  910 */
128'h05bbfff7871b04e462630037871beb05, /*  911 */
128'h96b2920166a20206961300e586bb40f4, /*  912 */
128'hb7319c3d01368023fff7c79301271a63, /*  913 */
128'h4603962a1088920102071613b7c12785, /*  914 */
128'h0789bddd4545b7e900c68023377dfc96, /*  915 */
128'h07850007470397369281020416936722, /*  916 */
128'hf8227139b709fe9465e3fee78fa32405, /*  917 */
128'h84ae842ae456e852ec4efc06f04af426, /*  918 */
128'h00b44783000917630005091bfb4fe0ef, /*  919 */
128'h790274a2854a744270e20007891bcf89, /*  920 */
128'h009777634818808261216aa26a4269e2, /*  921 */
128'h00042623445884bae3918b8900a44783, /*  922 */
128'h00a44783c81cfcf778e34818445ce4bd, /*  923 */
128'hf793445c4481bf7d00f405230207e793, /*  924 */
128'h099300a44783fc960ee34c50d3e51ff7, /*  925 */
128'hc50385ce4685601cc3850407f7930304, /*  926 */
128'hf79300a44783ed512501213040ef0017, /*  927 */
128'h0017c50386264685601c00f40523fbf7, /*  928 */
128'h6008bf59cc44ed3525011c1040ef85ce, /*  929 */
128'hfff4869b377dc7290097999b00254783, /*  930 */
128'h413007bb02c6ed630337563b0336d6bb, /*  931 */
128'h4a855a7dd1c19c9dc45c27814c0c8ff9, /*  932 */
128'hd7b51ff4f793c45c9fa5445c0499ea63, /*  933 */
128'h9ca90094d49bcd112501c87fe0ef6008, /*  934 */
128'h47850005059b814ff0efe595484cbfb1, /*  935 */
128'h57fdbded490900f405a3478900f59763, /*  936 */
128'hc84cb5ed490500f405a3478500f59763, /*  937 */
128'he0efcb818b89600800a44783b765cc0c, /*  938 */
128'hc4bfe0efbf6984cee5990005059bfddf, /*  939 */
128'h4f9c601cfabafee3fd4588e30005059b, /*  940 */
128'h013787bb413484bbcc0c445cfaf5fae3, /*  941 */
128'h842ac52de42ef822fc067139b7bdc45c, /*  942 */
128'h67e2e1152501fe6fe0ef0828002c4601, /*  943 */
128'h250197cff0eff01c101ce01c852265a2, /*  944 */
128'h4515e7898bc100b5c783cd996c0ce529, /*  945 */
128'he30fe0ef0007c50367e2a02d00043023, /*  946 */
128'h00f414230067d7838522458167e2c448, /*  947 */
128'h70e2f971fcf50be347912501cbdfe0ef, /*  948 */
128'hfcf501e34791bfdd4525808261217442, /*  949 */
128'h2501dbafe0ef842ae406e0221141b7c1, /*  950 */
128'h717980820141640260a200043023e119, /*  951 */
128'hd98fe0ef892e842af406e84aec26f022, /*  952 */
128'he0ef8522458100091f63e8890005049b, /*  953 */
128'h64e269428526740270a20005049bc5ff, /*  954 */
128'hb32ff0ef852245810224302380826145, /*  955 */
128'h852285ca00042a2302f5136347912501, /*  956 */
128'h47912501f8bfe0ef85224581c68fe0ef, /*  957 */
128'hbf6584aad16dbf7d00042a2300f51663, /*  958 */
128'hf0a21028002c460184aee42aeca67159, /*  959 */
128'h083c65a2e00d0005041bedafe0eff486, /*  960 */
128'h6786e8010005041b872ff0efe4be1028, /*  961 */
128'h70a68522c10fe0ef102885a6c489cf81, /*  962 */
128'hf0a27159bfcd44198082616564e67406, /*  963 */
128'he0d28522002c46018b2ee42af85a8432, /*  964 */
128'hec66f062f45efc56e4cee8caeca6f486, /*  965 */
128'h2c836000000a1c6300050a1be7cfe0ef, /*  966 */
128'h00fb202302f76263ffec871b481c0184, /*  967 */
128'h7ae26a0669a6694664e68552740670a6, /*  968 */
128'h00044b83808261656ce27c027ba27b42, /*  969 */
128'h85ca4a8559fd4481490902fb9f634785, /*  970 */
128'h09550863093508632501a55fe0ef8522, /*  971 */
128'h00544783fef963e329054c1c2485e111, /*  972 */
128'hb74d009b202300f402a30017e793c804, /*  973 */
128'h1afd4c0944814981490110000ab7504c, /*  974 */
128'h2501d10fe0ef0015899b852200099e63, /*  975 */
128'h038b9163200009930344091385cee921, /*  976 */
128'he3918fd90087979b0009470300194783, /*  977 */
128'h854ab745fc0c94e33cfd39f909092485, /*  978 */
128'he1116582015575332501abcfe0efe02e, /*  979 */
128'hbfbd4a09b7494a05b7c539f109112485, /*  980 */
128'h842ae04aec06e426e8221101bfad8a2a, /*  981 */
128'hcb9100b44783e4910005049bbc4fe0ef, /*  982 */
128'h610564a269028526644260e20007849b, /*  983 */
128'h48144458cf390027f71300a447838082, /*  984 */
128'h600800f40523c8180207e793fed772e3, /*  985 */
128'hc53900042a232501a58ff0ef484cef01, /*  986 */
128'h091b94dfe0ef4c0cbf7d84aa00a405a3, /*  987 */
128'h06374c0cb7dd450502f9146357fd0005, /*  988 */
128'h85ca6008f9792501b37fe0ef167d1000, /*  989 */
128'h45094785b769449db7e12501a1cff0ef, /*  990 */
128'h00a44783fcf96ae34d1c6008fcf900e3, /*  991 */
128'h0017c50346854c50601cdba50407f793, /*  992 */
128'h00a44783f55d25015f0040ef03040593, /*  993 */
128'h4605e42a7175b7b100f40523fbf7f793, /*  994 */
128'hca0fe0eff8cafca6e122e5061008002c, /*  995 */
128'he3bfe0efe0be1008081c65a2e9052501, /*  996 */
128'h0207f79300b7c78345196786e1052501, /*  997 */
128'hcb810014f79300b5c483c59975e2eb89, /*  998 */
128'h790280826149794674e6640a60aa451d, /*  999 */
128'h88c1cc0d0005041bad8fe0ef00094503, /* 1000 */
128'h100c02800613fc878de301492783c89d, /* 1001 */
128'h951fe0efcaa200a8458996cfe0ef00a8, /* 1002 */
128'hd94d2501836ff0ef00a84581f1612501, /* 1003 */
128'hf15525019f5fe0ef1008faf518e34791, /* 1004 */
128'h85a27502bf612501f20fe0ef7502e411, /* 1005 */
128'h4605e42a7171b769d575250191cff0ef, /* 1006 */
128'he152e54ee94aed26f506f1221028002c, /* 1007 */
128'hbd0fe0efe8eaece6f0e2f4def8dafcd6, /* 1008 */
128'he4be1028083c65a21c0414630005041b, /* 1009 */
128'h176347911c0409630005041bd67fe0ef, /* 1010 */
128'h9f630207f79300b7c783441967a61af4, /* 1011 */
128'h02630005091bb45fe0ef458175221807, /* 1012 */
128'h0b63440557fd16f90f63440947851809, /* 1013 */
128'h160414630005041ba98fe0ef752216f9, /* 1014 */
128'h0a13f6efe0ef85220109549b85ca7422, /* 1015 */
128'he0ef855200050c1b4581200006130344, /* 1016 */
128'h248188cfe0ef855202000593462d898f, /* 1017 */
128'h0fa30104949b0109199b0ff4fb1347c1, /* 1018 */
128'h0b930104d49b021007930109d99b02f4, /* 1019 */
128'hd99b046007930ff97a9304f4062302e0, /* 1020 */
128'h0a230200061304f406a30084d49b0089, /* 1021 */
128'h07a305540723040405a3040405230374, /* 1022 */
128'h0544051385d2049404a3056404230534, /* 1023 */
128'h00074603468d05740aa3772280efe0ef, /* 1024 */
128'h0723478100f69363571400d6166357d2, /* 1025 */
128'h06f4042327810107d79b0107969b06f4, /* 1026 */
128'h0086d69b0107d79b0106d69b0107979b, /* 1027 */
128'h00274b8306f404a306d407a30087d79b, /* 1028 */
128'h0005041bf59fe0ef1028040b99634c85, /* 1029 */
128'h0210071300e785a3752247416786e835, /* 1030 */
128'h00078ba300078b230460071300e78c23, /* 1031 */
128'h01678a2301378da301578d2300e78ca3, /* 1032 */
128'h041bd5afe0ef00f50223478500978aa3, /* 1033 */
128'h022303852823001c0d1b7522a82d0005, /* 1034 */
128'h20000613ec090005041b8dcfe0ef0195, /* 1035 */
128'h8c6a0ffbfb93f61fd0ef3bfd85524581, /* 1036 */
128'h70aa8522f25fe0ef85ca7522441db749, /* 1037 */
128'h7ba67b467ae66a0a69aa694a64ea740a, /* 1038 */
128'h7159b7c544218082614d6d466ce67c06, /* 1039 */
128'h10284605002c843284aee42aeca6f0a2, /* 1040 */
128'h1028083c65a2e13125019cafe0eff486, /* 1041 */
128'hc783451967a6e9152501b65fe0efe4be, /* 1042 */
128'h00b74783c30d6706e39d0207f79300b7, /* 1043 */
128'h008705a38c3d027474138c658cbd7522, /* 1044 */
128'h740670a62501c9efe0ef00f502234785, /* 1045 */
128'h002c4605e02ee42a71718082616564e6, /* 1046 */
128'h0005079b964fe0efed26f122f5060088, /* 1047 */
128'hf0be083cf4be008865a2678612079663, /* 1048 */
128'hc703778610079a630005079baf7fe0ef, /* 1049 */
128'h479165e61007126302077713479900b7, /* 1050 */
128'h0613e55fd0ef102805ad46550e058e63, /* 1051 */
128'hf05fd0ef850ae49fd0ef10a8008c0280, /* 1052 */
128'h079baadfe0ef10a865820c054d6347ad, /* 1053 */
128'hdc5fe0ef10a80ce793634711cbf90005, /* 1054 */
128'h851302a10593464d648aefc50005079b, /* 1055 */
128'h0207e793640602814783e0dfd0ef00d4, /* 1056 */
128'h8bc100b4c78300f40223478500f485a3, /* 1057 */
128'h85a60004450306f7086357d64736cbbd, /* 1058 */
128'h059bcaefe0ef85220005059bf2dfd0ef, /* 1059 */
128'h0005079bfc3fd0ef8522c5a547890005, /* 1060 */
128'h02f69d630557468302e007936706efb1, /* 1061 */
128'h27810107d79b06f707230107969b57d6, /* 1062 */
128'h0087d79b0107d79b0107979b06f70423, /* 1063 */
128'h07a3478506f704a30086d69b0106d69b, /* 1064 */
128'h0005079be24fe0ef008800f7022306d7, /* 1065 */
128'h740a70aa0005079bb50fe0ef6506e791, /* 1066 */
128'he8a2711dbfcd47a18082614d853e64ea, /* 1067 */
128'h810fe0efec861028002c4605842ee42a, /* 1068 */
128'h9abfe0efe4be1028083c65a2e9292501, /* 1069 */
128'h0207f79300b7c783451967a6e1292501, /* 1070 */
128'h00e78b23752200645703cb856786eb95, /* 1071 */
128'h00e78c230044570300e78ba30087571b, /* 1072 */
128'he0ef00f50223478500e78ca30087571b, /* 1073 */
128'he4a6711d80826125644660e62501ad6f, /* 1074 */
128'he8a208284601002c893284aee42ae0ca, /* 1075 */
128'h4581c4b9e0510005041bf9bfd0efec86, /* 1076 */
128'h08284585e5592501ca8fe0efd2020828, /* 1077 */
128'hd0ef8526462d75c2e93d2501b8ffe0ef, /* 1078 */
128'h000700230200061346ad00b48713ca1f, /* 1079 */
128'h97a6938117820007869bfff6879bce89, /* 1080 */
128'h656202090a63fec783e3177d0007c783, /* 1081 */
128'h470d6562e0150005041be69fd0ef510c, /* 1082 */
128'h0270079300e684630005468304300793, /* 1083 */
128'h852200a92023c29fd0ef953e03478793, /* 1084 */
128'h1563479180826125690664a6644660e6, /* 1085 */
128'he42a711db7d5842abf550004802300f5, /* 1086 */
128'h041bee3fd0efec86e8a21028002c4605, /* 1087 */
128'h02061793460100010c2366a2ec550005, /* 1088 */
128'hea2902000593eba10007c78397b69381, /* 1089 */
128'he8410005041bbd6fe0efda0210284581, /* 1090 */
128'h01814783e1792501abbfe0ef10284585, /* 1091 */
128'h07136786bc7fd0ef082c462dc3dd6506, /* 1092 */
128'h8ba300078b230460071300e78c230210, /* 1093 */
128'hbf45863eb74d2605a06100e78ca30007, /* 1094 */
128'h000747039736930102079713fff6079b, /* 1095 */
128'h07f00e9343658e2e4781082cfeb706e3, /* 1096 */
128'h91411542f9f7051b27850006c70348b1, /* 1097 */
128'h05130000651793411742370100a36c63, /* 1098 */
128'h8522441900eef863a82100070f1b8ee5, /* 1099 */
128'h48030505bfcdf36d80826125644660e6, /* 1100 */
128'h00fe06b3b7cdffe81be3060805630005, /* 1101 */
128'h752200f500235795a885078500c68023, /* 1102 */
128'hb7c10005041b8fefe0ef00f502234785, /* 1103 */
128'he0ef1028dbd50181478302f51b634791, /* 1104 */
128'h4581020006136506f4450005041ba55f, /* 1105 */
128'h6786ae5fd0ef082c462d6506b07fd0ef, /* 1106 */
128'hf91780e3b751842abf1900e785a34721, /* 1107 */
128'h93811782f4c7e5e30585068500e58023, /* 1108 */
128'h4703f8d771e30007869b020006134729, /* 1109 */
128'h05052e83bf89eaf71de30e5007930181, /* 1110 */
128'hec22110105c528830585230305452e03, /* 1111 */
128'h87f2869a8646040502938f2ae44ae826, /* 1112 */
128'h8dfd00c6c5b306ef8f9300004f978876, /* 1113 */
128'h008fa403000f2583000fa38300b64733, /* 1114 */
128'h004f2703ff4fa3839db9007585bb0fc1, /* 1115 */
128'h0105e8330198581b0078159b0105883b, /* 1116 */
128'h8e6d00f6c6339f3100f805bb0077073b, /* 1117 */
128'h0146561b00c6171b9e39008f23838e35, /* 1118 */
128'hc6b300d383bb00c5873b008383bb8e59, /* 1119 */
128'hd39b007686bb8ebd00cf24038ef900b7, /* 1120 */
128'hffcfa4039fa100d3e6b30116969b00f6, /* 1121 */
128'h9fa1007777338f2d0007061b00d703bb, /* 1122 */
128'h0f418f5d0167171b00a7579b9f3d8f2d, /* 1123 */
128'hf45f17e300e387bb0003869b0005881b, /* 1124 */
128'hfe8f8f9300004f970b05859300004597, /* 1125 */
128'h00cf7f3300d7cf330b02829300004297, /* 1126 */
128'h0025c4030015c383000faf0301e6c733, /* 1127 */
128'h972a070a93aa038a0005c70300ef0f3b, /* 1128 */
128'h083b004fa70300ef0f3b942a040a4318, /* 1129 */
128'h0003a70301b8581b9e3900581f1b010f, /* 1130 */
128'h8e7501e7c6339f3100f80f3b010f6833, /* 1131 */
128'h0176561b0096139b008fa7039e398e3d, /* 1132 */
128'h05919f3500cf03bb00c3e63340189eb9, /* 1133 */
128'h0fc101e6c6b3fff5c4838efd007f46b3, /* 1134 */
128'h9fb900e6941b94aa048affcfa7039eb9, /* 1135 */
128'hc7339fb900d3843b8ec140980126d69b, /* 1136 */
128'h00c7579b9f3d0077473301e777330083, /* 1137 */
128'h069b0003861b000f081b8f5d0147171b, /* 1138 */
128'h0f1300004f17f25599e300e407bb0004, /* 1139 */
128'h010fc403f3c38393000043978ffafc6f, /* 1140 */
128'h00c2c4b3942a040a00d7c2b30003a703, /* 1141 */
128'h048a0043a4039f21011fc4839f254000, /* 1142 */
128'h171b012fc4830107083b40809e2194aa, /* 1143 */
128'h0083a4039e210107683301c8581b0048, /* 1144 */
128'h863b9ea194aa00e2c2b3048a00f8073b, /* 1145 */
128'h0156561b013fc90300b6129b408000c2, /* 1146 */
128'hffc3a4839c3500c702bb03c100c2e633, /* 1147 */
128'h941b992a9ea1090a0056c6b300e7c6b3, /* 1148 */
128'h843b8ec1000924830106d69b9fa50106, /* 1149 */
128'h9f3d8f219fa5005747330007081b00d2, /* 1150 */
128'h0002861b0f918f5d0177171b0097579b, /* 1151 */
128'h00004297f5f592e300e407bb0004069b, /* 1152 */
128'ha70300d745b38f5dfff64713eb428293, /* 1153 */
128'h020f45839f2d022f4403021f43830002, /* 1154 */
128'h9f2d942a040a418c95aa058a93aa038a, /* 1155 */
128'ha5839e2d0068171b0107083b0042a583, /* 1156 */
128'h9db100f8073b0107683301a8581b0003, /* 1157 */
128'h139b0082a5839e2d8e3d8e59fff6c613, /* 1158 */
128'h03bb00c3e633400c9ead0166561b00a6, /* 1159 */
128'h0075e5b3fff7c593023f44839ead00c7, /* 1160 */
128'h00f5969b048a9db5ffc2a4038db902c1, /* 1161 */
128'h00b385bb40809fa18dd50115d59b94aa, /* 1162 */
128'h007747339fa18f4dfff747130007081b, /* 1163 */
128'h861b0f118f5d0157171b00b7579b9f3d, /* 1164 */
128'h6462f3ef9de300e587bb0005869b0003, /* 1165 */
128'h00c8863b00d306bb00fe07bb010e883b, /* 1166 */
128'h6105692264c2cd70cd34c97c05052823, /* 1167 */
128'he85af44ef84afc26e0a2715d653c8082, /* 1168 */
128'h84aa97b203f7f413ec56f052e486e45e, /* 1169 */
128'h07bb04000b9304000b13e53c893289ae, /* 1170 */
128'h0a1b00f974639381178200078a1b408b, /* 1171 */
128'h0084853385ce020ada93020a1a930009, /* 1172 */
128'h99d64159093348d020ef0144043b8656, /* 1173 */
128'h60a6b7c997824401852660bc01741763, /* 1174 */
128'h6ba26b426ae27a0279a2794274e26406, /* 1175 */
128'h842a03f7f793f0227179653c80826161, /* 1176 */
128'hf800071300178513e84af406e44eec26, /* 1177 */
128'h40a9863b449d0400099300e7802397a2, /* 1178 */
128'h3d5020ef95224581920116020006091b, /* 1179 */
128'h97828522603cfc1c078e643c0124f563, /* 1180 */
128'h69a2694264e2740270a2fd24fde34501, /* 1181 */
128'h3423639cc34787930000679780826145, /* 1182 */
128'hed3c639cc2c7879300006797e93c0405, /* 1183 */
128'h059311018082e13cb6c7879300000797, /* 1184 */
128'h669747013cb020efec06850a46410505, /* 1185 */
128'h45413825859300005597e72686930000, /* 1186 */
128'h0047d613070506890007c78300e107b3, /* 1187 */
128'h8f230007c78397ae000646038bbd962e, /* 1188 */
128'h0000651760e2fca71de3fef68fa3fec6, /* 1189 */
128'h0808842ae122717580826105e3450513, /* 1190 */
128'hf0ef080885a26622f71ff0efe42ee506, /* 1191 */
128'h60aaf83ff0ef0808f01ff0ef0808e85f, /* 1192 */
128'h00d70d63711c46a1595880826149640a, /* 1193 */
128'h80824501cf980200071300d717634691, /* 1194 */
128'he426e82211018082556dbfe50007ac23, /* 1195 */
128'h469702f5026384ae842a200007b7ec06, /* 1196 */
128'h85930000559708800613c62686930000, /* 1197 */
128'hfc2409f030ef2f650513000055172e65, /* 1198 */
128'h6100e82211018082610564a2644260e2, /* 1199 */
128'h469702f4026384ae200007b7ec06e426, /* 1200 */
128'h85930000559702f00613c3a686930000, /* 1201 */
128'he00405f030ef2b650513000055172a65, /* 1202 */
128'h6100e82211018082610564a2644260e2, /* 1203 */
128'h469702f4026384ae200007b7ec06e426, /* 1204 */
128'h85930000559703600613c0a686930000, /* 1205 */
128'he40401f030ef27650513000055172665, /* 1206 */
128'h6104e42611018082610564a2644260e2, /* 1207 */
128'h669702f48263842e200007b7ec06e822, /* 1208 */
128'h85930000559703e00613bb2686930000, /* 1209 */
128'h14027de030ef23650513000055172265, /* 1210 */
128'h11018082610564a2644260e2e8809001, /* 1211 */
128'h8263842e200007b7ec06e8226104e426, /* 1212 */
128'h559704500613b66686930000669702f4, /* 1213 */
128'h30ef1f250513000055171e2585930000, /* 1214 */
128'h610564a2644260e2ec809001140279a0, /* 1215 */
128'h200007b7ec06e4266100e82211018082, /* 1216 */
128'h0613b52686930000469702f4026384ae, /* 1217 */
128'h05130000551719e585930000559704c0, /* 1218 */
128'h610564a2644260e2f004756030ef1ae5, /* 1219 */
128'h200007b7ec06e4266100e82211018082, /* 1220 */
128'h0613b22686930000469702f4026384ae, /* 1221 */
128'h05130000551715e58593000055970530, /* 1222 */
128'h610564a2644260e2f404716030ef16e5, /* 1223 */
128'hf04af426f82200053983ec4e71398082, /* 1224 */
128'h02f984638436893284ae200007b7fc06, /* 1225 */
128'h0000559705a00613ae86869300004697, /* 1226 */
128'h30efe43a124505130000551711458593, /* 1227 */
128'h0029191b8b0589890014159b67226ca0, /* 1228 */
128'h88a10125e5b30034949b8dd900497913, /* 1229 */
128'h69e2790274a202b9b8238dc5744270e2, /* 1230 */
128'h4605468147057100e022114180826121, /* 1231 */
128'hf0ef45818522f7dff0efe40645818522, /* 1232 */
128'hf67ff0ef45814605468547058522f35f, /* 1233 */
128'h01414501640260a2d97ff0ef45816008, /* 1234 */
128'h3c23460546814705e022e40611418082, /* 1235 */
128'h8522f39ff0ef842a4581040530230205, /* 1236 */
128'h46054685470545818522ef1ff0ef4581, /* 1237 */
128'hf06f0141458160a264026008f23ff0ef, /* 1238 */
128'h200007b7ec06e8226104e4261101d4df, /* 1239 */
128'h0613a12686930000469702f48263842e, /* 1240 */
128'h05130000551702e58593000055970610, /* 1241 */
128'h644260e2fc80904114425e6030ef03e5, /* 1242 */
128'hec06e8226104e42611018082610564a2, /* 1243 */
128'h86930000469702f48263842e200007b7, /* 1244 */
128'h5517fea5859300005597068006139de6, /* 1245 */
128'h8c7d17fd67855a2030efffa505130000, /* 1246 */
128'he82211018082610564a2644260e2e0a0, /* 1247 */
128'h02f4026384ae200007b7ec06e4266100, /* 1248 */
128'h0000559706f006139a86869300004697, /* 1249 */
128'h55c030effb45051300005517fa458593, /* 1250 */
128'he04a11018082610564a2644260e2e424, /* 1251 */
128'h842a200007b7ec06e426e82200053903, /* 1252 */
128'h0613972686930000469702f9026384ae, /* 1253 */
128'h051300005517f5e58593000055970760, /* 1254 */
128'h644260e2c84404993c23516030eff6e5, /* 1255 */
128'heca67100f0a2715980826105690264a2, /* 1256 */
128'hf062f45ef85afc56e0d2e4cef486e8ca, /* 1257 */
128'he03084b2892e0005d783020408a3ec66, /* 1258 */
128'h9c636d6020ef00c9051345814611d01c, /* 1259 */
128'h07b700043983bf5ff0ef458560080e04, /* 1260 */
128'h44810049278316f99a6304043a032000, /* 1261 */
128'h4c1c4485e391448d8b89c7090017f713, /* 1262 */
128'h8b85008a2783000a09638cdd03243c23, /* 1263 */
128'h45814605468147050144e49316078663, /* 1264 */
128'h2583be1ff0ef85224581d71ff0ef8522, /* 1265 */
128'hc4fff0ef8ecc0c1300004c1785220089, /* 1266 */
128'hf0efe8aa0a1300005a17852200095583, /* 1267 */
128'hf0ef85224581cbdff0ef852285a6c81f, /* 1268 */
128'hd27ff0ef85224581460546854705cf5f, /* 1269 */
128'h4585e93ff0ef852224058593000f45b7, /* 1270 */
128'h009899b785220d89b583cd1ff0ef8522, /* 1271 */
128'h5a9768198993eb7ff0ef25810015e593, /* 1272 */
128'h64e6740670a6efe9485ce4aa8a930000, /* 1273 */
128'h6ce27c027ba27b427ae26a0669a66946, /* 1274 */
128'hdb7ff0efe024852244cc808261654501, /* 1275 */
128'hee079be38b85449cdf3ff0ef8522488c, /* 1276 */
128'h458163900107e683654100043883603c, /* 1277 */
128'h6e89f005051300ff0e37431147014781, /* 1278 */
128'h183b070500371f1b00064803ec0689e3, /* 1279 */
128'h0067036316fd060527810107e7b301e8, /* 1280 */
128'h981b010767330187971b0187d81bf2e5, /* 1281 */
128'h8fe9010767330087d79b01c878330087, /* 1282 */
128'h9746938183751782170200be873b8fd9, /* 1283 */
128'h869300003697b765470147812585e31c, /* 1284 */
128'h5517d6a58593000055971490061378e6, /* 1285 */
128'h00c4e493bd85322030efd7a505130000, /* 1286 */
128'h3597000b1d633b7d20000bb78b4ebd61, /* 1287 */
128'h00efd6a5051300005517772585930000, /* 1288 */
128'h061386e20179096300043903b7117020, /* 1289 */
128'h485c070934832e2030ef855685d20f20, /* 1290 */
128'h37830209370312048e6324818cfd4c81, /* 1291 */
128'hcc5cf9200793c7817c1c00f76f630c89, /* 1292 */
128'hb27ff0ef85224581b6fff0ef85224581, /* 1293 */
128'hff397913852201442903c3950044f793, /* 1294 */
128'h0000551785cad47ff0ef85ca00896913, /* 1295 */
128'h2903c3950084f79368c000efd0c50513, /* 1296 */
128'hf0ef85ca00496913ff39791385220144, /* 1297 */
128'h664000efd0c505130000551785cad1ff, /* 1298 */
128'h8c630384390300043c83cfb50014f793, /* 1299 */
128'h85d209c006136de6869300003697017c, /* 1300 */
128'h3c2300492783cba97c1c236030ef8556, /* 1301 */
128'h018c871308e69f630037f693470d0204, /* 1302 */
128'hff87051363104591480d468100c90793, /* 1303 */
128'h8361ff87370301068763c3900086161b, /* 1304 */
128'h603cfeb690e30791872a2685c3988f51, /* 1305 */
128'hc85c9bf9485cc85c0027e793485ccbb5, /* 1306 */
128'h01748c63040439036004cc9d4c858889, /* 1307 */
128'h855685d20ca006136786869300003697, /* 1308 */
128'h0089278300090963040430231b8030ef, /* 1309 */
128'h9bf54c85485cb4dff0ef8522ef8d8b85, /* 1310 */
128'h4505d80c8ee3c47ff0ef8522484cc85c, /* 1311 */
128'h2623000cb783dbd98b85bd955e1020ef, /* 1312 */
128'h97a667a1bf41b1dff0ef8522b77100f9, /* 1313 */
128'h8913fa978de394be00093c8301096483, /* 1314 */
128'h3a6020efe43e002c46218566639c0087, /* 1315 */
128'h0513717908b041635535b7dd87ca0ca1, /* 1316 */
128'h892e84b2e44ef406e84aec26f0220480, /* 1317 */
128'h0000351785a2cc1d5551842a0a8030ef, /* 1318 */
128'h5517862285aa89aa791010ef5e450513, /* 1319 */
128'h07b702098b6350a000efbda505130000, /* 1320 */
128'hcb990024f793f40401242423e01c2000, /* 1321 */
128'h69a2694264e2740270a24501c45c4789, /* 1322 */
128'hb7e5c45c4785d4fd4501888580826145, /* 1323 */
128'h458146098082bff9557d090030ef8522, /* 1324 */
128'h953e050e200007b7f73ff06f20000537, /* 1325 */
128'he4066380e0221141711c808225016108, /* 1326 */
128'h580686930000369702f40263200007b7, /* 1327 */
128'h00005517abc585930000559734c00613, /* 1328 */
128'h557de3914505703c074030efacc50513, /* 1329 */
128'h4501842ae822110180820141640260a2, /* 1330 */
128'h60e26622644285a24df010efe42eec06, /* 1331 */
128'hf4062000051371797a00006f61054685, /* 1332 */
128'h84aa7af020efe052e44ee84aec26f022, /* 1333 */
128'h0001b5030b6030efb305051300005517, /* 1334 */
128'h212010ef842a49d010ef4501457010ef, /* 1335 */
128'h404000ef638cb165051300005517681c, /* 1336 */
128'h3f4000efb14505130000551706f44583, /* 1337 */
128'h15c20085d59bb1e5051300005517546c, /* 1338 */
128'h0000551706c44583583c3de000ef91c1, /* 1339 */
128'h0187d61b0107d69b0087d71bb1450513, /* 1340 */
128'h00ef26010ff6f6930ff7f7930ff77713, /* 1341 */
128'h3a4000efb0450513000055175c0c3b20, /* 1342 */
128'h00005597c789a8e5859300005597545c, /* 1343 */
128'h384000efaf45051300005517a7c58593, /* 1344 */
128'h55977448006030efb005051300005517, /* 1345 */
128'h584c19c42783db9fb0ef08a585930000, /* 1346 */
128'h061300005617e789a586061300005617, /* 1347 */
128'h8526346000efade5051300005517de66, /* 1348 */
128'h0a1300005a174481ed5ff0ef84264581, /* 1349 */
128'hf79320000913ade9899300005997adea, /* 1350 */
128'h00044583318000ef855285a6e78901f4, /* 1351 */
128'h0405306000ef819100f5f6132485854e, /* 1352 */
128'h2f4000ef0145051300005517fd249fe3, /* 1353 */
128'h614545016a0269a2694264e2740270a2, /* 1354 */
128'hb7033bb0206face50513000055178082, /* 1355 */
128'h278540f707b30003b6830083b7830103, /* 1356 */
128'h00f3b8230017079300d7fe6393811782, /* 1357 */
128'h80820007802345050103b78300a70023, /* 1358 */
128'h020596130103b7830083b70380824501, /* 1359 */
128'hf5638e9dfff706930003b7038f999201, /* 1360 */
128'hb70340a786bb87aa9d9dfff7059b00c6, /* 1361 */
128'h06938082852e0007002300b6e6630103, /* 1362 */
128'h00d7002307850007c68300d3b8230017, /* 1363 */
128'h488540a0053be681000556634881bfe9, /* 1364 */
128'h4e250ff6f81304100693c21906100693, /* 1365 */
128'h0ff3751302b6733b0005061b385986ba, /* 1366 */
128'h0ff5751302b6563b0305051b046e6763, /* 1367 */
128'h051340e685bbfe718532fea68fa30685, /* 1368 */
128'h802302d007930008876302f5e9630300, /* 1369 */
128'h000680230015559b40e6853b068500f6, /* 1370 */
128'h053b808200b61b63fff5081b86ba2581, /* 1371 */
128'h07bbb7d92585fea68fa30685bf5d00a8, /* 1372 */
128'h0006c8830007c30397ba9381178240c8, /* 1373 */
128'h7119b7f1068501178023006680232605, /* 1374 */
128'he4d6e8d2eccef4a6f8a2597d011cf0ca, /* 1375 */
128'hf82af02ef42afc3e843684b2e0dafc86, /* 1376 */
128'h0209591303000a9306c00a1302500993, /* 1377 */
128'h0017079bc52d8f1d0004c50377a27742, /* 1378 */
128'h04850135086304d7ff63938117827682, /* 1379 */
128'h0f630014c503bfe1e7bff0ef02010393, /* 1380 */
128'hcb9d0004c78303551063478104890545, /* 1381 */
128'h478100f6f36346a50ff7f793fd07879b, /* 1382 */
128'heb6306d50f630640069304890014c503, /* 1383 */
128'h09630630079304d50f630580069302a6, /* 1384 */
128'h6a4669e6790674a6744670e6f55d08f5, /* 1385 */
128'h0024c503808261090007051b6b066aa6, /* 1386 */
128'h00a76c6306e50e6307300713b74d048d, /* 1387 */
128'h4685003800840b13f6e51ee307000713, /* 1388 */
128'h0780071302e5006307500713a00d4601, /* 1389 */
128'h4685003800840b13fa850613f6e510e3, /* 1390 */
128'h00840b13f8b50693a81145c100163613, /* 1391 */
128'he37ff0ef400845a946010016b6930038, /* 1392 */
128'ha809ddbff0ef0028020103930005059b, /* 1393 */
128'hd93ff0ef00840b130201039300044503, /* 1394 */
128'h852201247433600000840b13b5fd845a, /* 1395 */
128'hb7f18522020103930005059b4db010ef, /* 1396 */
128'he4c6e0c2fc3ef83aec061034f436715d, /* 1397 */
128'hf032715d8082616160e2e8dff0efe436, /* 1398 */
128'hfc3ef83aec06100005931014862ef436, /* 1399 */
128'h8082616160e2e69ff0efe436e4c6e0c2, /* 1400 */
128'h100005931234862afe36fa32f62e710d, /* 1401 */
128'he436eec6eac2e6bee2baea22ee060808, /* 1402 */
128'h60f285220bd020ef0808842ae3fff0ef, /* 1403 */
128'h03630087b303679c691c808261356452, /* 1404 */
128'h979304b7ee63479d8082450183020003, /* 1405 */
128'h439c97ba83f90ce70713000037170205, /* 1406 */
128'h2483795c878297bae426e822ec061101, /* 1407 */
128'h9381020497930c5010ef7540f55c08c5, /* 1408 */
128'h61054501e91c64a2644260e202f457b3, /* 1409 */
128'h058e05e135f1bfd9617cbfe97d5c8082, /* 1410 */
128'h11418082557d8082557db7e9659c95aa, /* 1411 */
128'h681c00055e63ff5ff0ef842ae406e022, /* 1412 */
128'h60a264028522000307630207b303679c, /* 1413 */
128'h557d80820141640260a2450183020141, /* 1414 */
128'h879300003797150200a7eb6347ad8082, /* 1415 */
128'h05130000451780826108953e81750567, /* 1416 */
128'h715d83020007b303679c691c80826fe5, /* 1417 */
128'h078517824785d23e47d502f1102347a1, /* 1418 */
128'hd402e486100c200007930030e83ee42e, /* 1419 */
128'h07374d148082616160a6fd3ff0efcc3e, /* 1420 */
128'h2381308345018082450100e6fe634004, /* 1421 */
128'h01138082240101132281348323013403, /* 1422 */
128'h342385a2980101f1041322813823dc01, /* 1423 */
128'hf579f95ff0ef1a05348322113c232291, /* 1424 */
128'h0dd4c70302f71c630a0447830a04c703, /* 1425 */
128'h0c0447830c04c70302f716630dd44783, /* 1426 */
128'h00f71a630e0447830e04c70302f71063, /* 1427 */
128'hd55156f010ef0d4485130d4405934611, /* 1428 */
128'h3e800513842af0227179b761fb600513, /* 1429 */
128'h00011023858a4601852267e020eff406, /* 1430 */
128'h7d000513e509842af21ff0efc202c402, /* 1431 */
128'h717980826145740270a28522660020ef, /* 1432 */
128'hc402c23ef406f022478500f110234785, /* 1433 */
128'h87934ad4008007b745386914c195842a, /* 1434 */
128'h400006b78f75600006b78ff58ff9f807, /* 1435 */
128'hec9ff0ef8522858a4601c43e8fd98f55, /* 1436 */
128'h711d80826145740270a2c43c47b2e119, /* 1437 */
128'he0ca07c55783c23e47d500f1102347b5, /* 1438 */
128'h6a056989fdf949370107979bf852fc4e, /* 1439 */
128'h4495c43e842e8aaaec86f456e4a6e8a2, /* 1440 */
128'h858a4601e00a0a13e009899308090913, /* 1441 */
128'hc7891005f79345b2ed0de73ff0ef8556, /* 1442 */
128'h4517c78d0125f7b3054793630135f7b3, /* 1443 */
128'h60e6fba00513d4bff0ef55a505130000, /* 1444 */
128'h808261257aa27a4279e2690664a66446, /* 1445 */
128'h00f057630014079b347dfe04c6e334fd, /* 1446 */
128'hfc8049e34501b75556c020ef3e800513, /* 1447 */
128'hf9200513d09ff0ef5305051300004517, /* 1448 */
128'h00f1102347c17139e7a919c52783bf7d, /* 1449 */
128'h842af426fc06f822858a460147d5c42e, /* 1450 */
128'hcb918b891b842783c11dde3ff0efc23e, /* 1451 */
128'h34fdc901dcdff0ef8522858a46014495, /* 1452 */
128'hbfd545018082612174a2744270e2f8ed, /* 1453 */
128'h4785e8a2ec86e0cae4a6711d80824501, /* 1454 */
128'h102302c9270347c906d7f66384b6892a, /* 1455 */
128'he42e4755d432cf3108c92783260102f1, /* 1456 */
128'hc83eca26d23a854a100c47850030cc3e, /* 1457 */
128'h47b10497f0634785e529842ad75ff0ef, /* 1458 */
128'hd23ed402854a100c47f5460102f11023, /* 1459 */
128'hf0ef48a5051300004517c11dd55ff0ef, /* 1460 */
128'h80826125690664a6644660e68522c43f, /* 1461 */
128'hb7d50004841bb74d02f6063bbf6147c5, /* 1462 */
128'hec4ef04af426f822fc067139b7c54401, /* 1463 */
128'h8ab684b28a2e4148842ace05e456e852, /* 1464 */
128'ha0ef852200b44583c11d892a482010ef, /* 1465 */
128'h00b67a63014485b3681000054d638d7f, /* 1466 */
128'ha0894481bd9ff0ef4405051300004517, /* 1467 */
128'h378389a6f96decdff0ef854a08c92583, /* 1468 */
128'h865286a2844e0089f3630207e4030109, /* 1469 */
128'h08c96783fc851ae3f01ff0ef854a85d6, /* 1470 */
128'hfc0999e39aa2028784339a22408989b3, /* 1471 */
128'h6aa26a4269e274a279028526744270e2, /* 1472 */
128'hc23e47f500f110234799713980826121, /* 1473 */
128'h8ed10106161b8edd030007b70086969b, /* 1474 */
128'h858a4601440dc43684aafc06f426f822, /* 1475 */
128'hf0ef85263e800593e919c53ff0ef8526, /* 1476 */
128'hfc79347d8082612174a2744270e2d91f, /* 1477 */
128'h23213823bffc07b7db0101134d18bfcd, /* 1478 */
128'h342322913c2324813023241134239fb9, /* 1479 */
128'h01f104131ce7f56349013ffc07372331, /* 1480 */
128'h1e051863892ac09ff0ef84aa85a29801, /* 1481 */
128'hb02365e020ef20000513e7991a04b783, /* 1482 */
128'h85a2200006131e0503631a04b5031aa4, /* 1483 */
128'h37171cf76b6347210c044783123010ef, /* 1484 */
128'h400407b753b897ba078ac02707130000, /* 1485 */
128'h67050d44278300e7fd63cc981ff78793, /* 1486 */
128'hf8dc00d773630147d69307a680070713, /* 1487 */
128'hf9938b8506f48f2309b449830a044783, /* 1488 */
128'h80a30b344783c7890e244783e7810019, /* 1489 */
128'h4783c7898b890a04478300098a6308f4, /* 1490 */
128'h8613091407130e24478306f48fa309c4, /* 1491 */
128'h468109d405130a844783fcdc07c60c84, /* 1492 */
128'h0087979b00074583fff74783e0fc07c6, /* 1493 */
128'h4685c39197aeffe745839fad0105959b, /* 1494 */
128'h0dd4478302f585b30e04458300098c63, /* 1495 */
128'hfca714e30621070de21c07ce02b787b3, /* 1496 */
128'h979b468508d4470308e4478304098f63, /* 1497 */
128'h470397ba08c447039fb90087171b0107, /* 1498 */
128'h07ce02e787b30dd4478302f707330e04, /* 1499 */
128'h171b0187979b08a4470308b44783f8fc, /* 1500 */
128'h47039fb90087171b089447039fb90107, /* 1501 */
128'h4783f4fc07a6c319f4fc54d89fb90884, /* 1502 */
128'hce81e3918bfd09c44783c7898b850a04, /* 1503 */
128'hed35e0bff0ef852645850af006134685, /* 1504 */
128'h8b850e0446830af447830af407a34785, /* 1505 */
128'h8663c79954dc08f4aa2300a6979bc7b9, /* 1506 */
128'h969b0dd44783f8dc07a60d4427830009, /* 1507 */
128'h80230a74478308d4ac2302f686bb00a6, /* 1508 */
128'h23813483854a240134032481308308f4, /* 1509 */
128'h50fc8082250101132281398323013903, /* 1510 */
128'h278527058bfd8b7d0057d79b00a7d71b, /* 1511 */
128'h1a04b503892abf4d08f4aa2302f707bb, /* 1512 */
128'hbf555951bf651a04b0234c0020efd169, /* 1513 */
128'h2281382322113c23dc010113bf455929, /* 1514 */
128'he16302f5886347892321302322913423, /* 1515 */
128'h230134032381308354a9c585468102b7, /* 1516 */
128'h80822401011322813483220139038526, /* 1517 */
128'h0613842e4685fef760e34705ffc5879b, /* 1518 */
128'h059bf57184aad1fff0ef892a45850b90, /* 1519 */
128'h85a2980101f10413f1e9258199f5ffe4, /* 1520 */
128'h0493f7d50b944783e51998dff0ef854a, /* 1521 */
128'he44ee84aec267179b74d84aab75ddf40, /* 1522 */
128'h0079f6930ff5f99308154783f022f406, /* 1523 */
128'hf0ef84aa45850b3006138edd892e9be1, /* 1524 */
128'h00091c6300f51e63842a57b5c519cc7f, /* 1525 */
128'h15e010ef8526842a875ff0ef852685ca, /* 1526 */
128'h69a2694264e2740270a28522013505a3, /* 1527 */
128'h2881382328113c23d601011380826145, /* 1528 */
128'h2741382327313c232921302328913423, /* 1529 */
128'h2581382325713c232761302327513423, /* 1530 */
128'he963478923b13c2325a1302325913423, /* 1531 */
128'h07b79f3dbff7879bbffc07b74d180ac7, /* 1532 */
128'h0000451784ae8b32892abfe787933ffc, /* 1533 */
128'h0016779307e9460300e7eb6304450513, /* 1534 */
128'h0413f96ff0ef0665051300004517e7b9, /* 1535 */
128'h2881348329013403298130838522f840, /* 1536 */
128'h26813a8327013a032781398328013903, /* 1537 */
128'h24813c8325013c0325813b8326013b03, /* 1538 */
128'h270380822a01011323813d8324013d03, /* 1539 */
128'h0045aa83db4503e50513000045170989, /* 1540 */
128'hf7bb0005ac83e79102eaf7bb060a8163, /* 1541 */
128'hf24ff0ef0445051300004517cb8902ec, /* 1542 */
128'he3994b8502eadabb02c92783bf415429, /* 1543 */
128'h478189d6856200c488138c0a009c9c9b, /* 1544 */
128'h02e8f33b0017859b000828834e114e85, /* 1545 */
128'hee4ff0ef03c505130000451700030d63, /* 1546 */
128'h202302e8d33bb7f14b814a814c81b7c1, /* 1547 */
128'h8b850107c78397a6078e020880630065, /* 1548 */
128'h09bb0ffbfb9300dbebb300be96bbcb89, /* 1549 */
128'h000b8963fbc596e387ae051108210133, /* 1550 */
128'h0a13f00600e301e50513000045178a09, /* 1551 */
128'h842af94ff0ef854a85d2fe0a7a1302f1, /* 1552 */
128'h0106161b09ea478309fa4603ee0519e3, /* 1553 */
128'h01367a63963e09da47839e3d0087979b, /* 1554 */
128'hb5c1e56ff0ef00e505130000451785ce, /* 1555 */
128'hc71989b60017f7130a7a46830084c783, /* 1556 */
128'h450547010016e993c3990fe6f9938b89, /* 1557 */
128'h0017581b4b189726070e0017059b4611, /* 1558 */
128'h0027571b00b517bb0208046300187813, /* 1559 */
128'hd99b4187d79b8b050189999b0187979b, /* 1560 */
128'h92e3872e0ff9f99300f9e9b3c70d4189, /* 1561 */
128'h4517ef898b850a6a478302d98263fcc5, /* 1562 */
128'hfff7c793b591268020effc2505130000, /* 1563 */
128'h4517cb898b8509ba4783bfd100f9f9b3, /* 1564 */
128'h02e3b51d547ddbaff0efff2505130000, /* 1565 */
128'h0af006134685e3958b850afa4783e20b, /* 1566 */
128'h0afa07a34785e569a21ff0ef854a4585, /* 1567 */
128'h0880049308f92a2300a7979b0e0a4783, /* 1568 */
128'h86260ff6f69301acd6bb08c00d934d01, /* 1569 */
128'h0ff4f4932485ed499f1ff0ef854a4585, /* 1570 */
128'h019ad6bb08f00d134c81ffb492e32d21, /* 1571 */
128'he9359cbff0ef854a458586260ff6f693, /* 1572 */
128'h0d934d61ffa492e32ca10ff4f4932485, /* 1573 */
128'hd6bb45858656000c26834c818aa609b0, /* 1574 */
128'h2a85e13999dff0ef854a0ff6f6930196, /* 1575 */
128'h0ff4f493248dffac90e30ffafa932ca1, /* 1576 */
128'h854a458509c0061386defdb498e30c11, /* 1577 */
128'h0a7a4783d4fb0de34785ed19975ff0ef, /* 1578 */
128'hf0ef854a458509b00613468501379b63, /* 1579 */
128'h854a45850a70061386cebb3d842a957f, /* 1580 */
128'he406e0221141b32ddd79842a945ff0ef, /* 1581 */
128'hb303679c681c00055e63804ff0ef842a, /* 1582 */
128'h8302014160a264028522000307630187, /* 1583 */
128'hfc06f426713980820141640260a24505, /* 1584 */
128'h5529478500f5866384aa4791f04af822, /* 1585 */
128'h07c4d78300f110230370079304f59263, /* 1586 */
128'hc24a8526858a46010107979b4955842e, /* 1587 */
128'hc24a00f110234799ed19d52ff0efc43e, /* 1588 */
128'h8526858a4601c43e478900f41f634791, /* 1589 */
128'h80826121790274a2744270e2d34ff0ef, /* 1590 */
128'h4f5c6918ee09b7cdc402fef414e34785, /* 1591 */
128'h00e7f46385be27814f1887ae00f5f363, /* 1592 */
128'h8082c2cff06f02c50823dd0c0007059b, /* 1593 */
128'hf8a2070d4b9c711910000737691c8082, /* 1594 */
128'hfc5ee0dae4d6e8d2eccef0caf4a6fc86, /* 1595 */
128'hc509f11ff0ef842ac17c8fd9f466f862, /* 1596 */
128'h0000451702042423eb8d6b9c679c681c, /* 1597 */
128'h744670e6f8500493bacff0efe0450513, /* 1598 */
128'h7be26b066aa66a4669e674a679068526, /* 1599 */
128'hf0eff3e54481541c808261097ca27c42, /* 1600 */
128'h2c2302f4082347851af42c23478df93f, /* 1601 */
128'h3b5010ef7d000513ba2ff0ef85220204, /* 1602 */
128'h2783f94584aa97826b9c679c8522681c, /* 1603 */
128'h478508f422231a04282318042e230884, /* 1604 */
128'hf0ef852245814601b72ff0ef8522d85c, /* 1605 */
128'h00ef8522f14984aacf2ff0ef8522f1df, /* 1606 */
128'h8737681c00f1102347a1000505a345d0, /* 1607 */
128'h0aa00713e3991aa007138ff94bdc00ff, /* 1608 */
128'hbf8ff0efc23ec43a8522858a460147d5, /* 1609 */
128'h07b700f715630aa0079300c14703e911, /* 1610 */
128'h0a934a55037009933e900913cc1c8002, /* 1611 */
128'h40000cb780020c3700ff8bb74b050290, /* 1612 */
128'hf0efc402c252013110238522858a4601, /* 1613 */
128'hc25a4bdc015110234c18681ce13dbb6f, /* 1614 */
128'hc43e0197e7b301871563c43e0177f7b3, /* 1615 */
128'hca6347b2ed1db8eff0ef8522858a4601, /* 1616 */
128'h2c5010ef3e80051306090863397d0007, /* 1617 */
128'h8001073700e68563800207374c14bf45, /* 1618 */
128'h06041e23d45c8b8541e7d79bc43ccc18, /* 1619 */
128'h02f51f63f9200793b55d18f40ca34785, /* 1620 */
128'hed09c34ff0ef85224581c04ff0ef8522, /* 1621 */
128'h4585bfd118f40c2347850007d663443c, /* 1622 */
128'hc805051300004517d965c1cff0ef8522, /* 1623 */
128'h551cb58584aab595fa100493a10ff0ef, /* 1624 */
128'hfed6e352e74eeb4aef26f706f3227161, /* 1625 */
128'he3b54401e6eeeaeaeee6f2e2f6defada, /* 1626 */
128'hc783c7b1199bc783193010ef45018baa, /* 1627 */
128'h460104f110234789e7b5180b8ca3198b, /* 1628 */
128'h842aabaff0efc482c2be855e008c479d, /* 1629 */
128'h46014495cf818b851b8ba783120500e3, /* 1630 */
128'h34fd100503e3842aaa0ff0ef855e008c, /* 1631 */
128'h842ad99ff0ef855ea031020ba423f4fd, /* 1632 */
128'h6a1a69ba695a64fa741a70ba8522d55d, /* 1633 */
128'h615d6db66d566cf67c167bb67b567af6, /* 1634 */
128'h855e0407c163180b8c23048ba7838082, /* 1635 */
128'h908102051493101010ef4501b16ff0ef, /* 1636 */
128'hf155842ab36ff0ef855e45853e800913, /* 1637 */
128'h6ee30dd010ef85260007cc63048ba783, /* 1638 */
128'h400007b7bfe916b010ef0640051312a9, /* 1639 */
128'ha6238b8541e7d79b048ba78300fbac23, /* 1640 */
128'h1aa60f63450dbf0506fb9e23478502fb, /* 1641 */
128'h40010637a029400406370ea61ee34511, /* 1642 */
128'h29978a9d0036d61b00cbac234006061b, /* 1643 */
128'h460396ce964e068a8a3d212989930000, /* 1644 */
128'h02d606bb018ba88345051086a6830f86, /* 1645 */
128'ha823180bae231a0ba8238a0500c7d61b, /* 1646 */
128'h8abd0107d69b08dba22308dba42304cb, /* 1647 */
128'h090ba8231408dc63090ba62300d5183b, /* 1648 */
128'h003f06b70107979b14068e6302cba683, /* 1649 */
128'h07854721938117828fd98ff50107571b, /* 1650 */
128'hb0230a0bbc23030787b300e797b30709, /* 1651 */
128'hb0230c0bbc230c0bb8230c0bb4230c0b, /* 1652 */
128'ha6230107d463200007930afbb8230e0b, /* 1653 */
128'ha82300e7f46320000793090ba70308fb, /* 1654 */
128'h471100e78e63577d04cba783c21508fb, /* 1655 */
128'hc4be04e11023855e008c46010107979b, /* 1656 */
128'h07cbd78304f11023479d902ff0efc282, /* 1657 */
128'hc4bec2ca855e008c0107979b46014955, /* 1658 */
128'h08fbaa234785e40516e3842a8e4ff0ef, /* 1659 */
128'h1ae3842ac9aff0ef855e08fb80a357fd, /* 1660 */
128'he0ef855e00b545830f7000ef855ee205, /* 1661 */
128'h54075a63018ba703e0051fe3842affbf, /* 1662 */
128'h10230370079304fba0232789100007b7, /* 1663 */
128'h855e0107979b108c460107cbd78306f1, /* 1664 */
128'h04934905d2caed05880ff0efd4bed2ca, /* 1665 */
128'h06f11023988102091a93033007930bf1, /* 1666 */
128'he826855e108c08104b210a854a11d482, /* 1667 */
128'hfe0a16e33a7dc131850ff0efd05aec56, /* 1668 */
128'hbd9940030637a7a940020637bb45842a, /* 1669 */
128'hb54d08bba82300b515bb89bd0165d59b, /* 1670 */
128'h8fd501e7569b8ff50027979b16f16685, /* 1671 */
128'h05374098b5558b1d938100f7571b1782, /* 1672 */
128'h8fd50087161b0187179b0187569b00ff, /* 1673 */
128'h8ef1f00706138fd167410087569b8e69, /* 1674 */
128'h169b0187559b40d804fbaa2327818fd5, /* 1675 */
128'h8ecd0087571b8de90087159b8ecd0187, /* 1676 */
128'h00638b3d0187d71b04ebac238f558f71, /* 1677 */
128'h00ebac238001073720d7026346892127, /* 1678 */
128'h20000737040ba7830007596302d79713, /* 1679 */
128'h1863800107b7018ba70304fba0238fd9, /* 1680 */
128'h040ba903639cd1678793000047971ef7, /* 1681 */
128'h00002497020d1a13044ba783f0be4d05, /* 1682 */
128'h83f979130ff1079300f9793302c48493, /* 1683 */
128'h77b300e797bb478540980a05fe07fc13, /* 1684 */
128'h0b1b4a81017d8b3716078563278100f9, /* 1685 */
128'h00f977b340dc0007ac8397d6109c840b, /* 1686 */
128'h8d6345a1400007b7140781630197f7b3, /* 1687 */
128'h100005b700fc88634591200007b700fc, /* 1688 */
128'h8daa971ff0ef855e0015b59340bc85b3, /* 1689 */
128'h073700ec8d6347a1400007370e051c63, /* 1690 */
128'h40fc8cb3100007b700ec886347912000, /* 1691 */
128'h409cdfdfe0ef855e02fbaa23001cb793, /* 1692 */
128'h102347994d850ce79163470d01a78663, /* 1693 */
128'he7b317c12d81810007b7d33e47d50af1, /* 1694 */
128'he162855e110c040007930110d53e00fd, /* 1695 */
128'h8bbd010c4783e941e91fe0efc93ee552, /* 1696 */
128'ha58314079a631afba823409c09b79463, /* 1697 */
128'h18fbae2308bba2230017b79317ed088b, /* 1698 */
128'hfe07fd930ff10793947ff0ef855e4601, /* 1699 */
128'h4601475507cbd7830af1102303700793, /* 1700 */
128'hd53ee03ad33a8cee855e110c0107979b, /* 1701 */
128'hd33a0af1102347b56702e915e35fe0ef, /* 1702 */
128'he43e855e110c0110040007134791d502, /* 1703 */
128'h0e050c63e0dfe0efe03ac93ae552e16e, /* 1704 */
128'ha823017d85b74785f3ed37fd670267a2, /* 1705 */
128'h840585934601180bae23096ba2231afb, /* 1706 */
128'h04a1eafa94e347a10a918c9ff0ef855e, /* 1707 */
128'h00003517e6f49fe3ea87879300002797, /* 1708 */
128'h1737b61ddf400413cbdfe0ef75c50513, /* 1709 */
128'h00ebac2380020737b519a007071b8001, /* 1710 */
128'h4905bbc580030737de075ee303079713, /* 1711 */
128'h3ac54a159881190201000ab70ff10493, /* 1712 */
128'h47d508f110234799020a08633a7d0905, /* 1713 */
128'hf426c556855e010c040007931030c33e, /* 1714 */
128'h83a54cdcd0051ce3d61fe0efdc3ef84a, /* 1715 */
128'h0087961bf006869366c144dcfbe18b85, /* 1716 */
128'h040ba70302e796938fd18ff50087d79b, /* 1717 */
128'h472db35d04fba02300876793da06d9e3, /* 1718 */
128'h2583974e837902079713eaf768e34581, /* 1719 */
128'h869300ff0537040d859366c1b5451187, /* 1720 */
128'h0187971b0187d61b0d91000da783f006, /* 1721 */
128'h8ff58f510087d79b8e690087961b8f51, /* 1722 */
128'h46a5008ca703fdb59ee3fefdae238fd9, /* 1723 */
128'h06b7018ba60300f6f8638bbd00c7579b, /* 1724 */
128'h078acfa686930000269704d61c638003, /* 1725 */
128'ha68308fbae230087171b1487a78397b6, /* 1726 */
128'hd71b8fd10186d61b8ff917fd67c100cc, /* 1727 */
128'h3e800613c305c38d03f7771327810126, /* 1728 */
128'h06bb02f757bb8a8d0106d69b02e6073b, /* 1729 */
128'haa231b0ba7830adba2230afba02302d6, /* 1730 */
128'h08fba62320000793c79919cba7831afb, /* 1731 */
128'h062300051523484000ef855e08fba823, /* 1732 */
128'h8793ccccd6b7aaaab7b708cba7030005, /* 1733 */
128'h00d036b327818ef98ff9ccc68693aaa7, /* 1734 */
128'h0f068693f0f0f6b79fb500f037b30686, /* 1735 */
128'h8693ff0106b79fb5068a00d036b38ef9, /* 1736 */
128'h161376c19fb5068e00d036b38ef9f006, /* 1737 */
128'hb783d11c9fb9071200e037338f750207, /* 1738 */
128'hd68307abd70302c7d7b3ed1092010a8b, /* 1739 */
128'h598585930000359784aa06fbc603074b, /* 1740 */
128'h070ba803a95fe0effef5362302450513, /* 1741 */
128'h0108571b0088579b06cbc603077bc883, /* 1742 */
128'h0ff777130ff878130ff7f7930188569b, /* 1743 */
128'he0ef04d4851357658593000035972681, /* 1744 */
128'h85135725859300003597074ba603a5ff, /* 1745 */
128'he0ef8a3d8abd0146561b0106569b0624, /* 1746 */
128'hb8d102fba42347856dc010ef8526a3ff, /* 1747 */
128'hb683400407b704fba0232785100007b7, /* 1748 */
128'h4f05051300003517e691ecf76ce31a0b, /* 1749 */
128'hc78304fba0230017079b70000737bb95, /* 1750 */
128'hce910027f6931adba42303f7f6930c46, /* 1751 */
128'ha70304eba0230217071bc68900c7f693, /* 1752 */
128'ha783c7998b8504eba02301076713040b, /* 1753 */
128'ha783040baa0304fba02300c7e793040b, /* 1754 */
128'h249700fa7a33855e4601088ba583044b, /* 1755 */
128'h00002b174a85db4ff0efbaa484930000, /* 1756 */
128'h409cbeec8c9300002c974c2dbbcb0b13, /* 1757 */
128'h00002917cbb5278100fa77b300fa97bb, /* 1758 */
128'h4703409c10000db720000d37b9c90913, /* 1759 */
128'h270340dc04f718630017b79317ed0049, /* 1760 */
128'h061300894683c3a18ff900fa77b30009, /* 1761 */
128'hc131debfe0ef855e0fb6f69345850b70, /* 1762 */
128'ha783ddbfe0ef855e45850b7006134681, /* 1763 */
128'haa2308fba223180bae231a0ba823088b, /* 1764 */
128'h04a1fb9911e30931973fe0ef855e035b, /* 1765 */
128'h925fe0ef3c45051300003517f7649fe3, /* 1766 */
128'h00d789634721400006b700092783bb6d, /* 1767 */
128'haa230017b71341b787b301a786634711, /* 1768 */
128'h808ff0ef855e408c933fe0ef855e02eb, /* 1769 */
128'ha823409ce79d0046f79300892683f941, /* 1770 */
128'ha2230017b79317ed088ba583ef8d1afb, /* 1771 */
128'h855ecb0ff0ef855e460118fbae2308bb, /* 1772 */
128'h0b7006130ff6f693bb91fd319fdfe0ef, /* 1773 */
128'h65e34581b7c9f521d31fe0ef855e4585, /* 1774 */
128'hbf6d11872583974e837902079713fcfc, /* 1775 */
128'h1023478d6da000ef06cb851300ec4641, /* 1776 */
128'hc4be0107979b008c460107cbd78304f1, /* 1777 */
128'hec051b63842a96ffe0efc2be47d5855e, /* 1778 */
128'h06fb9e2304e157830007d663018ba783, /* 1779 */
128'h460107cbd783c2be479d04f1102347a5, /* 1780 */
128'h842a93bfe0efc4be855e0107979b008c, /* 1781 */
128'h018ba50345e6475647c646b6ea051163, /* 1782 */
128'h06bba42306eba22306fba02304dbae23, /* 1783 */
128'h45098a3d01a6d61bf2c51a6340000637, /* 1784 */
128'h0637f0a609634505f0c543638ca602e3, /* 1785 */
128'hf06ffa100413f0eff06f2006061b4001, /* 1786 */
128'h8082557d8082557d80824501c56ce54f, /* 1787 */
128'h439c8ee7879300004797808218b50d23, /* 1788 */
128'h00004717842ae406e02247851141ef9d, /* 1789 */
128'h5563ae2fe0ef852212a000ef8cf72c23, /* 1790 */
128'h13e000ef02c00513fc5ff0ef85220005, /* 1791 */
128'h4501808201414501640260a20dc000ef, /* 1792 */
128'h90636394631c8a670713000047178082, /* 1793 */
128'he406372505130000351785aa114102e7, /* 1794 */
128'ha60380820141853e478160a2f60fe0ef, /* 1795 */
128'h41488082853ebfd187b600a604630fc7, /* 1796 */
128'h10354703c105fbdff0efe42eec061101, /* 1797 */
128'h0c630ff007930815470302b7006365a2, /* 1798 */
128'h610560e25535eb3fe06f610560e200f7, /* 1799 */
128'he4261101bfcdf8400513bfe545018082, /* 1800 */
128'hf0ef842acd09f7dff0ef84aee822ec06, /* 1801 */
128'h64a2644260e2e0800f840413e501cf0f, /* 1802 */
128'h6907879300003797bfd5553580826105, /* 1803 */
128'h80820f8505138082c3980015071b4388, /* 1804 */
128'h37971101808243886787879300003797, /* 1805 */
128'h84beec06e4266380e8227da787930000, /* 1806 */
128'h47838082610564a2644260e200941763, /* 1807 */
128'h3797b7d56000a9cff0ef8522c78119a4, /* 1808 */
128'ha72300003797e79ce39c7aa787930000, /* 1809 */
128'h67987927879300003797e50880826207, /* 1810 */
128'h3497e4a6711d8082e308e518e11ce788, /* 1811 */
128'hf456f852fc4e6080e8a277a484930000, /* 1812 */
128'h89aae0caec86e06ae466e862ec5ef05a, /* 1813 */
128'h250a8a9300003a97260a0a1300003a17, /* 1814 */
128'h258b8b9300003b97258b0b1300003b17, /* 1815 */
128'h15634d297b4c8c9300002c9700050c1b, /* 1816 */
128'h7aa27a4279e2690664a660e664460294, /* 1817 */
128'h0513000035176d026ca26c426be27b02, /* 1818 */
128'h4c1cc7914901541cddcfe06f61252fe5, /* 1819 */
128'h855a0fc42603681c89560007c3638952, /* 1820 */
128'he0ef855e85ca00090663dbefe0ef638c, /* 1821 */
128'hda4fe0ef856685e200978e63601cdb2f, /* 1822 */
128'h222010ef73c505130000251701a98863, /* 1823 */
128'h4401e04ae426ec06e8221101b7716000, /* 1824 */
128'hcbad511ccbbd4d5ccfad44014d1cc141, /* 1825 */
128'h1c00059384aa892ec7ad639cc7bd651c, /* 1826 */
128'h4799c57c57fdcd21842a0f8010ef4505, /* 1827 */
128'h03253023e90410f502a347850ef52c23, /* 1828 */
128'h91c78793fffff797e65ff0ef04052823, /* 1829 */
128'h18f430231b6787930000179716f43c23, /* 1830 */
128'h2e23681c18f434231a67879300001797, /* 1831 */
128'he99ff0ef10f400230247c78385220ea4, /* 1832 */
128'h106f80826105690264a2644260e28522, /* 1833 */
128'h65186294611c38e68693000036970b40, /* 1834 */
128'h0127d713e11897360017671302d786b3, /* 1835 */
128'h17bb40f007b300f7553b93ed836d8f3d, /* 1836 */
128'h5f05051300003517808225018d5d00f7, /* 1837 */
128'h842afefff0efe022e4061141fc3ff06f, /* 1838 */
128'h2501640260a28d410105151bfe9ff0ef, /* 1839 */
128'h041bfdbff0efe022e406114180820141, /* 1840 */
128'h60a28d4115029001fd1ff0ef14020005, /* 1841 */
128'h0785fff5c703058587aa808201416402, /* 1842 */
128'h00c7896387aa962a8082fb75fee78fa3, /* 1843 */
128'h8082fb65fee78fa30785fff5c7030585, /* 1844 */
128'hc7030585eb09001786930007c70387aa, /* 1845 */
128'hb7d587b68082fb75fee78fa30785fff5, /* 1846 */
128'h001786930007c70387b68082e21987aa, /* 1847 */
128'h0fa300178713fff5c6830585963efb7d, /* 1848 */
128'h8082000780a300c715638082e291fed7, /* 1849 */
128'h07bbfff5c783000547030585b7cd87ba, /* 1850 */
128'hf37d0505e3994187d79b0187979b40f7, /* 1851 */
128'h0585a839478100c59463962e8082853e, /* 1852 */
128'h0187979b40f707bbfff5c78300054703, /* 1853 */
128'hf5938082853eff790505e3994187d79b, /* 1854 */
128'h0505c399808200b79363000547830ff5, /* 1855 */
128'h9363000547830ff5f59380824501bfcd, /* 1856 */
128'h0007c70387aabfcd0505dffd808200b7, /* 1857 */
128'he8221101bfcd0785808240a78533e701, /* 1858 */
128'hf593952265a2fe5ff0efec06842ae42e, /* 1859 */
128'hfe857be3157d00b78663000547830ff5, /* 1860 */
128'h856387aa95aa80826105644260e24501, /* 1861 */
128'h0785808240a78533e7010007c70300b7, /* 1862 */
128'hea9940c785330007c68387aa862ab7fd, /* 1863 */
128'hfe081be3000748030705fed80fe38082, /* 1864 */
128'h0007c60387aa86aabfcd872eb7d50785, /* 1865 */
128'h4803070500c80a638082ea1140d78533, /* 1866 */
128'hbff90785bfd5872e8082fe081be30007, /* 1867 */
128'h0785fee68fe380824501eb1900054703, /* 1868 */
128'h1101bfd587aeb7e50505fafd0007c683, /* 1869 */
128'h00003797e519842a84aeec06e426e822, /* 1870 */
128'hf9dff0ef85a68522cc1163803ec78793, /* 1871 */
128'h3c07b82300003797ef8100044783942a, /* 1872 */
128'h85a68082610564a2644260e285224401, /* 1873 */
128'h0023c78100054783c519f9fff0ef8522, /* 1874 */
128'h1101bfd93aa7b2230000379705050005, /* 1875 */
128'hf0ef8526842ac891e822ec066104e426, /* 1876 */
128'h644260e2e008050500050023c501f73f, /* 1877 */
128'hcf9900054783c11d8082610564a28526, /* 1878 */
128'h8082e3110017c703ce810007c68387aa, /* 1879 */
128'h80824501b7e5078900d780a300e78023, /* 1880 */
128'h808204c79063963e87aacb9d00757793, /* 1881 */
128'h469d00c508b3872aff6d377d8fd507a2, /* 1882 */
128'h87335761003657930106ef6340e88833, /* 1883 */
128'h0ff5f6934725bfc1963a97aa078e02e7, /* 1884 */
128'hfeb78fa30785bfe1fef73c230721bfd1, /* 1885 */
128'h87aacb9d8b9d00a5e7b300b50a63bf6d, /* 1886 */
128'h07a1ff8738030721808202c79e63963e, /* 1887 */
128'h00365713ff06e8e340f88833ff07bc23, /* 1888 */
128'h00e507b3963e95ba070e02f707b357e1, /* 1889 */
128'h0585bfe1469d00c508b387aa872ebfc1, /* 1890 */
128'hf0227179bf65fee78fa30785fff5c703, /* 1891 */
128'hf0efe02ee84af406e432ec26852e842a, /* 1892 */
128'h00c564636582892ace1184aa6622dcdf, /* 1893 */
128'h0023f79ff0ef944a864a8522fff60913, /* 1894 */
128'h8082614564e269428526740270a20004, /* 1895 */
128'hf57ff0ef00a5e963842ae406e0221141, /* 1896 */
128'h00c506b395b280820141640260a28522, /* 1897 */
128'h0005c78315fdd7e500e587b340b60733, /* 1898 */
128'h478100c51563962ab7fd00f6802316fd, /* 1899 */
128'hfbed9f990005c703000547838082853e, /* 1900 */
128'h4783808200c51363962ab7dd05850505, /* 1901 */
128'h842af0227179bfc50505feb78de30005, /* 1902 */
128'hd1fff0ef89aee84af406e44eec26852e, /* 1903 */
128'h0005091bd13ff0ef8522c8890005049b, /* 1904 */
128'h694264e2740270a28522440100995b63, /* 1905 */
128'hf0ef397d852285ce86268082614569a2, /* 1906 */
128'h14630ff5f593962abfe90405d175f8bf, /* 1907 */
128'h0be300150793000547038082450100c5, /* 1908 */
128'h00c7ef630ff5f59347c1b7ed853efeb7, /* 1909 */
128'h0007c7038082853e4781e60187aa2601, /* 1910 */
128'hc31d00757713b7f5367d0785feb71ce3, /* 1911 */
128'h0007c80387aa0007069b40e7873b47a1, /* 1912 */
128'h938102071793faf5078536fdfcb81ce3, /* 1913 */
128'h0107179300b7e733008597938e1d953e, /* 1914 */
128'h87aa27018edd00365713020796938fd9, /* 1915 */
128'h0785f8b71fe30007c703d24d8a1deb11, /* 1916 */
128'h00d80a63008785130007b803bfcd367d, /* 1917 */
128'hbfa5fef51be30785f8b712e30007c703, /* 1918 */
128'h079300054703e7a9419cb7f1377d87aa, /* 1919 */
128'h8793000017970015470308f711630300, /* 1920 */
128'h071bc6898a850006c68300e786b3cf67, /* 1921 */
128'h470304d71b63078006930ff777130207, /* 1922 */
128'h47c1c3b10447f7930007c78397ba0025, /* 1923 */
128'h07930005470302f71c6347c14198c19c, /* 1924 */
128'h0713000017170015478302f716630300, /* 1925 */
128'h0207879bc7098b0500074703973eca67, /* 1926 */
128'h8082050900e79363078007130ff7f793, /* 1927 */
128'h006c842ee8221101bf6d47a9bf7d47a1, /* 1928 */
128'h1817468100c16583f63ff0efc632ec06, /* 1929 */
128'h06330007079b00054703c62808130000, /* 1930 */
128'hec0500089863044678930006460300f8, /* 1931 */
128'h8b6300467893808261058536644260e2, /* 1932 */
128'h050502d586b3feb7f4e3fd07879b0008, /* 1933 */
128'h0ff7f793fe07079bc6098a09b7d196be, /* 1934 */
128'hf426f8227139b7e1e008b7cdfc97879b, /* 1935 */
128'hf0ef84b2842ae42e00063023f04afc06, /* 1936 */
128'h790274a2744270e25529e90165a2b0df, /* 1937 */
128'hf5dff0ef8522082c892a862e80826121, /* 1938 */
128'h07858f81cb010007c703fe8782e367e2, /* 1939 */
128'hb7e94501e088fcf718e347a9fd279be3, /* 1940 */
128'hf2dff06f00e6846302d0071300054683, /* 1941 */
128'h40a0053360a2f23ff0efe40605051141, /* 1942 */
128'hf0dff0ef842ee406e022114180820141, /* 1943 */
128'hea6302d704630007c70304b00693601c, /* 1944 */
128'h0141640260a202d70e630470069300e6, /* 1945 */
128'h16e306b0069302d7076304d006938082, /* 1946 */
128'hfce69fe3052a069007130017c683fed7, /* 1947 */
128'he01c078d00e69863042007130027c683, /* 1948 */
128'he8221101bfd50789bff1052a052ab7e9, /* 1949 */
128'h00c16583e0fff0efc632ec06006c842e, /* 1950 */
128'h079b00054703b0e80813000018174681, /* 1951 */
128'h9863044678930006460300f806330007, /* 1952 */
128'h7893808261058536644260e2ec050008, /* 1953 */
128'h86b3feb7f4e3fd07879b00088b630046, /* 1954 */
128'hfe07079bc6098a09b7d196be050502d5, /* 1955 */
128'h1141b7e1e008b7cdfc97879b0ff7f793, /* 1956 */
128'h04b00693601cf87ff0ef842ee406e022, /* 1957 */
128'h0470069300e6ea6302d704630007c703, /* 1958 */
128'h04d0069380820141640260a202d70e63, /* 1959 */
128'h0017c683fed716e306b0069302d70763, /* 1960 */
128'h07130027c683fce69fe3052a06900713, /* 1961 */
128'h052a052ab7e9e01c078d00e698630420, /* 1962 */
128'he589842ae406e0221141bfd50789bff1, /* 1963 */
128'h00001797fff5c70300a405b395bff0ef, /* 1964 */
128'h8b1100074703973efff58513a3478793, /* 1965 */
128'h7ae3157d80820141557d640260a2e719, /* 1966 */
128'hf77d8b1100074703973e00054703fea4, /* 1967 */
128'hd7dff06f014105054581462960a26402, /* 1968 */
128'h0723812100a107a31141fa5ff06f4581, /* 1969 */
128'h45a9462547818082014100e1550300a1, /* 1970 */
128'hf693fd07069b8082853ee31900054703, /* 1971 */
128'hfd07879b9fb902f587bb00d667630ff6, /* 1972 */
128'h00a04563842ee406e0221141bff90505, /* 1973 */
128'hf0ef357d02b455bb45a900b7f86347a5, /* 1974 */
128'h0513014160a2640202a4753b4529fe7f, /* 1975 */
128'h33230000371707fe47854ac0006f0305, /* 1976 */
128'he82211018082f6f7332300003717f6f7, /* 1977 */
128'h85aa84ae862ee426f584041300003417, /* 1978 */
128'he00c95a660e2600ca2fff0efec066008, /* 1979 */
128'h87930000379711418082610564a26442, /* 1980 */
128'h638cf2278793000037976380e022f267, /* 1981 */
128'hba5fd0ef9d81e4068005051300003517, /* 1982 */
128'h11418302014160a2640283220000100f, /* 1983 */
128'h557d008503638f2fa0ef8432e406e022, /* 1984 */
128'hf22271698082450180820141640260a2, /* 1985 */
128'hea4aee26f606852289aae64e01258413, /* 1986 */
128'hf0ef852600a404b30505fe8ff0ef892e, /* 1987 */
128'h0793fff5071bee5ff0ef95260505fdcf, /* 1988 */
128'h8522e8a7a9230000379704e7ee631ff0, /* 1989 */
128'hf0ef5ba505130000251784aafbaff0ef, /* 1990 */
128'hf0ef852204a7f2630ff007939526facf, /* 1991 */
128'hf8eff0ef59c5051300002517842af9cf, /* 1992 */
128'haf5fd0ef764505130000251700a405b3, /* 1993 */
128'h07938082615569b2695264f2741270b2, /* 1994 */
128'h10000613b755e2f72b23000037172000, /* 1995 */
128'h55858593000025978cdff0ef850a4581, /* 1996 */
128'h096302f0079301294703e54ff0ef850a, /* 1997 */
128'he64ff0ef850a736585930000259700f7, /* 1998 */
128'hdf07879300003797e5cff0ef850a85a2, /* 1999 */
128'ha85fd0ef71c5051300002517858a4390, /* 2000 */
128'hdcf73c2300003717451101f417934405, /* 2001 */
128'h00003797defff0efdcf73c2300003717, /* 2002 */
128'h942300003797de1ff0ef4501baa79a23, /* 2003 */
128'hf0ef854eb9c58593000035974611baa7, /* 2004 */
128'he8221101b799d8879d2300003797eb1f, /* 2005 */
128'h892a08c7df638432478de04ae426ec06, /* 2006 */
128'h956325010004d783da3ff0ef84ae450d, /* 2007 */
128'hd783d8dff0efd6a555030000351708a7, /* 2008 */
128'h00448513ffc4059b06a79a6325010024, /* 2009 */
128'h9b2300003797d71ff0ef4511dfdff0ef, /* 2010 */
128'h4611d5dff0efd3a5550300003517b2a7, /* 2011 */
128'hb185859300003597b2a7912300003797, /* 2012 */
128'h00003597256000ef4535e2dff0ef854a, /* 2013 */
128'h00ef02000513d6fff0ef4515d105d583, /* 2014 */
128'h27850007d783cfa78793000037972400, /* 2015 */
128'hce07879300003797cef7162300003717, /* 2016 */
128'h62850513000025170087cf63278d439c, /* 2017 */
128'hf06f6105690264a260e26442971fd0ef, /* 2018 */
128'h717980826105690264a2644260e2d9bf, /* 2019 */
128'hc78300f10fa347090105c783f022f406, /* 2020 */
128'h470d00e78e6301e1578300f10f230115, /* 2021 */
128'h608505130000251770a2740202e78a63, /* 2022 */
128'h5e05051300002517842a91ffd06f6145, /* 2023 */
128'h614570a265a27402852290ffd0efe42e, /* 2024 */
128'hf06f614505c170a241907402d8dff06f, /* 2025 */
128'h30232291342322813823dc010113ebff, /* 2026 */
128'h0028218006134581893284ae842a2321, /* 2027 */
128'h08282040061385a6eccff0ef22113c23, /* 2028 */
128'hf63ff0ef8522002cf0eff0efe802c44a, /* 2029 */
128'h22013903228134832301340323813083, /* 2030 */
128'hcb81bf67d78300003797808224010113, /* 2031 */
128'h8082cf5ff06f9de58593000035974611, /* 2032 */
128'h7763878e1041e703468000efe4061141, /* 2033 */
128'h10a7a22310e1a02327051001a70300e5, /* 2034 */
128'h01418d5d91011782150260a21007e783, /* 2035 */
128'h84aae426e822ec061101808245018082, /* 2036 */
128'h07b33e8007933a4000ef842afc1ff0ef, /* 2037 */
128'h8d0502a7d533644260e29101150202f4, /* 2038 */
128'hf95ff0efe022e40611418082610564a2, /* 2039 */
128'h07b324078793000f47b7378000ef842a, /* 2040 */
128'h02a7d533014191011502640260a202f4, /* 2041 */
128'hf0ef84aae04ae426e822ec0611018082, /* 2042 */
128'h000f443702a48533346000ef892af63f, /* 2043 */
128'hf45ff0ef0405944a0285543324040413, /* 2044 */
128'h80826105690264a2644260e2fe856ee3, /* 2045 */
128'h842ae04aec06e822009894b7e4261101, /* 2046 */
128'h0433854a89260084f363892268048493, /* 2047 */
128'h690264a2644260e2f47dfa1ff0ef4124, /* 2048 */
128'h808200054503808200b5002380826105, /* 2049 */
128'h07378082020575130147c503100007b7, /* 2050 */
128'h00a70023dfe50207f793014747831000, /* 2051 */
128'h8623f800071300078223100007b78082, /* 2052 */
128'h8623470d0007822300e78023476d00e7, /* 2053 */
128'h88230200071300e78423fc70071300e7, /* 2054 */
128'h00044503842ae406e0221141808200e7, /* 2055 */
128'h0405fa5ff0ef80820141640260a2e509, /* 2056 */
128'h811100f577139c67879300001797b7f5, /* 2057 */
128'h00e580a30007c7830007470397aa973e, /* 2058 */
128'h8121842a002ce8221101808200f58023, /* 2059 */
128'h4503f65ff0ef00814503fd1ff0efec06, /* 2060 */
128'hfb7ff0ef0ff47513002cf5dff0ef0091, /* 2061 */
128'hf43ff0ef00914503f4bff0ef00814503, /* 2062 */
128'he84aec26f022717980826105644260e2, /* 2063 */
128'h7513002c0089553b54e14461892af406, /* 2064 */
128'hf13ff0ef346100814503f81ff0ef0ff5, /* 2065 */
128'h740270a2fe9410e3f0bff0ef00914503, /* 2066 */
128'he84aec26f022717980826145694264e2, /* 2067 */
128'h002c0089553354e103800413892af406, /* 2068 */
128'hf0ef346100814503f3fff0ef0ff57513, /* 2069 */
128'h70a2fe9410e3ec9ff0ef00914503ed1f, /* 2070 */
128'hec06002c110180826145694264e27402, /* 2071 */
128'h00914503ea7ff0ef00814503f13ff0ef, /* 2072 */
128'h43050000100f8082610560e2e9fff0ef, /* 2073 */
128'h8593000025974605da0101138302037e, /* 2074 */
128'h382324113c2395650513000035170765, /* 2075 */
128'h2501ebbfa0ef25213023249134232481, /* 2076 */
128'h3083db6fd0ef2be5051300002517c115, /* 2077 */
128'h01132401390324813483250134032581, /* 2078 */
128'hd94fd0ef2bc505130000251780822601, /* 2079 */
128'hed3fa0ef08082ce58593000025974605, /* 2080 */
128'h0000291704e20bf00493ed2144012501, /* 2081 */
128'h95a66605007491810204159338c90913, /* 2082 */
128'hdf3ff0ef4521ed19250183afb0ef0808, /* 2083 */
128'hde3ff0ef0007c50397ca8b8d00c4579b, /* 2084 */
128'h2501ceefb0ef54020808fbe19c3d47b2, /* 2085 */
128'h00002517bf852965051300002517c919, /* 2086 */
128'hfa858593000025974605b79d27450513, /* 2087 */
128'h051300002517c5112501e03fa0ef4501, /* 2088 */
128'h85a20184961386a20bf00493b7a12865, /* 2089 */
128'h00002517ce8fd0ef2885051300002517, /* 2090 */
128'h90ef0184951385a2cdcfd0ef2c450513, /* 2091 */
128'h051300002517c981c62e0005059b9bef, /* 2092 */
128'ha785051300002517b721cbefd0ef2be5, /* 2093 */
128'h1141900200000023eb7ff0efcb0fd0ef, /* 2094 */
128'h0513000f4537a001e05ff0efe4062501, /* 2095 */
128'h7f870713000027178082450180822405, /* 2096 */
128'he30895360017869300756513157d631c, /* 2097 */
128'h110102b506338082953e055e10d00513, /* 2098 */
128'hc509842afd1ff0efe4328532ec06e822, /* 2099 */
128'h6105644260e28522a4cff0ef45816622, /* 2100 */
128'he40625a5051300002517114180828082, /* 2101 */
128'h450160a2fe1fc0ef20000537c30fd0ef, /* 2102 */
128'hb0002573808245018082450180820141, /* 2103 */
128'h862e86b287361141808202f5553347a9, /* 2104 */
128'hbf4fd0efe406246505130000251785aa, /* 2105 */
128'h952e842ae0221141a001d57ff0ef4505, /* 2106 */
128'h640260a29522408007b3f57ff0efe406, /* 2107 */
128'h45058082450580824505808201418d7d, /* 2108 */
128'h00c684bb842ef406ec26f02271798082, /* 2109 */
128'h80826145450164e2740270a200961863, /* 2110 */
128'h200404136622f33fc0efe432852285b2, /* 2111 */
128'h808245098082450980824509bff92605, /* 2112 */
128'hf06f8082450180824501808280828082, /* 2113 */
128'hf0efe4064780e022400007b71141c57f, /* 2114 */
128'h2401c3bff0efb265051300002517c15f, /* 2115 */
128'h579bb46fd0efb26505130000251785a2, /* 2116 */
128'h8522a00100e787634705c78927810074, /* 2117 */
128'h00000000bfcd923f90efbfe5d45ff0ef, /* 2118 */
128'h00000000000000000000000000000000, /* 2119 */
128'h00000000000000000000000000000000, /* 2120 */
128'h00000000000000000000000000000000, /* 2121 */
128'h00000000000000000000000000000000, /* 2122 */
128'h00000000000000000000000000000000, /* 2123 */
128'h00000000000000000000000000000000, /* 2124 */
128'h00000000000000000000000000000000, /* 2125 */
128'h00000000000000000000000000000000, /* 2126 */
128'h00000000000000000000000000000000, /* 2127 */
128'h08082828282828080808080808080808, /* 2128 */
128'h08080808080808080808080808080808, /* 2129 */
128'h101010101010101010101010101010a0, /* 2130 */
128'h10101010101004040404040404040404, /* 2131 */
128'h01010101010101010141414141414110, /* 2132 */
128'h10101010100101010101010101010101, /* 2133 */
128'h02020202020202020242424242424210, /* 2134 */
128'h08101010100202020202020202020202, /* 2135 */
128'h00000000000000000000000000000000, /* 2136 */
128'h00000000000000000000000000000000, /* 2137 */
128'h101010101010101010101010101010a0, /* 2138 */
128'h10101010101010101010101010101010, /* 2139 */
128'h01010101010101010101010101010101, /* 2140 */
128'h02010101010101011001010101010101, /* 2141 */
128'h02020202020202020202020202020202, /* 2142 */
128'h02020202020202021002020202020202, /* 2143 */
128'hc1bdceee242070dbe8c7b756d76aa478, /* 2144 */
128'hfd469501a83046134787c62af57c0faf, /* 2145 */
128'h895cd7beffff5bb18b44f7af698098d8, /* 2146 */
128'h49b40821a679438efd9871936b901122, /* 2147 */
128'he9b6c7aa265e5a51c040b340f61e2562, /* 2148 */
128'he7d3fbc8d8a1e68102441453d62f105d, /* 2149 */
128'h455a14edf4d50d87c33707d621e1cde6, /* 2150 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /* 2151 */
128'hfde5380c6d9d61228771f681fffa3942, /* 2152 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /* 2153 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /* 2154 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /* 2155 */
128'hfc93a039ab9423a7432aff97f4292244, /* 2156 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /* 2157 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /* 2158 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /* 2159 */
128'h0c07020d08030e09040f0a05000b0601, /* 2160 */
128'h020f0c090603000d0a0704010e0b0805, /* 2161 */
128'h09020b040d060f08010a030c050e0700, /* 2162 */
128'h6c5f7465735f64735f63736972776f6c, /* 2163 */
128'h6e67696c615f64730000000000006465, /* 2164 */
128'h645f6b6c635f64730000000000000000, /* 2165 */
128'h69747465735f64730000000000007669, /* 2166 */
128'h735f646d635f6473000000000000676e, /* 2167 */
128'h74657365725f64730000000074726174, /* 2168 */
128'h6e636b6c625f64730000000000000000, /* 2169 */
128'h69736b6c625f64730000000000000074, /* 2170 */
128'h6f656d69745f6473000000000000657a, /* 2171 */
128'h655f7172695f64730000000000007475, /* 2172 */
128'h5f63736972776f6c000000000000006e, /* 2173 */
128'h00000000646d635f74726174735f6473, /* 2174 */
128'h746e695f746961775f63736972776f6c, /* 2175 */
128'h000000000067616c665f747075727265, /* 2176 */
128'h00007172695f64735f63736972776f6c, /* 2177 */
128'h695f646d635f64735f63736972776f6c, /* 2178 */
128'h5f63736972776f6c0000000000007172, /* 2179 */
128'h007172695f646e655f617461645f6473, /* 2180 */
128'h0000000087fe88880000000087fe9f48, /* 2181 */
128'h004c4b40004c4b400030000020000000, /* 2182 */
128'h6d6d5f6472616f62000000020000ffff, /* 2183 */
128'h0000000087fe4e880064637465675f63, /* 2184 */
128'h0000000087fe4cf40000000087fe4a96, /* 2185 */
128'h00000000000000000000000000000000, /* 2186 */
128'hffffcf76ffffcf72ffffcf72ffffcf4c, /* 2187 */
128'hffffcf7affffcf7affffcf7affffcf7a, /* 2188 */
128'h0000000087fea2a00000000087fea290, /* 2189 */
128'h0000000087fea2c80000000087fea2b0, /* 2190 */
128'h0000000087fea2f80000000087fea2e0, /* 2191 */
128'h0000000087fea3280000000087fea310, /* 2192 */
128'h0000000087fea3580000000087fea340, /* 2193 */
128'h0000000087fea3880000000087fea370, /* 2194 */
128'h40040300400402004004010040040000, /* 2195 */
128'h40050000400405004004040140040400, /* 2196 */
128'h30000000000000030000000040050100, /* 2197 */
128'h60000000000000053000000000000001, /* 2198 */
128'h70000000000000027000000000000004, /* 2199 */
128'h00000001400000007000000000000000, /* 2200 */
128'h00000005000000012000000000000006, /* 2201 */
128'h20000000000000020000000040000000, /* 2202 */
128'h00000000100000000000000100000000, /* 2203 */
128'h1e19140f0d0c0a000000000000000000, /* 2204 */
128'h000186a00000271050463c37322d2823, /* 2205 */
128'h017d7840017d784000989680000f4240, /* 2206 */
128'h031975000319750002faf080018cba80, /* 2207 */
128'h02faf08005f5e10002faf080017d7840, /* 2208 */
128'h00000020000000000bebc2000c65d400, /* 2209 */
128'h00000200000001000000008000000040, /* 2210 */
128'h00002000000010000000080000000400, /* 2211 */
128'h0000c000000080000000600000004000, /* 2212 */
128'h37363534333231300002000000010000, /* 2213 */
128'h2043534952776f4c4645444342413938, /* 2214 */
128'h746f6f622d7520646573696d696e696d, /* 2215 */
128'h00000000647261432d445320726f6620, /* 2216 */
128'h3809000038000000100c0000edfe0dd0, /* 2217 */
128'h00000000100000001100000028000000, /* 2218 */
128'h000000000000000000090000d8020000, /* 2219 */
128'h00000000010000000000000000000000, /* 2220 */
128'h02000000000000000400000003000000, /* 2221 */
128'h020000000f0000000400000003000000, /* 2222 */
128'h2c6874651b0000001400000003000000, /* 2223 */
128'h007665642d657261622d656e61697261, /* 2224 */
128'h2c687465260000001000000003000000, /* 2225 */
128'h0100000000657261622d656e61697261, /* 2226 */
128'h1a0000000300000000006e65736f6863, /* 2227 */
128'h303140747261752f636f732f2c000000, /* 2228 */
128'h0000003030323531313a303030303030, /* 2229 */
128'h00000000737570630100000002000000, /* 2230 */
128'h01000000000000000400000003000000, /* 2231 */
128'h000000000f0000000400000003000000, /* 2232 */
128'h40787d01380000000400000003000000, /* 2233 */
128'h03000000000000304075706301000000, /* 2234 */
128'h0300000080f0fa024b00000004000000, /* 2235 */
128'h03000000007570635b00000004000000, /* 2236 */
128'h03000000000000006700000004000000, /* 2237 */
128'h0000000079616b6f6b00000005000000, /* 2238 */
128'h2c6874651b0000001200000003000000, /* 2239 */
128'h000000766373697200656e6169726120, /* 2240 */
128'h34367672720000000b00000003000000, /* 2241 */
128'h0b000000030000000000757363616d69, /* 2242 */
128'h0000393376732c76637369727c000000, /* 2243 */
128'h01000000850000000000000003000000, /* 2244 */
128'h6f72746e6f632d747075727265746e69, /* 2245 */
128'h04000000030000000000000072656c6c, /* 2246 */
128'h0000000003000000010000008f000000, /* 2247 */
128'h1b0000000f00000003000000a0000000, /* 2248 */
128'h000063746e692d7570632c7663736972, /* 2249 */
128'h02000000b50000000400000003000000, /* 2250 */
128'h02000000bb0000000400000003000000, /* 2251 */
128'h01000000020000000200000002000000, /* 2252 */
128'h0030303030303030384079726f6d656d, /* 2253 */
128'h6f6d656d5b0000000700000003000000, /* 2254 */
128'h67000000100000000300000000007972, /* 2255 */
128'h00000040000000000000008000000000, /* 2256 */
128'h000000007364656c0100000002000000, /* 2257 */
128'h6f6970671b0000000a00000003000000, /* 2258 */
128'h72616568010000000000007364656c2d, /* 2259 */
128'h0300000000000064656c2d7461656274, /* 2260 */
128'h0100000001000000c30000000c000000, /* 2261 */
128'hc90000000a0000000300000000000000, /* 2262 */
128'h03000000000000746165627472616568, /* 2263 */
128'h0200000002000000df00000000000000, /* 2264 */
128'h040000000300000000636f7301000000, /* 2265 */
128'h04000000030000000200000000000000, /* 2266 */
128'h1f00000003000000020000000f000000, /* 2267 */
128'h622d656e616972612c6874651b000000, /* 2268 */
128'h622d656c706d697300636f732d657261, /* 2269 */
128'hf6000000000000000300000000007375, /* 2270 */
128'h30303030303240746e696c6301000000, /* 2271 */
128'h1b0000000d0000000300000000000030, /* 2272 */
128'h0000000030746e696c632c7663736972, /* 2273 */
128'h02000000fd0000001000000003000000, /* 2274 */
128'h03000000070000000200000003000000, /* 2275 */
128'h00000002000000006700000010000000, /* 2276 */
128'h080000000300000000000c0000000000, /* 2277 */
128'h02000000006c6f72746e6f6311010000, /* 2278 */
128'h6f632d747075727265746e6901000000, /* 2279 */
128'h303030303030634072656c6c6f72746e, /* 2280 */
128'h00000000040000000300000000000000, /* 2281 */
128'h8f000000040000000300000000000000, /* 2282 */
128'h1b0000000c0000000300000001000000, /* 2283 */
128'h03000000003063696c702c7663736972, /* 2284 */
128'h1000000003000000a000000000000000, /* 2285 */
128'h020000000b00000002000000fd000000, /* 2286 */
128'h67000000100000000300000009000000, /* 2287 */
128'h00000004000000000000000c00000000, /* 2288 */
128'h070000001b0100000400000003000000, /* 2289 */
128'h030000002e0100000400000003000000, /* 2290 */
128'h03000000b50000000400000003000000, /* 2291 */
128'h03000000bb0000000400000003000000, /* 2292 */
128'h6f632d67756265640100000002000000, /* 2293 */
128'h030000000000304072656c6c6f72746e, /* 2294 */
128'h65642c76637369721b00000010000000, /* 2295 */
128'h0800000003000000003331302d677562, /* 2296 */
128'h03000000ffff000002000000fd000000, /* 2297 */
128'h00000000000000006700000010000000, /* 2298 */
128'h08000000030000000010000000000000, /* 2299 */
128'h02000000006c6f72746e6f6311010000, /* 2300 */
128'h30303030303031407472617501000000, /* 2301 */
128'h1b000000080000000300000000000030, /* 2302 */
128'h1000000003000000003035373631736e, /* 2303 */
128'h00000000000000100000000067000000, /* 2304 */
128'h4b000000040000000300000000100000, /* 2305 */
128'h39010000040000000300000080f0fa02, /* 2306 */
128'h47010000040000000300000000c20100, /* 2307 */
128'h58010000040000000300000003000000, /* 2308 */
128'h63010000040000000300000001000000, /* 2309 */
128'h6d010000040000000300000002000000, /* 2310 */
128'h2d737078010000000200000004000000, /* 2311 */
128'h00000000303030303030303240697073, /* 2312 */
128'h786e6c781b0000002800000003000000, /* 2313 */
128'h00622e30302e322d6970732d7370782c, /* 2314 */
128'h302e322d6970732d7370782c786e6c78, /* 2315 */
128'h00000000040000000300000000612e30, /* 2316 */
128'h0f000000040000000300000001000000, /* 2317 */
128'h47010000040000000300000000000000, /* 2318 */
128'h58010000080000000300000003000000, /* 2319 */
128'h10000000030000000200000002000000, /* 2320 */
128'h00000000000000200000000067000000, /* 2321 */
128'h7a010000080000000300000000100000, /* 2322 */
128'h040000000300000000377865746e696b, /* 2323 */
128'h04000000030000000100000086010000, /* 2324 */
128'h04000000030000000100000096010000, /* 2325 */
128'h040000000300000008000000a7010000, /* 2326 */
128'h40636d6d0100000004000000be010000, /* 2327 */
128'h1b0000000d0000000300000000000030, /* 2328 */
128'h00000000746f6c732d6970732d636d6d, /* 2329 */
128'h00000000670000000400000003000000, /* 2330 */
128'h20bcbe00cd0100000400000003000000, /* 2331 */
128'he40c0000df0100000800000003000000, /* 2332 */
128'hee0100000000000003000000e40c0000, /* 2333 */
128'h72776f6c010000000200000002000000, /* 2334 */
128'h3030303030303033406874652d637369, /* 2335 */
128'h1b0000000c0000000300000000000000, /* 2336 */
128'h03000000006874652d63736972776f6c, /* 2337 */
128'h006b726f7774656e5b00000008000000, /* 2338 */
128'h03000000470100000400000003000000, /* 2339 */
128'h03000000580100000800000003000000, /* 2340 */
128'hf9010000060000000300000000000000, /* 2341 */
128'h100000000300000000007fe3023e1800, /* 2342 */
128'h00000000000000300000000067000000, /* 2343 */
128'h6f697067010000000200000000800000, /* 2344 */
128'h03000000000000303030303030303440, /* 2345 */
128'h03000000020000000b02000004000000, /* 2346 */
128'h7370782c786e6c781b00000015000000, /* 2347 */
128'h00000000612e30302e312d6f6970672d, /* 2348 */
128'h03000000170200000000000003000000, /* 2349 */
128'h00000040000000006700000010000000, /* 2350 */
128'h04000000030000000000010000000000, /* 2351 */
128'h04000000030000000000000027020000, /* 2352 */
128'h04000000030000000000000037020000, /* 2353 */
128'h04000000030000000000000049020000, /* 2354 */
128'h0400000003000000000000005b020000, /* 2355 */
128'h0400000003000000080000006f020000, /* 2356 */
128'h0400000003000000080000007f020000, /* 2357 */
128'h04000000030000000000000090020000, /* 2358 */
128'h040000000300000001000000a7020000, /* 2359 */
128'h0400000003000000ffffffffb4020000, /* 2360 */
128'h0400000003000000ffffffffc5020000, /* 2361 */
128'h040000000300000001000000b5000000, /* 2362 */
128'h020000000200000001000000bb000000, /* 2363 */
128'h73736572646461230900000002000000, /* 2364 */
128'h6c65632d657a69732300736c6c65632d, /* 2365 */
128'h6f6d00656c62697461706d6f6300736c, /* 2366 */
128'h00687461702d74756f647473006c6564, /* 2367 */
128'h6e6575716572662d65736162656d6974, /* 2368 */
128'h6e6575716572662d6b636f6c63007963, /* 2369 */
128'h7200657079745f656369766564007963, /* 2370 */
128'h2c766373697200737574617473006765, /* 2371 */
128'h626c7400657079742d756d6d00617369, /* 2372 */
128'h7075727265746e69230074696c70732d, /* 2373 */
128'h7075727265746e6900736c6c65632d74, /* 2374 */
128'h6e696c0072656c6c6f72746e6f632d74, /* 2375 */
128'h736f69706700656c646e6168702c7875, /* 2376 */
128'h742d746c75616665642c78756e696c00, /* 2377 */
128'h74732d6e696174657200726567676972, /* 2378 */
128'h6172006465646e65707375732d657461, /* 2379 */
128'h2d73747075727265746e69007365676e, /* 2380 */
128'h6d616e2d676572006465646e65747865, /* 2381 */
128'h6972702d78616d2c7663736972007365, /* 2382 */
128'h7665646e2c766373697200797469726f, /* 2383 */
128'h690064656570732d746e657272756300, /* 2384 */
128'h00746e657261702d747075727265746e, /* 2385 */
128'h732d6765720073747075727265746e69, /* 2386 */
128'h746469772d6f692d6765720074666968, /* 2387 */
128'h6c7800796c696d61662c786e6c780068, /* 2388 */
128'h6c780074736978652d6f6669662c786e, /* 2389 */
128'h7800737469622d73732d6d756e2c786e, /* 2390 */
128'h726566736e6172742d6d756e2c786e6c, /* 2391 */
128'h722d6b63732c786e6c7800737469622d, /* 2392 */
128'h6572662d78616d2d697073006f697461, /* 2393 */
128'h722d656761746c6f760079636e657571, /* 2394 */
128'h70772d656c6261736964007365676e61, /* 2395 */
128'h65726464612d63616d2d6c61636f6c00, /* 2396 */
128'h6700736c6c65632d6f69706723007373, /* 2397 */
128'h780072656c6c6f72746e6f632d6f6970, /* 2398 */
128'h7800737475706e692d6c6c612c786e6c, /* 2399 */
128'h322d737475706e692d6c6c612c786e6c, /* 2400 */
128'h75616665642d74756f642c786e6c7800, /* 2401 */
128'h6665642d74756f642c786e6c7800746c, /* 2402 */
128'h6f6970672c786e6c7800322d746c7561, /* 2403 */
128'h6f6970672c786e6c780068746469772d, /* 2404 */
128'h746e692c786e6c780068746469772d32, /* 2405 */
128'h7800746e65736572702d747075727265, /* 2406 */
128'h786e6c78006c6175642d73692c786e6c, /* 2407 */
128'h6e6c7800746c75616665642d6972742c, /* 2408 */
128'h00322d746c75616665642d6972742c78, /* 2409 */
128'h0000000000203a642520656369766544, /* 2410 */
128'h00203a6425206563697665642073250a, /* 2411 */
128'h00000000203a6425206563697665440a, /* 2412 */
128'h000a656369766564206e776f6e6b6e75, /* 2413 */
128'h00000a2973252c73252870756b6f6f6c, /* 2414 */
128'h7265206c616e7265746e692070636864, /* 2415 */
128'h00000000000000000a7025202c726f72, /* 2416 */
128'h5145525f5043484420676e69646e6553, /* 2417 */
128'h4b434120504348440000000a54534555, /* 2418 */
128'h696c432050434844000000000000000a, /* 2419 */
128'h203a7373657264644120504920746e65, /* 2420 */
128'h0000000a64252e64252e64252e642520, /* 2421 */
128'h73657264644120504920726576726553, /* 2422 */
128'h0a64252e64252e64252e642520203a73, /* 2423 */
128'h6120726574756f520000000000000000, /* 2424 */
128'h252e64252e642520203a737365726464, /* 2425 */
128'h6b73616d2074654e0000000a64252e64, /* 2426 */
128'h64252e642520203a7373657264646120, /* 2427 */
128'h697420657361654c000a64252e64252e, /* 2428 */
128'h00000000000000000a6425203d20656d, /* 2429 */
128'h00000a22732522203d206e69616d6f64, /* 2430 */
128'h00000a22732522203d20726576726573, /* 2431 */
128'h000000000a44455050494b53204b4341, /* 2432 */
128'h000000000000000a4b414e2050434844, /* 2433 */
128'h73657264646120646574736575716552, /* 2434 */
128'h0000000000000a646573756665722073, /* 2435 */
128'h000000000000000a732520726f727245, /* 2436 */
128'h6e6f6974706f2064656c646e61686e75, /* 2437 */
128'h656c646e61686e55000000000a642520, /* 2438 */
128'h64252065646f63706f20504348442064, /* 2439 */
128'h20676e69646e6553000000000000000a, /* 2440 */
128'h000a595245564f435349445f50434844, /* 2441 */
128'h00000000000a29732528726f72726570, /* 2442 */
128'h3a2043414d2073250000000030687465, /* 2443 */
128'h3a583230253a583230253a5832302520, /* 2444 */
128'h000a583230253a583230253a58323025, /* 2445 */
128'h484420646e65732074276e646c756f43, /* 2446 */
128'h206e6f20595245564f43534944205043, /* 2447 */
128'h00000a7325203a732520656369766564, /* 2448 */
128'h5043484420726f6620676e6974696157, /* 2449 */
128'h2020202020202020000a524546464f5f, /* 2450 */
128'h00000000000063250000000000000020, /* 2451 */
128'h0000000000202020000000000000002e, /* 2452 */
128'h0000000000000a0a0000005832302520, /* 2453 */
128'h3a646c697542202c0000000073257325, /* 2454 */
128'h00000000000073250000000000732520, /* 2455 */
128'h000000000000000073257a4820756c25, /* 2456 */
128'h00000000646c252e0000000000756c25, /* 2457 */
128'h6574794220756c250073257a48632520, /* 2458 */
128'h00732542696325200000000000732573, /* 2459 */
128'h00786c6c2a30252000003a786c383025, /* 2460 */
128'h5b6e6f6974636553000a732520202020, /* 2461 */
128'h75716572206e656c000000203a5d6425, /* 2462 */
128'h6175746361202c5825203d2064657269, /* 2463 */
128'h25287970636d656d000a7825203d206c, /* 2464 */
128'h00000a3b29782578302c782578302c78, /* 2465 */
128'h782578302c302c7825287465736d656d, /* 2466 */
128'h464f5f4f4c43414d00000000000a3b29, /* 2467 */
128'h464f5f494843414d0000000054455346, /* 2468 */
128'h46464f5f524c50540000000054455346, /* 2469 */
128'h46464f5f534346540000000000544553, /* 2470 */
128'h4c5254434f49444d0000000000544553, /* 2471 */
128'h46464f5f534346520054455346464f5f, /* 2472 */
128'h5346464f5f5253520000000000544553, /* 2473 */
128'h46464f5f444142520000000000005445, /* 2474 */
128'h46464f5f524c50520000000000544553, /* 2475 */
128'h000000003f3f3f3f0000000000544553, /* 2476 */
128'h000064252b54455346464f5f524c5052, /* 2477 */
128'h6f746f72502050490000000000000047, /* 2478 */
128'h00000000000000000a50495049203d20, /* 2479 */
128'h6f746f72502050490000000000000054, /* 2480 */
128'h6f746f7250205049000a504745203d20, /* 2481 */
128'h6165682074736574000a505550203d20, /* 2482 */
128'h6e6f6320747365740000000a3a726564, /* 2483 */
128'h6f746f7250205049000a3a73746e6574, /* 2484 */
128'h6f746f7250205049000a504449203d20, /* 2485 */
128'h6f746f725020504900000a5054203d20, /* 2486 */
128'h00000000000000000a50434344203d20, /* 2487 */
128'h6f746f72502050490000000000000036, /* 2488 */
128'h00000000000000000a50565352203d20, /* 2489 */
128'h000a455247203d206f746f7250205049, /* 2490 */
128'h000a505345203d206f746f7250205049, /* 2491 */
128'h00000a4841203d206f746f7250205049, /* 2492 */
128'h000a50544d203d206f746f7250205049, /* 2493 */
128'h5054454542203d206f746f7250205049, /* 2494 */
128'h6f746f72502050490000000000000a48, /* 2495 */
128'h000000000000000a5041434e45203d20, /* 2496 */
128'h6f746f7250205049000000000000004d, /* 2497 */
128'h00000000000000000a504d4f43203d20, /* 2498 */
128'h0a50544353203d206f746f7250205049, /* 2499 */
128'h6f746f72502050490000000000000000, /* 2500 */
128'h00000000000a4554494c504455203d20, /* 2501 */
128'h0a534c504d203d206f746f7250205049, /* 2502 */
128'h6f746f72502050490000000000000000, /* 2503 */
128'h6f746f7270205049000a574152203d20, /* 2504 */
128'h2820646574726f707075736e75203d20, /* 2505 */
128'h79745f6f746f7270000000000a297825, /* 2506 */
128'h0000000000000a78257830203d206570, /* 2507 */
128'h727265746e692064656c646e61686e75, /* 2508 */
128'h414d2070757465530000000a21747075, /* 2509 */
128'h6c25203d2043414d000a726464612043, /* 2510 */
128'h726464612043414d00000a786c253a78, /* 2511 */
128'h3a783230253a78323025203d20737365, /* 2512 */
128'h253a783230253a783230253a78323025, /* 2513 */
128'h74656e72656874450000000a2e783230, /* 2514 */
128'h757461747320747075727265746e6920, /* 2515 */
128'h00000000000000000a646c25203d2073, /* 2516 */
128'h20646564616f6c2065687420746f6f42, /* 2517 */
128'h00000000000a2e2e2e6d6172676f7270, /* 2518 */
128'h207265746f6f62202c657962646f6f47, /* 2519 */
128'h3d3c3b3a2c2b2a22000000000a2e2e2e, /* 2520 */
128'h3c3b3a2e2c2b2a2200007f7c5d5b3f3e, /* 2521 */
128'h3736353433323130007f7c5d5b3f3e3d, /* 2522 */
128'h00000000000000006665646362613938, /* 2523 */
128'h2e636d6d5f63736972776f6c2f637273, /* 2524 */
128'h20657361625f64730000000000000063, /* 2525 */
128'h00726464615f657361625f6473203d3d, /* 2526 */
128'h74207325203a64735f63736972776f6c, /* 2527 */
128'h6d65722064726143000a74756f656d69, /* 2528 */
128'h676e616863206b73616d202c6465766f, /* 2529 */
128'h000000000000000a6425206f74206465, /* 2530 */
128'h6d202c6465747265736e692064726143, /* 2531 */
128'h25206f74206465676e616863206b7361, /* 2532 */
128'h6165726320636d6d0000000000000a64, /* 2533 */
128'h2074736f68202c782520746120646574, /* 2534 */
128'h00000000007365590000000a7825203d, /* 2535 */
128'h00000000524444200000000000006f4e, /* 2536 */
128'h203a656369766544002020203a434d4d, /* 2537 */
128'h74636166756e614d00000000000a7325, /* 2538 */
128'h000000000a7825203a44492072657275, /* 2539 */
128'h00000000000000000a7825203a4d454f, /* 2540 */
128'h63256325632563256325203a656d614e, /* 2541 */
128'h65657053207375420000000000000a20, /* 2542 */
128'h706143206867694800000a6425203a64, /* 2543 */
128'h0000000000000a7325203a7974696361, /* 2544 */
128'h000000000000203a7974696361706143, /* 2545 */
128'h69622d6425203a687464695720737542, /* 2546 */
128'h000000203a78250a000000000a732574, /* 2547 */
128'h5f63736972776f6c0000007825782520, /* 2548 */
128'h6f57206f6c6c65480000000000006473, /* 2549 */
128'h732068637469775300000a0d21646c72, /* 2550 */
128'h000000000a5825203d20676e69747465, /* 2551 */
128'h206e776f6e6b6e5500000a0d70617274, /* 2552 */
128'h45207375746174530000000065646f6d, /* 2553 */
128'h0000000a583830257830203a726f7272, /* 2554 */
128'h20676e69746961772074756f656d6954, /* 2555 */
128'h00000000000a79646165722064726163, /* 2556 */
128'h646e6573206f74206c69616620636d6d, /* 2557 */
128'h0000000000000a646d6320706f747320, /* 2558 */
128'h65626d756e206b636f6c62203a434d4d, /* 2559 */
128'h207364656563786520786c2578302072, /* 2560 */
128'h00000000000a29786c2578302878616d, /* 2561 */
128'h7571657220342e34203d3e20434d4d65, /* 2562 */
128'h65636e61686e6520726f662064657269, /* 2563 */
128'h61657261206174616420726573752064, /* 2564 */
128'h656f642064726143000000000000000a, /* 2565 */
128'h61702074726f7070757320746f6e2073, /* 2566 */
128'h00000000000a676e696e6f6974697472, /* 2567 */
128'h656420746f6e2073656f642064726143, /* 2568 */
128'h70756f726720505720434820656e6966, /* 2569 */
128'h746164207265735500000a657a697320, /* 2570 */
128'h2061657261206465636e61686e652061, /* 2571 */
128'h2070756f726720505720434820746f6e, /* 2572 */
128'h0000000a64656e67696c6120657a6973, /* 2573 */
128'h6e206e6f697469747261702069255047, /* 2574 */
128'h732070756f726720505720434820746f, /* 2575 */
128'h000000000a64656e67696c6120657a69, /* 2576 */
128'h757320746f6e2073656f642064726143, /* 2577 */
128'h61206465636e61686e652074726f7070, /* 2578 */
128'h000000000000000a6574756269727474, /* 2579 */
128'h73206465636e61686e65206c61746f54, /* 2580 */
128'h6978616d207364656563786520657a69, /* 2581 */
128'h00000a297525203e20752528206d756d, /* 2582 */
128'h757320746f6e2073656f642064726143, /* 2583 */
128'h72746e6f632074736f682074726f7070, /* 2584 */
128'h206e6f697469747261702064656c6c6f, /* 2585 */
128'h74696c696261696c6572206574697277, /* 2586 */
128'h00000000000a73676e69747465732079, /* 2587 */
128'h7261702079646165726c612064726143, /* 2588 */
128'h000000000000000a64656e6f69746974, /* 2589 */
128'h6572702064726163206f6e203a434d4d, /* 2590 */
128'h64696420647261430000000a746e6573, /* 2591 */
128'h206f7420646e6f7073657220746f6e20, /* 2592 */
128'h0a217463656c657320656761746c6f76, /* 2593 */
128'h7420656c62616e750000000000000000, /* 2594 */
128'h0a65646f6d2061207463656c6573206f, /* 2595 */
128'h635f747865206f4e0000000000000000, /* 2596 */
128'h0000000000000a21646e756f66206473, /* 2597 */
128'h34302520726e532078363025206e614d, /* 2598 */
128'h63256325632563250000007834302578, /* 2599 */
128'h00000064252e64250000000063256325, /* 2600 */
128'h00000000000079636167656c20434d4d, /* 2601 */
128'h0000000000000079636167654c204453, /* 2602 */
128'h28206465657053206867694820434d4d, /* 2603 */
128'h20686769482044530000297a484d3632, /* 2604 */
128'h000000297a484d303528206465657053, /* 2605 */
128'h28206465657053206867694820434d4d, /* 2606 */
128'h3552444420434d4d0000297a484d3235, /* 2607 */
128'h00000000000000297a484d3235282032, /* 2608 */
128'h7a484d35322820323152445320534855, /* 2609 */
128'h32524453205348550000000000000029, /* 2610 */
128'h00000000000000297a484d3035282035, /* 2611 */
128'h484d3030312820303552445320534855, /* 2612 */
128'h3552444420534855000000000000297a, /* 2613 */
128'h00000000000000297a484d3035282030, /* 2614 */
128'h4d383032282034303152445320534855, /* 2615 */
128'h32282030303253480000000000297a48, /* 2616 */
128'h6976654420434d4d0000297a484d3030, /* 2617 */
128'h0a646e756f6620746f6e206425206563, /* 2618 */
128'h00000000434d4d650000000000000000, /* 2619 */
128'h00006425203a73250000000000004453, /* 2620 */
128'h0000000000636d6d0000002973252820, /* 2621 */
128'h6425203d206874676e656c20656c6946, /* 2622 */
128'h2074736575716552000000000000000a, /* 2623 */
128'h25202e676e6f6c206f6f742068746170, /* 2624 */
128'h000000000000002f00000000000a646c, /* 2625 */
128'h6b636f6c62202c22732522203a717277, /* 2626 */
128'h00000000000000000a64253d657a6973, /* 2627 */
128'h646e6520656c69662065766965636552, /* 2628 */
128'h775f656c646e61680000000000000a2e, /* 2629 */
128'h00000000000a2e64656c6c6163207172, /* 2630 */
128'h65706f2050544654206c6167656c6c49, /* 2631 */
128'h00000000000000000a2e6e6f69746172, /* 2632 */
128'h445320746e756f6d206f74206c696146, /* 2633 */
128'h000000000000000a2172657669726420, /* 2634 */
128'h6e69206e69622e746f6f622064616f4c, /* 2635 */
128'h0000000000000a79726f6d656d206f74, /* 2636 */
128'h00000000000000006e69622e746f6f62, /* 2637 */
128'h62206e65706f206f742064656c696146, /* 2638 */
128'h206f74206c6961660000000a21746f6f, /* 2639 */
128'h000000000021656c69662065736f6c63, /* 2640 */
128'h6420746e756f6d75206f74206c696166, /* 2641 */
128'h2520646564616f4c00000000216b7369, /* 2642 */
128'h726f6d656d206f742073657479622064, /* 2643 */
128'h6f726620782520737365726464612079, /* 2644 */
128'h642520666f206e69622e746f6f62206d, /* 2645 */
128'h00000000000000000a2e736574796220, /* 2646 */
128'h20524444206f7420666c652064616f6c, /* 2647 */
128'h6461657220666c65000a79726f6d656d, /* 2648 */
128'h646f6320687469772064656c69616620, /* 2649 */
128'h000000005c2d2f7c0000000064252065, /* 2650 */
128'h696620646573616220746f6f622d750a, /* 2651 */
128'h6c20746f6f6220656761747320747372, /* 2652 */
128'h6f6974726573736100000a726564616f, /* 2653 */
128'h6c6966202c64656c696166207325206e, /* 2654 */
128'h66202c642520656e696c202c73252065, /* 2655 */
128'h00000000000a7325206e6f6974636e75, /* 2656 */
128'hefcdab8967452301cccccccccccccccd, /* 2657 */
128'h10000000200000001032547698badcfe, /* 2658 */
128'h00000000000000005851f42d4c957f2d, /* 2659 */
128'h00000000000000000000000000000000, /* 2660 */
128'h00000000000000000000000000000000, /* 2661 */
128'h00000000000000000000000000000000, /* 2662 */
128'h00000000000000000000000000000000, /* 2663 */
128'h00000000000000000000000000000000, /* 2664 */
128'h00000000000000000000000000000000, /* 2665 */
128'h00000000000000000000000000000000, /* 2666 */
128'h00000000000000000000000000000000, /* 2667 */
128'h00000000000000000000000000000000, /* 2668 */
128'h00000000000000000000000000000000, /* 2669 */
128'h00000000000000000000000000000000, /* 2670 */
128'h00000000000000000000000000000000, /* 2671 */
128'h00004b4d47545045000000030f060301, /* 2672 */
128'h000000003000000000000000004b4d47, /* 2673 */
128'h00000000ffffffff0000000000000000, /* 2674 */
128'h0000646d635f6473000000000c000000, /* 2675 */
128'h00000000ffffffff00006772615f6473, /* 2676 */
128'h0000000087fea3d80000000087fea220, /* 2677 */
128'h0000000000000000ffffffff00000006, /* 2678 */
128'h0000000000000000000000000000008c, /* 2679 */
128'h00000000000000000000000000000000, /* 2680 */
128'h00000000000000000000000000000000, /* 2681 */
128'h00000000000000000000000000000000, /* 2682 */
128'h00000000000000000000000000000000, /* 2683 */
128'h00000000000000000000000000000000, /* 2684 */
128'h00000000000000000000000000000000, /* 2685 */
128'h00000000000000000000000000000000, /* 2686 */
128'h00000000000000000000000000000000, /* 2687 */
128'h00000000000000000000000000000000, /* 2688 */
128'h00000000000000000000000000000000, /* 2689 */
128'h00000000000000000000000000000000, /* 2690 */
128'h00000000000000000000000000000000, /* 2691 */
128'h00000000000000000000000000000000, /* 2692 */
128'h00000000000000000000000000000000, /* 2693 */
128'h00000000000000000000000000000000, /* 2694 */
128'h00000000000000000000000000000000, /* 2695 */
128'h00000000000000000000000000000000, /* 2696 */
128'h00000000000000000000000000000000, /* 2697 */
128'h00000000000000000000000000000000, /* 2698 */
128'h00000000000000000000000000000000, /* 2699 */
128'h00000000000000000000000000000000, /* 2700 */
128'h00000000000000000000000000000000, /* 2701 */
128'h00000000000000000000000000000000, /* 2702 */
128'h00000000000000000000000000000000, /* 2703 */
128'h00000000000000000000000000000000, /* 2704 */
128'h00000000000000000000000000000000, /* 2705 */
128'h00000000000000000000000000000000, /* 2706 */
128'h00000000000000000000000000000000, /* 2707 */
128'h00000000000000000000000000000000, /* 2708 */
128'h00000000000000000000000000000000, /* 2709 */
128'h00000000000000000000000000000000, /* 2710 */
128'h00000000000000000000000000000000, /* 2711 */
128'h00000000000000000000000000000000, /* 2712 */
128'h00000000000000000000000000000000, /* 2713 */
128'h00000000000000000000000000000000, /* 2714 */
128'h00000000000000000000000000000000, /* 2715 */
128'h00000000000000000000000000000000, /* 2716 */
128'h00000000000000000000000000000000, /* 2717 */
128'h00000000000000000000000000000000, /* 2718 */
128'h00000000000000000000000000000000, /* 2719 */
128'h00000000000000000000000000000000, /* 2720 */
128'h00000000000000000000000000000000, /* 2721 */
128'h00000000000000000000000000000000, /* 2722 */
128'h00000000000000000000000000000000, /* 2723 */
128'h00000000000000000000000000000000, /* 2724 */
128'h00000000000000000000000000000000, /* 2725 */
128'h00000000000000000000000000000000, /* 2726 */
128'h00000000000000000000000000000000, /* 2727 */
128'h00000000000000000000000000000000, /* 2728 */
128'h00000000000000000000000000000000, /* 2729 */
128'h00000000000000000000000000000000, /* 2730 */
128'h00000000000000000000000000000000, /* 2731 */
128'h00000000000000000000000000000000, /* 2732 */
128'h00000000000000000000000000000000, /* 2733 */
128'h00000000000000000000000000000000, /* 2734 */
128'h00000000000000000000000000000000, /* 2735 */
128'h00000000000000000000000000000000, /* 2736 */
128'h00000000000000000000000000000000, /* 2737 */
128'h00000000000000000000000000000000, /* 2738 */
128'h00000000000000000000000000000000, /* 2739 */
128'h00000000000000000000000000000000, /* 2740 */
128'h00000000000000000000000000000000, /* 2741 */
128'h00000000000000000000000000000000, /* 2742 */
128'h00000000000000000000000000000000, /* 2743 */
128'h00000000000000000000000000000000, /* 2744 */
128'h00000000000000000000000000000000, /* 2745 */
128'h00000000000000000000000000000000, /* 2746 */
128'h00000000000000000000000000000000, /* 2747 */
128'h00000000000000000000000000000000, /* 2748 */
128'h00000000000000000000000000000000, /* 2749 */
128'h00000000000000000000000000000000, /* 2750 */
128'h00000000000000000000000000000000, /* 2751 */
128'h00000000000000000000000000000000, /* 2752 */
128'h00000000000000000000000000000000, /* 2753 */
128'h00000000000000000000000000000000, /* 2754 */
128'h00000000000000000000000000000000, /* 2755 */
128'h00000000000000000000000000000000, /* 2756 */
128'h00000000000000000000000000000000, /* 2757 */
128'h00000000000000000000000000000000, /* 2758 */
128'h00000000000000000000000000000000, /* 2759 */
128'h00000000000000000000000000000000, /* 2760 */
128'h00000000000000000000000000000000, /* 2761 */
128'h00000000000000000000000000000000, /* 2762 */
128'h00000000000000000000000000000000, /* 2763 */
128'h00000000000000000000000000000000, /* 2764 */
128'h00000000000000000000000000000000, /* 2765 */
128'h00000000000000000000000000000000, /* 2766 */
128'h00000000000000000000000000000000, /* 2767 */
128'h00000000000000000000000000000000, /* 2768 */
128'h00000000000000000000000000000000, /* 2769 */
128'h00000000000000000000000000000000, /* 2770 */
128'h00000000000000000000000000000000, /* 2771 */
128'h00000000000000000000000000000000, /* 2772 */
128'h00000000000000000000000000000000, /* 2773 */
128'h00000000000000000000000000000000, /* 2774 */
128'h00000000000000000000000000000000, /* 2775 */
128'h00000000000000000000000000000000, /* 2776 */
128'h00000000000000000000000000000000, /* 2777 */
128'h00000000000000000000000000000000, /* 2778 */
128'h00000000000000000000000000000000, /* 2779 */
128'h00000000000000000000000000000000, /* 2780 */
128'h00000000000000000000000000000000, /* 2781 */
128'h00000000000000000000000000000000, /* 2782 */
128'h00000000000000000000000000000000, /* 2783 */
128'h00000000000000000000000000000000, /* 2784 */
128'h00000000000000000000000000000000, /* 2785 */
128'h00000000000000000000000000000000, /* 2786 */
128'h00000000000000000000000000000000, /* 2787 */
128'h00000000000000000000000000000000, /* 2788 */
128'h00000000000000000000000000000000, /* 2789 */
128'h00000000000000000000000000000000, /* 2790 */
128'h00000000000000000000000000000000, /* 2791 */
128'h00000000000000000000000000000000, /* 2792 */
128'h00000000000000000000000000000000, /* 2793 */
128'h00000000000000000000000000000000, /* 2794 */
128'h00000000000000000000000000000000, /* 2795 */
128'h00000000000000000000000000000000, /* 2796 */
128'h00000000000000000000000000000000, /* 2797 */
128'h00000000000000000000000000000000, /* 2798 */
128'h00000000000000000000000000000000, /* 2799 */
128'h00000000000000000000000000000000, /* 2800 */
128'h00000000000000000000000000000000, /* 2801 */
128'h00000000000000000000000000000000, /* 2802 */
128'h00000000000000000000000000000000, /* 2803 */
128'h00000000000000000000000000000000, /* 2804 */
128'h00000000000000000000000000000000, /* 2805 */
128'h00000000000000000000000000000000, /* 2806 */
128'h00000000000000000000000000000000, /* 2807 */
128'h00000000000000000000000000000000, /* 2808 */
128'h00000000000000000000000000000000, /* 2809 */
128'h00000000000000000000000000000000, /* 2810 */
128'h00000000000000000000000000000000, /* 2811 */
128'h00000000000000000000000000000000, /* 2812 */
128'h00000000000000000000000000000000, /* 2813 */
128'h00000000000000000000000000000000, /* 2814 */
128'h00000000000000000000000000000000, /* 2815 */
128'h00000000000000000000000000000000, /* 2816 */
128'h00000000000000000000000000000000, /* 2817 */
128'h00000000000000000000000000000000, /* 2818 */
128'h00000000000000000000000000000000, /* 2819 */
128'h00000000000000000000000000000000, /* 2820 */
128'h00000000000000000000000000000000, /* 2821 */
128'h00000000000000000000000000000000, /* 2822 */
128'h00000000000000000000000000000000, /* 2823 */
128'h00000000000000000000000000000000, /* 2824 */
128'h00000000000000000000000000000000, /* 2825 */
128'h00000000000000000000000000000000, /* 2826 */
128'h00000000000000000000000000000000, /* 2827 */
128'h00000000000000000000000000000000, /* 2828 */
128'h00000000000000000000000000000000, /* 2829 */
128'h00000000000000000000000000000000, /* 2830 */
128'h00000000000000000000000000000000, /* 2831 */
128'h00000000000000000000000000000000, /* 2832 */
128'h00000000000000000000000000000000, /* 2833 */
128'h00000000000000000000000000000000, /* 2834 */
128'h00000000000000000000000000000000, /* 2835 */
128'h00000000000000000000000000000000, /* 2836 */
128'h00000000000000000000000000000000, /* 2837 */
128'h00000000000000000000000000000000, /* 2838 */
128'h00000000000000000000000000000000, /* 2839 */
128'h00000000000000000000000000000000, /* 2840 */
128'h00000000000000000000000000000000, /* 2841 */
128'h00000000000000000000000000000000, /* 2842 */
128'h00000000000000000000000000000000, /* 2843 */
128'h00000000000000000000000000000000, /* 2844 */
128'h00000000000000000000000000000000, /* 2845 */
128'h00000000000000000000000000000000, /* 2846 */
128'h00000000000000000000000000000000, /* 2847 */
128'h00000000000000000000000000000000, /* 2848 */
128'h00000000000000000000000000000000, /* 2849 */
128'h00000000000000000000000000000000, /* 2850 */
128'h00000000000000000000000000000000, /* 2851 */
128'h00000000000000000000000000000000, /* 2852 */
128'h00000000000000000000000000000000, /* 2853 */
128'h00000000000000000000000000000000, /* 2854 */
128'h00000000000000000000000000000000, /* 2855 */
128'h00000000000000000000000000000000, /* 2856 */
128'h00000000000000000000000000000000, /* 2857 */
128'h00000000000000000000000000000000, /* 2858 */
128'h00000000000000000000000000000000, /* 2859 */
128'h00000000000000000000000000000000, /* 2860 */
128'h00000000000000000000000000000000, /* 2861 */
128'h00000000000000000000000000000000, /* 2862 */
128'h00000000000000000000000000000000, /* 2863 */
128'h00000000000000000000000000000000, /* 2864 */
128'h00000000000000000000000000000000, /* 2865 */
128'h00000000000000000000000000000000, /* 2866 */
128'h00000000000000000000000000000000, /* 2867 */
128'h00000000000000000000000000000000, /* 2868 */
128'h00000000000000000000000000000000, /* 2869 */
128'h00000000000000000000000000000000, /* 2870 */
128'h00000000000000000000000000000000, /* 2871 */
128'h00000000000000000000000000000000, /* 2872 */
128'h00000000000000000000000000000000, /* 2873 */
128'h00000000000000000000000000000000, /* 2874 */
128'h00000000000000000000000000000000, /* 2875 */
128'h00000000000000000000000000000000, /* 2876 */
128'h00000000000000000000000000000000, /* 2877 */
128'h00000000000000000000000000000000, /* 2878 */
128'h00000000000000000000000000000000, /* 2879 */
128'h00000000000000000000000000000000, /* 2880 */
128'h00000000000000000000000000000000, /* 2881 */
128'h00000000000000000000000000000000, /* 2882 */
128'h00000000000000000000000000000000, /* 2883 */
128'h00000000000000000000000000000000, /* 2884 */
128'h00000000000000000000000000000000, /* 2885 */
128'h00000000000000000000000000000000, /* 2886 */
128'h00000000000000000000000000000000, /* 2887 */
128'h00000000000000000000000000000000, /* 2888 */
128'h00000000000000000000000000000000, /* 2889 */
128'h00000000000000000000000000000000, /* 2890 */
128'h00000000000000000000000000000000, /* 2891 */
128'h00000000000000000000000000000000, /* 2892 */
128'h00000000000000000000000000000000, /* 2893 */
128'h00000000000000000000000000000000, /* 2894 */
128'h00000000000000000000000000000000, /* 2895 */
128'h00000000000000000000000000000000, /* 2896 */
128'h00000000000000000000000000000000, /* 2897 */
128'h00000000000000000000000000000000, /* 2898 */
128'h00000000000000000000000000000000, /* 2899 */
128'h00000000000000000000000000000000, /* 2900 */
128'h00000000000000000000000000000000, /* 2901 */
128'h00000000000000000000000000000000, /* 2902 */
128'h00000000000000000000000000000000, /* 2903 */
128'h00000000000000000000000000000000, /* 2904 */
128'h00000000000000000000000000000000, /* 2905 */
128'h00000000000000000000000000000000, /* 2906 */
128'h00000000000000000000000000000000, /* 2907 */
128'h00000000000000000000000000000000, /* 2908 */
128'h00000000000000000000000000000000, /* 2909 */
128'h00000000000000000000000000000000, /* 2910 */
128'h00000000000000000000000000000000, /* 2911 */
128'h00000000000000000000000000000000, /* 2912 */
128'h00000000000000000000000000000000, /* 2913 */
128'h00000000000000000000000000000000, /* 2914 */
128'h00000000000000000000000000000000, /* 2915 */
128'h00000000000000000000000000000000, /* 2916 */
128'h00000000000000000000000000000000, /* 2917 */
128'h00000000000000000000000000000000, /* 2918 */
128'h00000000000000000000000000000000, /* 2919 */
128'h00000000000000000000000000000000, /* 2920 */
128'h00000000000000000000000000000000, /* 2921 */
128'h00000000000000000000000000000000, /* 2922 */
128'h00000000000000000000000000000000, /* 2923 */
128'h00000000000000000000000000000000, /* 2924 */
128'h00000000000000000000000000000000, /* 2925 */
128'h00000000000000000000000000000000, /* 2926 */
128'h00000000000000000000000000000000, /* 2927 */
128'h00000000000000000000000000000000, /* 2928 */
128'h00000000000000000000000000000000, /* 2929 */
128'h00000000000000000000000000000000, /* 2930 */
128'h00000000000000000000000000000000, /* 2931 */
128'h00000000000000000000000000000000, /* 2932 */
128'h00000000000000000000000000000000, /* 2933 */
128'h00000000000000000000000000000000, /* 2934 */
128'h00000000000000000000000000000000, /* 2935 */
128'h00000000000000000000000000000000, /* 2936 */
128'h00000000000000000000000000000000, /* 2937 */
128'h00000000000000000000000000000000, /* 2938 */
128'h00000000000000000000000000000000, /* 2939 */
128'h00000000000000000000000000000000, /* 2940 */
128'h00000000000000000000000000000000, /* 2941 */
128'h00000000000000000000000000000000, /* 2942 */
128'h00000000000000000000000000000000, /* 2943 */
128'h00000000000000000000000000000000, /* 2944 */
128'h00000000000000000000000000000000, /* 2945 */
128'h00000000000000000000000000000000, /* 2946 */
128'h00000000000000000000000000000000, /* 2947 */
128'h00000000000000000000000000000000, /* 2948 */
128'h00000000000000000000000000000000, /* 2949 */
128'h00000000000000000000000000000000, /* 2950 */
128'h00000000000000000000000000000000, /* 2951 */
128'h00000000000000000000000000000000, /* 2952 */
128'h00000000000000000000000000000000, /* 2953 */
128'h00000000000000000000000000000000, /* 2954 */
128'h00000000000000000000000000000000, /* 2955 */
128'h00000000000000000000000000000000, /* 2956 */
128'h00000000000000000000000000000000, /* 2957 */
128'h00000000000000000000000000000000, /* 2958 */
128'h00000000000000000000000000000000, /* 2959 */
128'h00000000000000000000000000000000, /* 2960 */
128'h00000000000000000000000000000000, /* 2961 */
128'h00000000000000000000000000000000, /* 2962 */
128'h00000000000000000000000000000000, /* 2963 */
128'h00000000000000000000000000000000, /* 2964 */
128'h00000000000000000000000000000000, /* 2965 */
128'h00000000000000000000000000000000, /* 2966 */
128'h00000000000000000000000000000000, /* 2967 */
128'h00000000000000000000000000000000, /* 2968 */
128'h00000000000000000000000000000000, /* 2969 */
128'h00000000000000000000000000000000, /* 2970 */
128'h00000000000000000000000000000000, /* 2971 */
128'h00000000000000000000000000000000, /* 2972 */
128'h00000000000000000000000000000000, /* 2973 */
128'h00000000000000000000000000000000, /* 2974 */
128'h00000000000000000000000000000000, /* 2975 */
128'h00000000000000000000000000000000, /* 2976 */
128'h00000000000000000000000000000000, /* 2977 */
128'h00000000000000000000000000000000, /* 2978 */
128'h00000000000000000000000000000000, /* 2979 */
128'h00000000000000000000000000000000, /* 2980 */
128'h00000000000000000000000000000000, /* 2981 */
128'h00000000000000000000000000000000, /* 2982 */
128'h00000000000000000000000000000000, /* 2983 */
128'h00000000000000000000000000000000, /* 2984 */
128'h00000000000000000000000000000000, /* 2985 */
128'h00000000000000000000000000000000, /* 2986 */
128'h00000000000000000000000000000000, /* 2987 */
128'h00000000000000000000000000000000, /* 2988 */
128'h00000000000000000000000000000000, /* 2989 */
128'h00000000000000000000000000000000, /* 2990 */
128'h00000000000000000000000000000000, /* 2991 */
128'h00000000000000000000000000000000, /* 2992 */
128'h00000000000000000000000000000000, /* 2993 */
128'h00000000000000000000000000000000, /* 2994 */
128'h00000000000000000000000000000000, /* 2995 */
128'h00000000000000000000000000000000, /* 2996 */
128'h00000000000000000000000000000000, /* 2997 */
128'h00000000000000000000000000000000, /* 2998 */
128'h00000000000000000000000000000000, /* 2999 */
128'h00000000000000000000000000000000, /* 3000 */
128'h00000000000000000000000000000000, /* 3001 */
128'h00000000000000000000000000000000, /* 3002 */
128'h00000000000000000000000000000000, /* 3003 */
128'h00000000000000000000000000000000, /* 3004 */
128'h00000000000000000000000000000000, /* 3005 */
128'h00000000000000000000000000000000, /* 3006 */
128'h00000000000000000000000000000000, /* 3007 */
128'h00000000000000000000000000000000, /* 3008 */
128'h00000000000000000000000000000000, /* 3009 */
128'h00000000000000000000000000000000, /* 3010 */
128'h00000000000000000000000000000000, /* 3011 */
128'h00000000000000000000000000000000, /* 3012 */
128'h00000000000000000000000000000000, /* 3013 */
128'h00000000000000000000000000000000, /* 3014 */
128'h00000000000000000000000000000000, /* 3015 */
128'h00000000000000000000000000000000, /* 3016 */
128'h00000000000000000000000000000000, /* 3017 */
128'h00000000000000000000000000000000, /* 3018 */
128'h00000000000000000000000000000000, /* 3019 */
128'h00000000000000000000000000000000, /* 3020 */
128'h00000000000000000000000000000000, /* 3021 */
128'h00000000000000000000000000000000, /* 3022 */
128'h00000000000000000000000000000000, /* 3023 */
128'h00000000000000000000000000000000, /* 3024 */
128'h00000000000000000000000000000000, /* 3025 */
128'h00000000000000000000000000000000, /* 3026 */
128'h00000000000000000000000000000000, /* 3027 */
128'h00000000000000000000000000000000, /* 3028 */
128'h00000000000000000000000000000000, /* 3029 */
128'h00000000000000000000000000000000, /* 3030 */
128'h00000000000000000000000000000000, /* 3031 */
128'h00000000000000000000000000000000, /* 3032 */
128'h00000000000000000000000000000000, /* 3033 */
128'h00000000000000000000000000000000, /* 3034 */
128'h00000000000000000000000000000000, /* 3035 */
128'h00000000000000000000000000000000, /* 3036 */
128'h00000000000000000000000000000000, /* 3037 */
128'h00000000000000000000000000000000, /* 3038 */
128'h00000000000000000000000000000000, /* 3039 */
128'h00000000000000000000000000000000, /* 3040 */
128'h00000000000000000000000000000000, /* 3041 */
128'h00000000000000000000000000000000, /* 3042 */
128'h00000000000000000000000000000000, /* 3043 */
128'h00000000000000000000000000000000, /* 3044 */
128'h00000000000000000000000000000000, /* 3045 */
128'h00000000000000000000000000000000, /* 3046 */
128'h00000000000000000000000000000000, /* 3047 */
128'h00000000000000000000000000000000, /* 3048 */
128'h00000000000000000000000000000000, /* 3049 */
128'h00000000000000000000000000000000, /* 3050 */
128'h00000000000000000000000000000000, /* 3051 */
128'h00000000000000000000000000000000, /* 3052 */
128'h00000000000000000000000000000000, /* 3053 */
128'h00000000000000000000000000000000, /* 3054 */
128'h00000000000000000000000000000000, /* 3055 */
128'h00000000000000000000000000000000, /* 3056 */
128'h00000000000000000000000000000000, /* 3057 */
128'h00000000000000000000000000000000, /* 3058 */
128'h00000000000000000000000000000000, /* 3059 */
128'h00000000000000000000000000000000, /* 3060 */
128'h00000000000000000000000000000000, /* 3061 */
128'h00000000000000000000000000000000, /* 3062 */
128'h00000000000000000000000000000000, /* 3063 */
128'h00000000000000000000000000000000, /* 3064 */
128'h00000000000000000000000000000000, /* 3065 */
128'h00000000000000000000000000000000, /* 3066 */
128'h00000000000000000000000000000000, /* 3067 */
128'h00000000000000000000000000000000, /* 3068 */
128'h00000000000000000000000000000000, /* 3069 */
128'h00000000000000000000000000000000, /* 3070 */
128'h00000000000000000000000000000000, /* 3071 */
128'h00000000000000000000000000000000, /* 3072 */
128'h00000000000000000000000000000000, /* 3073 */
128'h00000000000000000000000000000000, /* 3074 */
128'h00000000000000000000000000000000, /* 3075 */
128'h00000000000000000000000000000000, /* 3076 */
128'h00000000000000000000000000000000, /* 3077 */
128'h00000000000000000000000000000000, /* 3078 */
128'h00000000000000000000000000000000, /* 3079 */
128'h00000000000000000000000000000000, /* 3080 */
128'h00000000000000000000000000000000, /* 3081 */
128'h00000000000000000000000000000000, /* 3082 */
128'h00000000000000000000000000000000, /* 3083 */
128'h00000000000000000000000000000000, /* 3084 */
128'h00000000000000000000000000000000, /* 3085 */
128'h00000000000000000000000000000000, /* 3086 */
128'h00000000000000000000000000000000, /* 3087 */
128'h00000000000000000000000000000000, /* 3088 */
128'h00000000000000000000000000000000, /* 3089 */
128'h00000000000000000000000000000000, /* 3090 */
128'h00000000000000000000000000000000, /* 3091 */
128'h00000000000000000000000000000000, /* 3092 */
128'h00000000000000000000000000000000, /* 3093 */
128'h00000000000000000000000000000000, /* 3094 */
128'h00000000000000000000000000000000, /* 3095 */
128'h00000000000000000000000000000000, /* 3096 */
128'h00000000000000000000000000000000, /* 3097 */
128'h00000000000000000000000000000000, /* 3098 */
128'h00000000000000000000000000000000, /* 3099 */
128'h00000000000000000000000000000000, /* 3100 */
128'h00000000000000000000000000000000, /* 3101 */
128'h00000000000000000000000000000000, /* 3102 */
128'h00000000000000000000000000000000, /* 3103 */
128'h00000000000000000000000000000000, /* 3104 */
128'h00000000000000000000000000000000, /* 3105 */
128'h00000000000000000000000000000000, /* 3106 */
128'h00000000000000000000000000000000, /* 3107 */
128'h00000000000000000000000000000000, /* 3108 */
128'h00000000000000000000000000000000, /* 3109 */
128'h00000000000000000000000000000000, /* 3110 */
128'h00000000000000000000000000000000, /* 3111 */
128'h00000000000000000000000000000000, /* 3112 */
128'h00000000000000000000000000000000, /* 3113 */
128'h00000000000000000000000000000000, /* 3114 */
128'h00000000000000000000000000000000, /* 3115 */
128'h00000000000000000000000000000000, /* 3116 */
128'h00000000000000000000000000000000, /* 3117 */
128'h00000000000000000000000000000000, /* 3118 */
128'h00000000000000000000000000000000, /* 3119 */
128'h00000000000000000000000000000000, /* 3120 */
128'h00000000000000000000000000000000, /* 3121 */
128'h00000000000000000000000000000000, /* 3122 */
128'h00000000000000000000000000000000, /* 3123 */
128'h00000000000000000000000000000000, /* 3124 */
128'h00000000000000000000000000000000, /* 3125 */
128'h00000000000000000000000000000000, /* 3126 */
128'h00000000000000000000000000000000, /* 3127 */
128'h00000000000000000000000000000000, /* 3128 */
128'h00000000000000000000000000000000, /* 3129 */
128'h00000000000000000000000000000000, /* 3130 */
128'h00000000000000000000000000000000, /* 3131 */
128'h00000000000000000000000000000000, /* 3132 */
128'h00000000000000000000000000000000, /* 3133 */
128'h00000000000000000000000000000000, /* 3134 */
128'h00000000000000000000000000000000, /* 3135 */
128'h00000000000000000000000000000000, /* 3136 */
128'h00000000000000000000000000000000, /* 3137 */
128'h00000000000000000000000000000000, /* 3138 */
128'h00000000000000000000000000000000, /* 3139 */
128'h00000000000000000000000000000000, /* 3140 */
128'h00000000000000000000000000000000, /* 3141 */
128'h00000000000000000000000000000000, /* 3142 */
128'h00000000000000000000000000000000, /* 3143 */
128'h00000000000000000000000000000000, /* 3144 */
128'h00000000000000000000000000000000, /* 3145 */
128'h00000000000000000000000000000000, /* 3146 */
128'h00000000000000000000000000000000, /* 3147 */
128'h00000000000000000000000000000000, /* 3148 */
128'h00000000000000000000000000000000, /* 3149 */
128'h00000000000000000000000000000000, /* 3150 */
128'h00000000000000000000000000000000, /* 3151 */
128'h00000000000000000000000000000000, /* 3152 */
128'h00000000000000000000000000000000, /* 3153 */
128'h00000000000000000000000000000000, /* 3154 */
128'h00000000000000000000000000000000, /* 3155 */
128'h00000000000000000000000000000000, /* 3156 */
128'h00000000000000000000000000000000, /* 3157 */
128'h00000000000000000000000000000000, /* 3158 */
128'h00000000000000000000000000000000, /* 3159 */
128'h00000000000000000000000000000000, /* 3160 */
128'h00000000000000000000000000000000, /* 3161 */
128'h00000000000000000000000000000000, /* 3162 */
128'h00000000000000000000000000000000, /* 3163 */
128'h00000000000000000000000000000000, /* 3164 */
128'h00000000000000000000000000000000, /* 3165 */
128'h00000000000000000000000000000000, /* 3166 */
128'h00000000000000000000000000000000, /* 3167 */
128'h00000000000000000000000000000000, /* 3168 */
128'h00000000000000000000000000000000, /* 3169 */
128'h00000000000000000000000000000000, /* 3170 */
128'h00000000000000000000000000000000, /* 3171 */
128'h00000000000000000000000000000000, /* 3172 */
128'h00000000000000000000000000000000, /* 3173 */
128'h00000000000000000000000000000000, /* 3174 */
128'h00000000000000000000000000000000, /* 3175 */
128'h00000000000000000000000000000000, /* 3176 */
128'h00000000000000000000000000000000, /* 3177 */
128'h00000000000000000000000000000000, /* 3178 */
128'h00000000000000000000000000000000, /* 3179 */
128'h00000000000000000000000000000000, /* 3180 */
128'h00000000000000000000000000000000, /* 3181 */
128'h00000000000000000000000000000000, /* 3182 */
128'h00000000000000000000000000000000, /* 3183 */
128'h00000000000000000000000000000000, /* 3184 */
128'h00000000000000000000000000000000, /* 3185 */
128'h00000000000000000000000000000000, /* 3186 */
128'h00000000000000000000000000000000, /* 3187 */
128'h00000000000000000000000000000000, /* 3188 */
128'h00000000000000000000000000000000, /* 3189 */
128'h00000000000000000000000000000000, /* 3190 */
128'h00000000000000000000000000000000, /* 3191 */
128'h00000000000000000000000000000000, /* 3192 */
128'h00000000000000000000000000000000, /* 3193 */
128'h00000000000000000000000000000000, /* 3194 */
128'h00000000000000000000000000000000, /* 3195 */
128'h00000000000000000000000000000000, /* 3196 */
128'h00000000000000000000000000000000, /* 3197 */
128'h00000000000000000000000000000000, /* 3198 */
128'h00000000000000000000000000000000, /* 3199 */
128'h00000000000000000000000000000000, /* 3200 */
128'h00000000000000000000000000000000, /* 3201 */
128'h00000000000000000000000000000000, /* 3202 */
128'h00000000000000000000000000000000, /* 3203 */
128'h00000000000000000000000000000000, /* 3204 */
128'h00000000000000000000000000000000, /* 3205 */
128'h00000000000000000000000000000000, /* 3206 */
128'h00000000000000000000000000000000, /* 3207 */
128'h00000000000000000000000000000000, /* 3208 */
128'h00000000000000000000000000000000, /* 3209 */
128'h00000000000000000000000000000000, /* 3210 */
128'h00000000000000000000000000000000, /* 3211 */
128'h00000000000000000000000000000000, /* 3212 */
128'h00000000000000000000000000000000, /* 3213 */
128'h00000000000000000000000000000000, /* 3214 */
128'h00000000000000000000000000000000, /* 3215 */
128'h00000000000000000000000000000000, /* 3216 */
128'h00000000000000000000000000000000, /* 3217 */
128'h00000000000000000000000000000000, /* 3218 */
128'h00000000000000000000000000000000, /* 3219 */
128'h00000000000000000000000000000000, /* 3220 */
128'h00000000000000000000000000000000, /* 3221 */
128'h00000000000000000000000000000000, /* 3222 */
128'h00000000000000000000000000000000, /* 3223 */
128'h00000000000000000000000000000000, /* 3224 */
128'h00000000000000000000000000000000, /* 3225 */
128'h00000000000000000000000000000000, /* 3226 */
128'h00000000000000000000000000000000, /* 3227 */
128'h00000000000000000000000000000000, /* 3228 */
128'h00000000000000000000000000000000, /* 3229 */
128'h00000000000000000000000000000000, /* 3230 */
128'h00000000000000000000000000000000, /* 3231 */
128'h00000000000000000000000000000000, /* 3232 */
128'h00000000000000000000000000000000, /* 3233 */
128'h00000000000000000000000000000000, /* 3234 */
128'h00000000000000000000000000000000, /* 3235 */
128'h00000000000000000000000000000000, /* 3236 */
128'h00000000000000000000000000000000, /* 3237 */
128'h00000000000000000000000000000000, /* 3238 */
128'h00000000000000000000000000000000, /* 3239 */
128'h00000000000000000000000000000000, /* 3240 */
128'h00000000000000000000000000000000, /* 3241 */
128'h00000000000000000000000000000000, /* 3242 */
128'h00000000000000000000000000000000, /* 3243 */
128'h00000000000000000000000000000000, /* 3244 */
128'h00000000000000000000000000000000, /* 3245 */
128'h00000000000000000000000000000000, /* 3246 */
128'h00000000000000000000000000000000, /* 3247 */
128'h00000000000000000000000000000000, /* 3248 */
128'h00000000000000000000000000000000, /* 3249 */
128'h00000000000000000000000000000000, /* 3250 */
128'h00000000000000000000000000000000, /* 3251 */
128'h00000000000000000000000000000000, /* 3252 */
128'h00000000000000000000000000000000, /* 3253 */
128'h00000000000000000000000000000000, /* 3254 */
128'h00000000000000000000000000000000, /* 3255 */
128'h00000000000000000000000000000000, /* 3256 */
128'h00000000000000000000000000000000, /* 3257 */
128'h00000000000000000000000000000000, /* 3258 */
128'h00000000000000000000000000000000, /* 3259 */
128'h00000000000000000000000000000000, /* 3260 */
128'h00000000000000000000000000000000, /* 3261 */
128'h00000000000000000000000000000000, /* 3262 */
128'h00000000000000000000000000000000, /* 3263 */
128'h00000000000000000000000000000000, /* 3264 */
128'h00000000000000000000000000000000, /* 3265 */
128'h00000000000000000000000000000000, /* 3266 */
128'h00000000000000000000000000000000, /* 3267 */
128'h00000000000000000000000000000000, /* 3268 */
128'h00000000000000000000000000000000, /* 3269 */
128'h00000000000000000000000000000000, /* 3270 */
128'h00000000000000000000000000000000, /* 3271 */
128'h00000000000000000000000000000000, /* 3272 */
128'h00000000000000000000000000000000, /* 3273 */
128'h00000000000000000000000000000000, /* 3274 */
128'h00000000000000000000000000000000, /* 3275 */
128'h00000000000000000000000000000000, /* 3276 */
128'h00000000000000000000000000000000, /* 3277 */
128'h00000000000000000000000000000000, /* 3278 */
128'h00000000000000000000000000000000, /* 3279 */
128'h00000000000000000000000000000000, /* 3280 */
128'h00000000000000000000000000000000, /* 3281 */
128'h00000000000000000000000000000000, /* 3282 */
128'h00000000000000000000000000000000, /* 3283 */
128'h00000000000000000000000000000000, /* 3284 */
128'h00000000000000000000000000000000, /* 3285 */
128'h00000000000000000000000000000000, /* 3286 */
128'h00000000000000000000000000000000, /* 3287 */
128'h00000000000000000000000000000000, /* 3288 */
128'h00000000000000000000000000000000, /* 3289 */
128'h00000000000000000000000000000000, /* 3290 */
128'h00000000000000000000000000000000, /* 3291 */
128'h00000000000000000000000000000000, /* 3292 */
128'h00000000000000000000000000000000, /* 3293 */
128'h00000000000000000000000000000000, /* 3294 */
128'h00000000000000000000000000000000, /* 3295 */
128'h00000000000000000000000000000000, /* 3296 */
128'h00000000000000000000000000000000, /* 3297 */
128'h00000000000000000000000000000000, /* 3298 */
128'h00000000000000000000000000000000, /* 3299 */
128'h00000000000000000000000000000000, /* 3300 */
128'h00000000000000000000000000000000, /* 3301 */
128'h00000000000000000000000000000000, /* 3302 */
128'h00000000000000000000000000000000, /* 3303 */
128'h00000000000000000000000000000000, /* 3304 */
128'h00000000000000000000000000000000, /* 3305 */
128'h00000000000000000000000000000000, /* 3306 */
128'h00000000000000000000000000000000, /* 3307 */
128'h00000000000000000000000000000000, /* 3308 */
128'h00000000000000000000000000000000, /* 3309 */
128'h00000000000000000000000000000000, /* 3310 */
128'h00000000000000000000000000000000, /* 3311 */
128'h00000000000000000000000000000000, /* 3312 */
128'h00000000000000000000000000000000, /* 3313 */
128'h00000000000000000000000000000000, /* 3314 */
128'h00000000000000000000000000000000, /* 3315 */
128'h00000000000000000000000000000000, /* 3316 */
128'h00000000000000000000000000000000, /* 3317 */
128'h00000000000000000000000000000000, /* 3318 */
128'h00000000000000000000000000000000, /* 3319 */
128'h00000000000000000000000000000000, /* 3320 */
128'h00000000000000000000000000000000, /* 3321 */
128'h00000000000000000000000000000000, /* 3322 */
128'h00000000000000000000000000000000, /* 3323 */
128'h00000000000000000000000000000000, /* 3324 */
128'h00000000000000000000000000000000, /* 3325 */
128'h00000000000000000000000000000000, /* 3326 */
128'h00000000000000000000000000000000, /* 3327 */
128'h00000000000000000000000000000000, /* 3328 */
128'h00000000000000000000000000000000, /* 3329 */
128'h00000000000000000000000000000000, /* 3330 */
128'h00000000000000000000000000000000, /* 3331 */
128'h00000000000000000000000000000000, /* 3332 */
128'h00000000000000000000000000000000, /* 3333 */
128'h00000000000000000000000000000000, /* 3334 */
128'h00000000000000000000000000000000, /* 3335 */
128'h00000000000000000000000000000000, /* 3336 */
128'h00000000000000000000000000000000, /* 3337 */
128'h00000000000000000000000000000000, /* 3338 */
128'h00000000000000000000000000000000, /* 3339 */
128'h00000000000000000000000000000000, /* 3340 */
128'h00000000000000000000000000000000, /* 3341 */
128'h00000000000000000000000000000000, /* 3342 */
128'h00000000000000000000000000000000, /* 3343 */
128'h00000000000000000000000000000000, /* 3344 */
128'h00000000000000000000000000000000, /* 3345 */
128'h00000000000000000000000000000000, /* 3346 */
128'h00000000000000000000000000000000, /* 3347 */
128'h00000000000000000000000000000000, /* 3348 */
128'h00000000000000000000000000000000, /* 3349 */
128'h00000000000000000000000000000000, /* 3350 */
128'h00000000000000000000000000000000, /* 3351 */
128'h00000000000000000000000000000000, /* 3352 */
128'h00000000000000000000000000000000, /* 3353 */
128'h00000000000000000000000000000000, /* 3354 */
128'h00000000000000000000000000000000, /* 3355 */
128'h00000000000000000000000000000000, /* 3356 */
128'h00000000000000000000000000000000, /* 3357 */
128'h00000000000000000000000000000000, /* 3358 */
128'h00000000000000000000000000000000, /* 3359 */
128'h00000000000000000000000000000000, /* 3360 */
128'h00000000000000000000000000000000, /* 3361 */
128'h00000000000000000000000000000000, /* 3362 */
128'h00000000000000000000000000000000, /* 3363 */
128'h00000000000000000000000000000000, /* 3364 */
128'h00000000000000000000000000000000, /* 3365 */
128'h00000000000000000000000000000000, /* 3366 */
128'h00000000000000000000000000000000, /* 3367 */
128'h00000000000000000000000000000000, /* 3368 */
128'h00000000000000000000000000000000, /* 3369 */
128'h00000000000000000000000000000000, /* 3370 */
128'h00000000000000000000000000000000, /* 3371 */
128'h00000000000000000000000000000000, /* 3372 */
128'h00000000000000000000000000000000, /* 3373 */
128'h00000000000000000000000000000000, /* 3374 */
128'h00000000000000000000000000000000, /* 3375 */
128'h00000000000000000000000000000000, /* 3376 */
128'h00000000000000000000000000000000, /* 3377 */
128'h00000000000000000000000000000000, /* 3378 */
128'h00000000000000000000000000000000, /* 3379 */
128'h00000000000000000000000000000000, /* 3380 */
128'h00000000000000000000000000000000, /* 3381 */
128'h00000000000000000000000000000000, /* 3382 */
128'h00000000000000000000000000000000, /* 3383 */
128'h00000000000000000000000000000000, /* 3384 */
128'h00000000000000000000000000000000, /* 3385 */
128'h00000000000000000000000000000000, /* 3386 */
128'h00000000000000000000000000000000, /* 3387 */
128'h00000000000000000000000000000000, /* 3388 */
128'h00000000000000000000000000000000, /* 3389 */
128'h00000000000000000000000000000000, /* 3390 */
128'h00000000000000000000000000000000, /* 3391 */
128'h00000000000000000000000000000000, /* 3392 */
128'h00000000000000000000000000000000, /* 3393 */
128'h00000000000000000000000000000000, /* 3394 */
128'h00000000000000000000000000000000, /* 3395 */
128'h00000000000000000000000000000000, /* 3396 */
128'h00000000000000000000000000000000, /* 3397 */
128'h00000000000000000000000000000000, /* 3398 */
128'h00000000000000000000000000000000, /* 3399 */
128'h00000000000000000000000000000000, /* 3400 */
128'h00000000000000000000000000000000, /* 3401 */
128'h00000000000000000000000000000000, /* 3402 */
128'h00000000000000000000000000000000, /* 3403 */
128'h00000000000000000000000000000000, /* 3404 */
128'h00000000000000000000000000000000, /* 3405 */
128'h00000000000000000000000000000000, /* 3406 */
128'h00000000000000000000000000000000, /* 3407 */
128'h00000000000000000000000000000000, /* 3408 */
128'h00000000000000000000000000000000, /* 3409 */
128'h00000000000000000000000000000000, /* 3410 */
128'h00000000000000000000000000000000, /* 3411 */
128'h00000000000000000000000000000000, /* 3412 */
128'h00000000000000000000000000000000, /* 3413 */
128'h00000000000000000000000000000000, /* 3414 */
128'h00000000000000000000000000000000, /* 3415 */
128'h00000000000000000000000000000000, /* 3416 */
128'h00000000000000000000000000000000, /* 3417 */
128'h00000000000000000000000000000000, /* 3418 */
128'h00000000000000000000000000000000, /* 3419 */
128'h00000000000000000000000000000000, /* 3420 */
128'h00000000000000000000000000000000, /* 3421 */
128'h00000000000000000000000000000000, /* 3422 */
128'h00000000000000000000000000000000, /* 3423 */
128'h00000000000000000000000000000000, /* 3424 */
128'h00000000000000000000000000000000, /* 3425 */
128'h00000000000000000000000000000000, /* 3426 */
128'h00000000000000000000000000000000, /* 3427 */
128'h00000000000000000000000000000000, /* 3428 */
128'h00000000000000000000000000000000, /* 3429 */
128'h00000000000000000000000000000000, /* 3430 */
128'h00000000000000000000000000000000, /* 3431 */
128'h00000000000000000000000000000000, /* 3432 */
128'h00000000000000000000000000000000, /* 3433 */
128'h00000000000000000000000000000000, /* 3434 */
128'h00000000000000000000000000000000, /* 3435 */
128'h00000000000000000000000000000000, /* 3436 */
128'h00000000000000000000000000000000, /* 3437 */
128'h00000000000000000000000000000000, /* 3438 */
128'h00000000000000000000000000000000, /* 3439 */
128'h00000000000000000000000000000000, /* 3440 */
128'h00000000000000000000000000000000, /* 3441 */
128'h00000000000000000000000000000000, /* 3442 */
128'h00000000000000000000000000000000, /* 3443 */
128'h00000000000000000000000000000000, /* 3444 */
128'h00000000000000000000000000000000, /* 3445 */
128'h00000000000000000000000000000000, /* 3446 */
128'h00000000000000000000000000000000, /* 3447 */
128'h00000000000000000000000000000000, /* 3448 */
128'h00000000000000000000000000000000, /* 3449 */
128'h00000000000000000000000000000000, /* 3450 */
128'h00000000000000000000000000000000, /* 3451 */
128'h00000000000000000000000000000000, /* 3452 */
128'h00000000000000000000000000000000, /* 3453 */
128'h00000000000000000000000000000000, /* 3454 */
128'h00000000000000000000000000000000, /* 3455 */
128'h00000000000000000000000000000000, /* 3456 */
128'h00000000000000000000000000000000, /* 3457 */
128'h00000000000000000000000000000000, /* 3458 */
128'h00000000000000000000000000000000, /* 3459 */
128'h00000000000000000000000000000000, /* 3460 */
128'h00000000000000000000000000000000, /* 3461 */
128'h00000000000000000000000000000000, /* 3462 */
128'h00000000000000000000000000000000, /* 3463 */
128'h00000000000000000000000000000000, /* 3464 */
128'h00000000000000000000000000000000, /* 3465 */
128'h00000000000000000000000000000000, /* 3466 */
128'h00000000000000000000000000000000, /* 3467 */
128'h00000000000000000000000000000000, /* 3468 */
128'h00000000000000000000000000000000, /* 3469 */
128'h00000000000000000000000000000000, /* 3470 */
128'h00000000000000000000000000000000, /* 3471 */
128'h00000000000000000000000000000000, /* 3472 */
128'h00000000000000000000000000000000, /* 3473 */
128'h00000000000000000000000000000000, /* 3474 */
128'h00000000000000000000000000000000, /* 3475 */
128'h00000000000000000000000000000000, /* 3476 */
128'h00000000000000000000000000000000, /* 3477 */
128'h00000000000000000000000000000000, /* 3478 */
128'h00000000000000000000000000000000, /* 3479 */
128'h00000000000000000000000000000000, /* 3480 */
128'h00000000000000000000000000000000, /* 3481 */
128'h00000000000000000000000000000000, /* 3482 */
128'h00000000000000000000000000000000, /* 3483 */
128'h00000000000000000000000000000000, /* 3484 */
128'h00000000000000000000000000000000, /* 3485 */
128'h00000000000000000000000000000000, /* 3486 */
128'h00000000000000000000000000000000, /* 3487 */
128'h00000000000000000000000000000000, /* 3488 */
128'h00000000000000000000000000000000, /* 3489 */
128'h00000000000000000000000000000000, /* 3490 */
128'h00000000000000000000000000000000, /* 3491 */
128'h00000000000000000000000000000000, /* 3492 */
128'h00000000000000000000000000000000, /* 3493 */
128'h00000000000000000000000000000000, /* 3494 */
128'h00000000000000000000000000000000, /* 3495 */
128'h00000000000000000000000000000000, /* 3496 */
128'h00000000000000000000000000000000, /* 3497 */
128'h00000000000000000000000000000000, /* 3498 */
128'h00000000000000000000000000000000, /* 3499 */
128'h00000000000000000000000000000000, /* 3500 */
128'h00000000000000000000000000000000, /* 3501 */
128'h00000000000000000000000000000000, /* 3502 */
128'h00000000000000000000000000000000, /* 3503 */
128'h00000000000000000000000000000000, /* 3504 */
128'h00000000000000000000000000000000, /* 3505 */
128'h00000000000000000000000000000000, /* 3506 */
128'h00000000000000000000000000000000, /* 3507 */
128'h00000000000000000000000000000000, /* 3508 */
128'h00000000000000000000000000000000, /* 3509 */
128'h00000000000000000000000000000000, /* 3510 */
128'h00000000000000000000000000000000, /* 3511 */
128'h00000000000000000000000000000000, /* 3512 */
128'h00000000000000000000000000000000, /* 3513 */
128'h00000000000000000000000000000000, /* 3514 */
128'h00000000000000000000000000000000, /* 3515 */
128'h00000000000000000000000000000000, /* 3516 */
128'h00000000000000000000000000000000, /* 3517 */
128'h00000000000000000000000000000000, /* 3518 */
128'h00000000000000000000000000000000, /* 3519 */
128'h00000000000000000000000000000000, /* 3520 */
128'h00000000000000000000000000000000, /* 3521 */
128'h00000000000000000000000000000000, /* 3522 */
128'h00000000000000000000000000000000, /* 3523 */
128'h00000000000000000000000000000000, /* 3524 */
128'h00000000000000000000000000000000, /* 3525 */
128'h00000000000000000000000000000000, /* 3526 */
128'h00000000000000000000000000000000, /* 3527 */
128'h00000000000000000000000000000000, /* 3528 */
128'h00000000000000000000000000000000, /* 3529 */
128'h00000000000000000000000000000000, /* 3530 */
128'h00000000000000000000000000000000, /* 3531 */
128'h00000000000000000000000000000000, /* 3532 */
128'h00000000000000000000000000000000, /* 3533 */
128'h00000000000000000000000000000000, /* 3534 */
128'h00000000000000000000000000000000, /* 3535 */
128'h00000000000000000000000000000000, /* 3536 */
128'h00000000000000000000000000000000, /* 3537 */
128'h00000000000000000000000000000000, /* 3538 */
128'h00000000000000000000000000000000, /* 3539 */
128'h00000000000000000000000000000000, /* 3540 */
128'h00000000000000000000000000000000, /* 3541 */
128'h00000000000000000000000000000000, /* 3542 */
128'h00000000000000000000000000000000, /* 3543 */
128'h00000000000000000000000000000000, /* 3544 */
128'h00000000000000000000000000000000, /* 3545 */
128'h00000000000000000000000000000000, /* 3546 */
128'h00000000000000000000000000000000, /* 3547 */
128'h00000000000000000000000000000000, /* 3548 */
128'h00000000000000000000000000000000, /* 3549 */
128'h00000000000000000000000000000000, /* 3550 */
128'h00000000000000000000000000000000, /* 3551 */
128'h00000000000000000000000000000000, /* 3552 */
128'h00000000000000000000000000000000, /* 3553 */
128'h00000000000000000000000000000000, /* 3554 */
128'h00000000000000000000000000000000, /* 3555 */
128'h00000000000000000000000000000000, /* 3556 */
128'h00000000000000000000000000000000, /* 3557 */
128'h00000000000000000000000000000000, /* 3558 */
128'h00000000000000000000000000000000, /* 3559 */
128'h00000000000000000000000000000000, /* 3560 */
128'h00000000000000000000000000000000, /* 3561 */
128'h00000000000000000000000000000000, /* 3562 */
128'h00000000000000000000000000000000, /* 3563 */
128'h00000000000000000000000000000000, /* 3564 */
128'h00000000000000000000000000000000, /* 3565 */
128'h00000000000000000000000000000000, /* 3566 */
128'h00000000000000000000000000000000, /* 3567 */
128'h00000000000000000000000000000000, /* 3568 */
128'h00000000000000000000000000000000, /* 3569 */
128'h00000000000000000000000000000000, /* 3570 */
128'h00000000000000000000000000000000, /* 3571 */
128'h00000000000000000000000000000000, /* 3572 */
128'h00000000000000000000000000000000, /* 3573 */
128'h00000000000000000000000000000000, /* 3574 */
128'h00000000000000000000000000000000, /* 3575 */
128'h00000000000000000000000000000000, /* 3576 */
128'h00000000000000000000000000000000, /* 3577 */
128'h00000000000000000000000000000000, /* 3578 */
128'h00000000000000000000000000000000, /* 3579 */
128'h00000000000000000000000000000000, /* 3580 */
128'h00000000000000000000000000000000, /* 3581 */
128'h00000000000000000000000000000000, /* 3582 */
128'h00000000000000000000000000000000, /* 3583 */
128'h00000000000000000000000000000000, /* 3584 */
128'h00000000000000000000000000000000, /* 3585 */
128'h00000000000000000000000000000000, /* 3586 */
128'h00000000000000000000000000000000, /* 3587 */
128'h00000000000000000000000000000000, /* 3588 */
128'h00000000000000000000000000000000, /* 3589 */
128'h00000000000000000000000000000000, /* 3590 */
128'h00000000000000000000000000000000, /* 3591 */
128'h00000000000000000000000000000000, /* 3592 */
128'h00000000000000000000000000000000, /* 3593 */
128'h00000000000000000000000000000000, /* 3594 */
128'h00000000000000000000000000000000, /* 3595 */
128'h00000000000000000000000000000000, /* 3596 */
128'h00000000000000000000000000000000, /* 3597 */
128'h00000000000000000000000000000000, /* 3598 */
128'h00000000000000000000000000000000, /* 3599 */
128'h00000000000000000000000000000000, /* 3600 */
128'h00000000000000000000000000000000, /* 3601 */
128'h00000000000000000000000000000000, /* 3602 */
128'h00000000000000000000000000000000, /* 3603 */
128'h00000000000000000000000000000000, /* 3604 */
128'h00000000000000000000000000000000, /* 3605 */
128'h00000000000000000000000000000000, /* 3606 */
128'h00000000000000000000000000000000, /* 3607 */
128'h00000000000000000000000000000000, /* 3608 */
128'h00000000000000000000000000000000, /* 3609 */
128'h00000000000000000000000000000000, /* 3610 */
128'h00000000000000000000000000000000, /* 3611 */
128'h00000000000000000000000000000000, /* 3612 */
128'h00000000000000000000000000000000, /* 3613 */
128'h00000000000000000000000000000000, /* 3614 */
128'h00000000000000000000000000000000, /* 3615 */
128'h00000000000000000000000000000000, /* 3616 */
128'h00000000000000000000000000000000, /* 3617 */
128'h00000000000000000000000000000000, /* 3618 */
128'h00000000000000000000000000000000, /* 3619 */
128'h00000000000000000000000000000000, /* 3620 */
128'h00000000000000000000000000000000, /* 3621 */
128'h00000000000000000000000000000000, /* 3622 */
128'h00000000000000000000000000000000, /* 3623 */
128'h00000000000000000000000000000000, /* 3624 */
128'h00000000000000000000000000000000, /* 3625 */
128'h00000000000000000000000000000000, /* 3626 */
128'h00000000000000000000000000000000, /* 3627 */
128'h00000000000000000000000000000000, /* 3628 */
128'h00000000000000000000000000000000, /* 3629 */
128'h00000000000000000000000000000000, /* 3630 */
128'h00000000000000000000000000000000, /* 3631 */
128'h00000000000000000000000000000000, /* 3632 */
128'h00000000000000000000000000000000, /* 3633 */
128'h00000000000000000000000000000000, /* 3634 */
128'h00000000000000000000000000000000, /* 3635 */
128'h00000000000000000000000000000000, /* 3636 */
128'h00000000000000000000000000000000, /* 3637 */
128'h00000000000000000000000000000000, /* 3638 */
128'h00000000000000000000000000000000, /* 3639 */
128'h00000000000000000000000000000000, /* 3640 */
128'h00000000000000000000000000000000, /* 3641 */
128'h00000000000000000000000000000000, /* 3642 */
128'h00000000000000000000000000000000, /* 3643 */
128'h00000000000000000000000000000000, /* 3644 */
128'h00000000000000000000000000000000, /* 3645 */
128'h00000000000000000000000000000000, /* 3646 */
128'h00000000000000000000000000000000, /* 3647 */
128'h00000000000000000000000000000000, /* 3648 */
128'h00000000000000000000000000000000, /* 3649 */
128'h00000000000000000000000000000000, /* 3650 */
128'h00000000000000000000000000000000, /* 3651 */
128'h00000000000000000000000000000000, /* 3652 */
128'h00000000000000000000000000000000, /* 3653 */
128'h00000000000000000000000000000000, /* 3654 */
128'h00000000000000000000000000000000, /* 3655 */
128'h00000000000000000000000000000000, /* 3656 */
128'h00000000000000000000000000000000, /* 3657 */
128'h00000000000000000000000000000000, /* 3658 */
128'h00000000000000000000000000000000, /* 3659 */
128'h00000000000000000000000000000000, /* 3660 */
128'h00000000000000000000000000000000, /* 3661 */
128'h00000000000000000000000000000000, /* 3662 */
128'h00000000000000000000000000000000, /* 3663 */
128'h00000000000000000000000000000000, /* 3664 */
128'h00000000000000000000000000000000, /* 3665 */
128'h00000000000000000000000000000000, /* 3666 */
128'h00000000000000000000000000000000, /* 3667 */
128'h00000000000000000000000000000000, /* 3668 */
128'h00000000000000000000000000000000, /* 3669 */
128'h00000000000000000000000000000000, /* 3670 */
128'h00000000000000000000000000000000, /* 3671 */
128'h00000000000000000000000000000000, /* 3672 */
128'h00000000000000000000000000000000, /* 3673 */
128'h00000000000000000000000000000000, /* 3674 */
128'h00000000000000000000000000000000, /* 3675 */
128'h00000000000000000000000000000000, /* 3676 */
128'h00000000000000000000000000000000, /* 3677 */
128'h00000000000000000000000000000000, /* 3678 */
128'h00000000000000000000000000000000, /* 3679 */
128'h00000000000000000000000000000000, /* 3680 */
128'h00000000000000000000000000000000, /* 3681 */
128'h00000000000000000000000000000000, /* 3682 */
128'h00000000000000000000000000000000, /* 3683 */
128'h00000000000000000000000000000000, /* 3684 */
128'h00000000000000000000000000000000, /* 3685 */
128'h00000000000000000000000000000000, /* 3686 */
128'h00000000000000000000000000000000, /* 3687 */
128'h00000000000000000000000000000000, /* 3688 */
128'h00000000000000000000000000000000, /* 3689 */
128'h00000000000000000000000000000000, /* 3690 */
128'h00000000000000000000000000000000, /* 3691 */
128'h00000000000000000000000000000000, /* 3692 */
128'h00000000000000000000000000000000, /* 3693 */
128'h00000000000000000000000000000000, /* 3694 */
128'h00000000000000000000000000000000, /* 3695 */
128'h00000000000000000000000000000000, /* 3696 */
128'h00000000000000000000000000000000, /* 3697 */
128'h00000000000000000000000000000000, /* 3698 */
128'h00000000000000000000000000000000, /* 3699 */
128'h00000000000000000000000000000000, /* 3700 */
128'h00000000000000000000000000000000, /* 3701 */
128'h00000000000000000000000000000000, /* 3702 */
128'h00000000000000000000000000000000, /* 3703 */
128'h00000000000000000000000000000000, /* 3704 */
128'h00000000000000000000000000000000, /* 3705 */
128'h00000000000000000000000000000000, /* 3706 */
128'h00000000000000000000000000000000, /* 3707 */
128'h00000000000000000000000000000000, /* 3708 */
128'h00000000000000000000000000000000, /* 3709 */
128'h00000000000000000000000000000000, /* 3710 */
128'h00000000000000000000000000000000, /* 3711 */
128'h00000000000000000000000000000000, /* 3712 */
128'h00000000000000000000000000000000, /* 3713 */
128'h00000000000000000000000000000000, /* 3714 */
128'h00000000000000000000000000000000, /* 3715 */
128'h00000000000000000000000000000000, /* 3716 */
128'h00000000000000000000000000000000, /* 3717 */
128'h00000000000000000000000000000000, /* 3718 */
128'h00000000000000000000000000000000, /* 3719 */
128'h00000000000000000000000000000000, /* 3720 */
128'h00000000000000000000000000000000, /* 3721 */
128'h00000000000000000000000000000000, /* 3722 */
128'h00000000000000000000000000000000, /* 3723 */
128'h00000000000000000000000000000000, /* 3724 */
128'h00000000000000000000000000000000, /* 3725 */
128'h00000000000000000000000000000000, /* 3726 */
128'h00000000000000000000000000000000, /* 3727 */
128'h00000000000000000000000000000000, /* 3728 */
128'h00000000000000000000000000000000, /* 3729 */
128'h00000000000000000000000000000000, /* 3730 */
128'h00000000000000000000000000000000, /* 3731 */
128'h00000000000000000000000000000000, /* 3732 */
128'h00000000000000000000000000000000, /* 3733 */
128'h00000000000000000000000000000000, /* 3734 */
128'h00000000000000000000000000000000, /* 3735 */
128'h00000000000000000000000000000000, /* 3736 */
128'h00000000000000000000000000000000, /* 3737 */
128'h00000000000000000000000000000000, /* 3738 */
128'h00000000000000000000000000000000, /* 3739 */
128'h00000000000000000000000000000000, /* 3740 */
128'h00000000000000000000000000000000, /* 3741 */
128'h00000000000000000000000000000000, /* 3742 */
128'h00000000000000000000000000000000, /* 3743 */
128'h00000000000000000000000000000000, /* 3744 */
128'h00000000000000000000000000000000, /* 3745 */
128'h00000000000000000000000000000000, /* 3746 */
128'h00000000000000000000000000000000, /* 3747 */
128'h00000000000000000000000000000000, /* 3748 */
128'h00000000000000000000000000000000, /* 3749 */
128'h00000000000000000000000000000000, /* 3750 */
128'h00000000000000000000000000000000, /* 3751 */
128'h00000000000000000000000000000000, /* 3752 */
128'h00000000000000000000000000000000, /* 3753 */
128'h00000000000000000000000000000000, /* 3754 */
128'h00000000000000000000000000000000, /* 3755 */
128'h00000000000000000000000000000000, /* 3756 */
128'h00000000000000000000000000000000, /* 3757 */
128'h00000000000000000000000000000000, /* 3758 */
128'h00000000000000000000000000000000, /* 3759 */
128'h00000000000000000000000000000000, /* 3760 */
128'h00000000000000000000000000000000, /* 3761 */
128'h00000000000000000000000000000000, /* 3762 */
128'h00000000000000000000000000000000, /* 3763 */
128'h00000000000000000000000000000000, /* 3764 */
128'h00000000000000000000000000000000, /* 3765 */
128'h00000000000000000000000000000000, /* 3766 */
128'h00000000000000000000000000000000, /* 3767 */
128'h00000000000000000000000000000000, /* 3768 */
128'h00000000000000000000000000000000, /* 3769 */
128'h00000000000000000000000000000000, /* 3770 */
128'h00000000000000000000000000000000, /* 3771 */
128'h00000000000000000000000000000000, /* 3772 */
128'h00000000000000000000000000000000, /* 3773 */
128'h00000000000000000000000000000000, /* 3774 */
128'h00000000000000000000000000000000, /* 3775 */
128'h00000000000000000000000000000000, /* 3776 */
128'h00000000000000000000000000000000, /* 3777 */
128'h00000000000000000000000000000000, /* 3778 */
128'h00000000000000000000000000000000, /* 3779 */
128'h00000000000000000000000000000000, /* 3780 */
128'h00000000000000000000000000000000, /* 3781 */
128'h00000000000000000000000000000000, /* 3782 */
128'h00000000000000000000000000000000, /* 3783 */
128'h00000000000000000000000000000000, /* 3784 */
128'h00000000000000000000000000000000, /* 3785 */
128'h00000000000000000000000000000000, /* 3786 */
128'h00000000000000000000000000000000, /* 3787 */
128'h00000000000000000000000000000000, /* 3788 */
128'h00000000000000000000000000000000, /* 3789 */
128'h00000000000000000000000000000000, /* 3790 */
128'h00000000000000000000000000000000, /* 3791 */
128'h00000000000000000000000000000000, /* 3792 */
128'h00000000000000000000000000000000, /* 3793 */
128'h00000000000000000000000000000000, /* 3794 */
128'h00000000000000000000000000000000, /* 3795 */
128'h00000000000000000000000000000000, /* 3796 */
128'h00000000000000000000000000000000, /* 3797 */
128'h00000000000000000000000000000000, /* 3798 */
128'h00000000000000000000000000000000, /* 3799 */
128'h00000000000000000000000000000000, /* 3800 */
128'h00000000000000000000000000000000, /* 3801 */
128'h00000000000000000000000000000000, /* 3802 */
128'h00000000000000000000000000000000, /* 3803 */
128'h00000000000000000000000000000000, /* 3804 */
128'h00000000000000000000000000000000, /* 3805 */
128'h00000000000000000000000000000000, /* 3806 */
128'h00000000000000000000000000000000, /* 3807 */
128'h00000000000000000000000000000000, /* 3808 */
128'h00000000000000000000000000000000, /* 3809 */
128'h00000000000000000000000000000000, /* 3810 */
128'h00000000000000000000000000000000, /* 3811 */
128'h00000000000000000000000000000000, /* 3812 */
128'h00000000000000000000000000000000, /* 3813 */
128'h00000000000000000000000000000000, /* 3814 */
128'h00000000000000000000000000000000, /* 3815 */
128'h00000000000000000000000000000000, /* 3816 */
128'h00000000000000000000000000000000, /* 3817 */
128'h00000000000000000000000000000000, /* 3818 */
128'h00000000000000000000000000000000, /* 3819 */
128'h00000000000000000000000000000000, /* 3820 */
128'h00000000000000000000000000000000, /* 3821 */
128'h00000000000000000000000000000000, /* 3822 */
128'h00000000000000000000000000000000, /* 3823 */
128'h00000000000000000000000000000000, /* 3824 */
128'h00000000000000000000000000000000, /* 3825 */
128'h00000000000000000000000000000000, /* 3826 */
128'h00000000000000000000000000000000, /* 3827 */
128'h00000000000000000000000000000000, /* 3828 */
128'h00000000000000000000000000000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00000000000000000000000000000000, /* 3840 */
128'h00000000000000000000000000000000, /* 3841 */
128'h00000000000000000000000000000000, /* 3842 */
128'h00000000000000000000000000000000, /* 3843 */
128'h00000000000000000000000000000000, /* 3844 */
128'h00000000000000000000000000000000, /* 3845 */
128'h00000000000000000000000000000000, /* 3846 */
128'h00000000000000000000000000000000, /* 3847 */
128'h00000000000000000000000000000000, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule

