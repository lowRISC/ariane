/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'h01111113fff1011b0000613711249463, /*    1 */
128'h00008297000280e70ce2829300008297, /*    2 */
128'h000280e713050513000005170f428293, /*    3 */
128'hbc5606130000c617fc05859300000597, /*    4 */
128'h000f4eb701169693fff6869b000066b7, /*    5 */
128'h0085b703fffe8e930005b703240e8e9b, /*    6 */
128'hff81011301b111130110011bfe0e9ae3, /*    7 */
128'h0085b70300e6b0230005b7030006b703, /*    8 */
128'h0185b70300e6b8230105b70300e6b423, /*    9 */
128'hfcc5cce3020686930205859300e6bc23, /*   10 */
128'h40b787b300d787b30147879300000797, /*   11 */
128'h30579073090787930000079700078067, /*   12 */
128'h3c8606130000c617c30585930000c597, /*   13 */
128'h0005bc230005b8230005b4230005b023, /*   14 */
128'h020004b772c090effec5c6e302058593, /*   15 */
128'h02000937004484930124a02300100913, /*   16 */
128'h3440297310500073ff24c6e34009091b, /*   17 */
128'hf1402973020004b7fe090ae300897913, /*   18 */
128'h0004a903000920230099093300291913, /*   19 */
128'h4009091b0200093700448493fe091ee3, /*   20 */
128'h1050007334102373342022f3ff24c6e3, /*   21 */
128'h41206d6f7266206f6c6c6548ffdff06f, /*   22 */
128'h617720657361656c502021656e616972, /*   23 */
128'h000a2e2e2e746e656d6f6d2061207469, /*   24 */
128'h00000000000000000000000000000000, /*   25 */
128'h00000000000000000000000000000000, /*   26 */
128'h00000000000000000000000000000000, /*   27 */
128'h00000000000000000000000000000000, /*   28 */
128'h00000000000000000000000000000000, /*   29 */
128'h00000000000000000000000000000000, /*   30 */
128'h00000000000000000000000000000000, /*   31 */
128'hd963454c0005cc635735c28587ae6914, /*   32 */
128'he21c97b6470102a787b30a00051300b7, /*   33 */
128'h853e85b200030563018533038082853a, /*   34 */
128'h838686930000c697b7edfda007138302, /*   35 */
128'h87930000c79762949d0707130000c717, /*   36 */
128'h87b30280069302d787bb878d8f999c67, /*   37 */
128'h47148082853a470100e7956397ba02d7, /*   38 */
128'hf0efe4061141b7f502870713fea68de3, /*   39 */
128'hbfe545018082014160a26108c509fbbf, /*   40 */
128'hf0efe852ec4ef04af426f822fc067139, /*   41 */
128'h0000ba17440144814985892acd31f9bf, /*   42 */
128'he091450100f44d6300c92783384a0a13, /*   43 */
128'h61216a4269e2790274a2744270e25535, /*   44 */
128'h67a2ed19f29ff0ef854a85a200308082, /*   45 */
128'h50ef8552000995632485cb990087c783, /*   46 */
128'h0513bf65240524c080ef498165224e60, /*   47 */
128'hf2dff0efe42ef406f0227179b7c1fda0, /*   48 */
128'h842aee7ff0ef083065a2c105fda00413, /*   49 */
128'h00f7096300c547030ff007936562e911, /*   50 */
128'h547980826145740270a28522212080ef, /*   51 */
128'hf0efec4ef04af426f822fc067139bfd5, /*   52 */
128'h0000a9970ff00913440184aacd01eebf, /*   53 */
128'h74a2744270e200f4496344dc4a498993, /*   54 */
128'hf0ef852685a200308082612169e27902, /*   55 */
128'h85a20127896300c7c78367a2ed09e83f, /*   56 */
128'hb7d924051ac080ef6522442050ef854e, /*   57 */
128'he8dff0ef892eec26f406e84af0227179, /*   58 */
128'he45ff0ef84aa85ca0030c11dfda00413, /*   59 */
128'h448505130000a517864a608ced01842a, /*   60 */
128'h740270a2852216e080ef6522404050ef, /*   61 */
128'hf406ec26f022717980826145694264e2, /*   62 */
128'h85a6842ac11dfda00413e47ff0ef84ae, /*   63 */
128'hcf63445c3cc050ef420505130000a517, /*   64 */
128'h5435134080ef41e505130000a51700f4, /*   65 */
128'h003085228082614564e2740270a28522, /*   66 */
128'h108080ef6522f565842adcfff0ef85a6, /*   67 */
128'h5479fcf71be30ff0079300c7c70367a2, /*   68 */
128'he50965a2de1ff0eff406e42e7179bfc1, /*   69 */
128'hf96dd97ff0ef08308082614570a24501, /*   70 */
128'he42eec064108842ae8221101bfc56562, /*   71 */
128'h852200030e6302053303c919db9ff0ef, /*   72 */
128'h60e2fda005138302610560e265a26442, /*   73 */
128'h0000b7977139bfdd4501808261056442, /*   74 */
128'h04130000b417f426f822639c5c478793, /*   75 */
128'h043b840d8c0574e484930000b4977564, /*   76 */
128'h892afc06e852ec4ef04a0280079302f4, /*   77 */
128'h942602f4043335ea0a130000aa1789ae, /*   78 */
128'h69e2790274a2744270e2450100849b63, /*   79 */
128'h2c8050ef855285ca6090808261216a42, /*   80 */
128'hbfc902848493c5016f5060ef854a608c, /*   81 */
128'hb7e16522f569cdbff0ef852685ce0030, /*   82 */
128'h84b68432e42efc06f04af426f8227139, /*   83 */
128'hcb5ff0ef083065a2c115cf7ff0ef893a, /*   84 */
128'h70e2978285a2615c862686ca6562e519, /*   85 */
128'hbfc5fda0051380826121790274a27442, /*   86 */
128'h84b68432e42efc06f04af426f8227139, /*   87 */
128'hc75ff0ef083065a2c115cb7ff0ef893a, /*   88 */
128'h70e2978285a2655c862686ca6562e519, /*   89 */
128'hbfc5fda0051380826121790274a27442, /*   90 */
128'hc7dff0ef84b2e42ef822fc06f4267139, /*   91 */
128'h701ce509c39ff0ef842a083065a2c105, /*   92 */
128'h8082612174a2744270e2978285a66562, /*   93 */
128'h2785c3190017f713419cbfcdfda00513, /*   94 */
128'hd71b8e5927a106220086571b419cc19c, /*   95 */
128'h0ff77713c19c0087d7138ed906a20086, /*   96 */
128'h122300d5112300c510238fd90087979b, /*   97 */
128'hf022f4067179419c80820005132300f5, /*   98 */
128'h419c00f510230457879b6785c19c27d1, /*   99 */
128'h0087979b0ff777130087d713c632842a, /*  100 */
128'hc4360509084c57fd460900f11a238fd9, /*  101 */
128'h05130161059346097df060ef00f11b23, /*  102 */
128'h00041323082c462147c17d1060ef0044, /*  103 */
128'h00f404a347c57bd060efec3e00840513, /*  104 */
128'h7a7060ef00c4051300041523006c4611, /*  105 */
128'h0144069379b060ef01040513002c4611, /*  106 */
128'hfed79ce39f31ffe7d6030789470187a2, /*  107 */
128'h9fb94107d71b9fb9934117424107579b, /*  108 */
128'h80826145740270a200f41523fff7c793, /*  109 */
128'h97b64721678563943e8787930000b797, /*  110 */
128'hc7bb27850077e793fff6079b8007bc23, /*  111 */
128'h678500f747630005071b6805450102e7, /*  112 */
128'h00e588b300351713808280c6b82396be, /*  113 */
128'hbfe1050501173023973697420008b883, /*  114 */
128'he406450185aa86220005841be0221141, /*  115 */
128'h717980820141640260a28522fa1ff0ef, /*  116 */
128'he436f4064619051984b2842aec26f022, /*  117 */
128'h6d7060ef85b64619852266a26e3060ef, /*  118 */
128'h00e4859b70a27402852200f4162347a1, /*  119 */
128'h6785737dc5010113fadff06f614564e2, /*  120 */
128'h38913c233a113423392138233a813023, /*  121 */
128'h3761382337513c233941302339313423, /*  122 */
128'h35a1382335913c233781302337713423, /*  123 */
128'hd00007b7943e747d978a911a35078793, /*  124 */
128'hf0040023e0040023ca040b23ce042023, /*  125 */
128'h00e7ea63892a5800073797aad0040023, /*  126 */
128'ha0017db040ef05e505130000a51785aa, /*  127 */
128'h871374fd678524f71d63478900054703, /*  128 */
128'h970a350787139abacd848a93970a3507, /*  129 */
128'h49818a368cb28baed0048c13cb848b13, /*  130 */
128'hcd03013907b395ca0f0985939c3a9b3a, /*  131 */
128'h89bb058902a0071329890f07c7830015, /*  132 */
128'h22e78f63471904f76b6326e78b6301a9, /*  133 */
128'hcc848513470d2ae78963470502f76263, /*  134 */
128'h40ef162505130000a51785be22e78763, /*  135 */
128'hfee794e3473d22e783634731bf4d7570, /*  136 */
128'h953e866ae0048513978a350787936785, /*  137 */
128'h03600713b769e00d00235a1060ef9d22, /*  138 */
128'h20e78e630330071300f76e6322e78163, /*  139 */
128'haac94605cb648513fae798e303500713, /*  140 */
128'hf8e79ce30ff0071324e7856303800713, /*  141 */
128'h8363479924f58363747d479500614583, /*  142 */
128'h16079263000ca7833af59f63478938f5, /*  143 */
128'h0593ce4405134985978a350a87936a85, /*  144 */
128'h8793529060ef013ca023953e46110109, /*  145 */
128'h953e461101490593ce840513978a350a, /*  146 */
128'h54e25a52f3c505130000a517513060ef, /*  147 */
128'hcf840913978a350a8793693040efde02, /*  148 */
128'h03a3478d49d060ef854a55fd4619993e, /*  149 */
128'h978a350a879346f115231350079300f1, /*  150 */
128'h46c1051385a6460594becb740493c2a6, /*  151 */
128'h879346f106a3032007934c1060efc0d2, /*  152 */
128'h051346114a1195becf040593978a350a, /*  153 */
128'h09a30360079349d060ef4741072346f1, /*  154 */
128'h461195becf440593978a350a879346f1, /*  155 */
128'h460557fd47b060ef47410a2347510513, /*  156 */
128'h0d23000103a346f10ca347b1051385a6, /*  157 */
128'h45810f00061310200793461060ef4731, /*  158 */
128'h1d23101007933ff060efde3e37a10513, /*  159 */
128'h36f10e233961051385de4799464136f1, /*  160 */
128'h679946f113232637879377e1433060ef, /*  161 */
128'h0413978a350a879346f1142335378793, /*  162 */
128'h051385a20440061304300693943ecec4, /*  163 */
128'h35e1051385a2460156fdba5ff0ef3721, /*  164 */
128'hcf3ff0ef0e8885de86ca5672bd9ff0ef, /*  165 */
128'h398134833a0134033a813083911a6305, /*  166 */
128'h37813a8338013a033881398339013903, /*  167 */
128'h35813c8336013c0336813b8337013b03, /*  168 */
128'h4611cd04851380823b01011335013d03, /*  169 */
128'h87936785a00d953e978a350787936785, /*  170 */
128'h60ef9d22953e866af0048513978a3507, /*  171 */
128'h377060ef85564611b3bdf00d00233850, /*  172 */
128'h978a350787936785bfdd855a4611b395, /*  173 */
128'hce04578335b060ef4611953ece048513, /*  174 */
128'h578300f411238fd90087979b0087d71b, /*  175 */
128'h00f410238fd90087979b0087d71bce24, /*  176 */
128'h866ab749cc048513bb39cef42023401c, /*  177 */
128'h2783b321d00d002331f060ef9d228562, /*  178 */
128'h0000a51700fa2023478512079a63000a, /*  179 */
128'h0e88010905934611491040efd4c50513, /*  180 */
128'hcb840513978a3504879364852f3060ef, /*  181 */
128'h353147032db060ef014905934611953e, /*  182 */
128'h0000a517350145833511460335214683, /*  183 */
128'h00a1468335015783451040efd1c50513, /*  184 */
128'h352157831cf71e230000b71700914603, /*  185 */
128'h0000b717d1c505130000a51700814583, /*  186 */
128'h01b1470341d040ef00b147031cf71323, /*  187 */
128'h0000a517018145830191460301a14683, /*  188 */
128'h0121468301314703401040efd1c50513, /*  189 */
128'hd20505130000a5170101458301114603, /*  190 */
128'h05130000a51755c2010157833e5040ef, /*  191 */
128'hb7170121578316f713230000b717d2e5, /*  192 */
128'hf6bb02f5d63b03c0079314f71e230000, /*  193 */
128'h02f5d5bbe107879b678502f6763b02f5, /*  194 */
128'h95bee0040593978a350487933a5040ef, /*  195 */
128'h3504879338d040efd08505130000a517, /*  196 */
128'hd00505130000a51795be978af0040593, /*  197 */
128'h40efd0a505130000a517bbf5375040ef, /*  198 */
128'h20234785de0794e3000a2783b3fd3670, /*  199 */
128'ha51734b040efcfe505130000a51700fa, /*  200 */
128'h35078793678533f040efd02505130000, /*  201 */
128'hd08505130000a51795be978ad0040593, /*  202 */
128'hb34d31b040efd0e505130000a517bf45, /*  203 */
128'hf852fc4ee0cae4a6e8a2ec86711d737d, /*  204 */
128'h6a85d22505130000a517911a89aaf456, /*  205 */
128'h0493978a020a8793747d2f3040efca02, /*  206 */
128'hb7970fb060ef852655fd461994beff84, /*  207 */
128'hc83e4a05fef40913439cdb2787930000, /*  208 */
128'h993e978a020a879312f11d2313500793, /*  209 */
128'h0793119060ef014107a31a68460585ca, /*  210 */
128'h020a879312f10f23479112f10ea30370, /*  211 */
128'h60ef13f10513461195beff040593978a, /*  212 */
128'h14f101a314510513460585ca57fd0f50, /*  213 */
128'h0fc007930db060ef000107a315410223, /*  214 */
128'h079060efca3e04a1051345810f000613, /*  215 */
128'h05134641479985ce04f1152310100793, /*  216 */
128'h2637879377e10ad060ef04f106230661, /*  217 */
128'h879312f11c2335378793679912f11b23, /*  218 */
128'h06930421051385a2943e1451978a020a, /*  219 */
128'h02e1051385a2821ff0ef044006130430, /*  220 */
128'h85ce86a610084652855ff0ef460156fd, /*  221 */
128'h64a66446450160e6911a630596fff0ef, /*  222 */
128'ha51785aa808261257aa27a4279e26906, /*  223 */
128'hf0a2f48671591cf0406fc12505130000, /*  224 */
128'h05a1051384aa81010113e4cee8caeca6, /*  225 */
128'h60efd602e83eec3ae442893689b2e046, /*  226 */
128'h6762747d97ba81078793101867850150, /*  227 */
128'h0521051385a2864a86ba943e7fc40413, /*  228 */
128'h863e86c285a267c26822f94ff0efd64e, /*  229 */
128'h85a6180856326882fc4ff0ef03e10513, /*  230 */
128'h7406450170a67f0101138ddff0ef86c6, /*  231 */
128'he222e606716d8082616569a6694664e6, /*  232 */
128'h00254703003547830045480300554883, /*  233 */
128'h85930000a597842a0005460300154683, /*  234 */
128'h852211b040efb76505130000a517b765, /*  235 */
128'h85930000a597860ac10d842ae01ff0ef, /*  236 */
128'h85220fb040efb7e505130000a517b565, /*  237 */
128'hb98505130000a51780826151641260b2, /*  238 */
128'h7159b7cd0dd040efe007a8230000b797, /*  239 */
128'hec66f062f45ef85afc56e0d2e4ceeca6, /*  240 */
128'h44818aae89aae46ee8caf0a2f486e86a, /*  241 */
128'hb70b0b130000ab17870a0a130000ba17, /*  242 */
128'h0000ac97b7cc0c130000ac1706000b93, /*  243 */
128'h035441630004841bfff58d1bb6cc8c93, /*  244 */
128'h7b427ae26a0669a6694664e6740670a6, /*  245 */
128'hc01d808261656da26d426ce27c027ba2, /*  246 */
128'hff04891305d040ef855ae39d00f47793, /*  247 */
128'h6a8505130000a51702879d630009079b, /*  248 */
128'hc583009987b303f040ef8552045040ef, /*  249 */
128'h126302b040efb16505130000a5170007, /*  250 */
128'h87b3a80500f979134d81fffd4913068d, /*  251 */
128'he7630ff7f793fe05879b0007c5830129, /*  252 */
128'h40ef8562b75d0905001040ef856600fb, /*  253 */
128'hff2dcce32d857ee040ef8552bfdd7f60, /*  254 */
128'h079b4124093b7de040ef00f4f913855a, /*  255 */
128'h40ef62a505130000a51700f45a630009, /*  256 */
128'h879b0007c583012987b3bf1504857c60, /*  257 */
128'h7a8040ef856600fbe7630ff7f793fe05, /*  258 */
128'hec267179bfdd79e040ef8562b7f10905, /*  259 */
128'ha697893289ae84b6f022f406e44ee84a, /*  260 */
128'ha68686930000a697c50931a686930000, /*  261 */
128'ha60606130000a617f187071300009717, /*  262 */
128'h5d6300098f63842a720040ef854a85a6, /*  263 */
128'ha48606130000a61786ce40a485bb0095, /*  264 */
128'h00f44463ffe4879b9c29702040ef954a, /*  265 */
128'ha18585930000a59700890533ffd4841b, /*  266 */
128'h69a2694264e2854a740270a22de060ef, /*  267 */
128'h7115f73ff06f4581862e86b280826145, /*  268 */
128'h002cfebff0efed8645050c800613002c, /*  269 */
128'h450160ee6ec040efa00505130000a517, /*  270 */
128'h6963862e9ff787133b9ad7b78082612d, /*  271 */
128'h079304a7676323f78713000f47b704a7, /*  272 */
128'h0000b7173e80079346890ca7fc633e70, /*  273 */
128'hec0600074903e04a973611019a470713, /*  274 */
128'h690264a260e2644202091663e426e822, /*  275 */
128'h6880406f61059a6505130000a51785aa, /*  276 */
128'hbf7d240787934685b7d9a00787934681, /*  277 */
128'h47293e800793c81502f555b302f57433, /*  278 */
128'h0713cf3902f4773346a547a90687e263, /*  279 */
128'h743302f457b30640071300877d630630, /*  280 */
128'h0000a517943e001444130324341302e4, /*  281 */
128'ha51785a2c80162e040ef84b295c50513, /*  282 */
128'h862660e2644261e040ef952505130000, /*  283 */
128'h6105942505130000a517690264a285ca, /*  284 */
128'hf46302f45733bf6102e454336040406f, /*  285 */
128'h0000a51785aabf554401bf51843a0086, /*  286 */
128'h86bb459958d94701862ebfa18fc50513, /*  287 */
128'h1702cf8500f557b3883e03c6879b02e8, /*  288 */
128'he426972e11018a6585930000b5979301, /*  289 */
128'h60e26442e495e04ae822ec0600074483, /*  290 */
128'h61058da505130000a51785aa690264a2, /*  291 */
128'h0000a51785aafab71ce327055940406f, /*  292 */
128'hfff7471301071733577db7f58c450513, /*  293 */
128'h03b6869b02e505334729c10d44018d79, /*  294 */
128'h746301045433942a472500d414334405, /*  295 */
128'h870505130000a51785be078514590087, /*  296 */
128'h05130000a51785a2c801542040ef8932, /*  297 */
128'h690285a6864a60e26442532040ef8665, /*  298 */
128'h5180406f610586e505130000a51764a2, /*  299 */
128'hf54ef94ae1a202c7073b8cbafce67155, /*  300 */
128'he162e55ee95aed56f152fd26e586f8ea, /*  301 */
128'hf66384368d3289ae892a04000793f4ee, /*  302 */
128'h4cc1000c956302ccdcbb04000c9300e7, /*  303 */
128'h001a849b020d1a13001d1a9b03acdcbb, /*  304 */
128'h00009b9781cb0b130000ab17020a5a13, /*  305 */
128'h4501e00d6dcc0c1300008c17784b8b93, /*  306 */
128'h6b4a6aea7a0a79aa794a74ea640e60ae, /*  307 */
128'h85ca808261697da67d467ce66c0a6baa, /*  308 */
128'h00040d9b47c040ef7d85051300009517, /*  309 */
128'h482146914781874e000c8d9b008cf463, /*  310 */
128'h9381020d979305b66b630007861b4889, /*  311 */
128'h083803bd06bb0d9de56399be034787b3, /*  312 */
128'h0b079c630006881b02e0089385ba4781, /*  313 */
128'h8c23e036794505130000951797ba1098, /*  314 */
128'h9281168241b4043b6682422040effa07, /*  315 */
128'h02dd1963b79d557dd13d0e2070ef9936, /*  316 */
128'h1602c19095aa26010828002795934310, /*  317 */
128'h67023ea040efe03ae43e855a85d69201, /*  318 */
128'h1963bf9d4691482107859752488967a2, /*  319 */
128'hbfd1e19095aa0828003795936310010d, /*  320 */
128'h164208280017959300075603011d1d63, /*  321 */
128'h082c00074603bf6d00c5902395aa9241, /*  322 */
128'he03e855eb76500c580230ff6761395be, /*  323 */
128'hbf253cfdfe97eae32785678210e070ef, /*  324 */
128'h0005450300cc053300074603bfdd4781, /*  325 */
128'h54634186561b0186161bc51909757513, /*  326 */
128'h87aa1582b70d07052785011700230006, /*  327 */
128'h8f8d25058082e21c00b7f46345019181, /*  328 */
128'h0088458189aa04000613fd4e7115bfd5, /*  329 */
128'hed5ef15af556f952e1cae5a6e9a2ed86, /*  330 */
128'h07130000a71767869982e16ae566e962, /*  331 */
128'h440106e79d63450983e107e263185be7, /*  332 */
128'h9b9766ab0b1300009b174a8503800a13, /*  333 */
128'h9d1708000cb780000c376a2b8b930000, /*  334 */
128'h450100f464630781578367ad0d130000, /*  335 */
128'h9dbd0028038006137786028a05bba091, /*  336 */
128'h855a85a2cfbd77c20957926347a29982, /*  337 */
128'h018487b374820409086379222b4040ef, /*  338 */
128'h40ef61a505130000951785a60397e863, /*  339 */
128'h7a4a79ea690e64ae644e60ee450d2960, /*  340 */
128'h8082612d6d0a6caa6c4a6bea7b0a7aaa, /*  341 */
128'h061b45c226c040ef856a86ca85a66642, /*  342 */
128'h79020097ff6377a274c2998285260009, /*  343 */
128'h862624a040ef855e85ca993e86268c9d, /*  344 */
128'h057e4505bfb12405060060ef854a4581, /*  345 */
128'h780707130000a7178082400005378082, /*  346 */
128'he30895360017869300756513157d631c, /*  347 */
128'h67858082953e057e450597aa20000537, /*  348 */
128'h871308a74463862a0ce5076382078713, /*  349 */
128'h496306e60b635c650513000095178087, /*  350 */
128'hc3ad5a250513000095178006079b04c7, /*  351 */
128'hc963622505130000951787f787936785, /*  352 */
128'h000095979e3d11417c07879b77fd04c7, /*  353 */
128'h40efe4066e4505130000a51761458593, /*  354 */
128'h808201416d4505130000a51760a21820, /*  355 */
128'h00e60a63574505130000951781078713, /*  356 */
128'hfaf612e3574505130000951781878793, /*  357 */
128'h09e35925051300009517830787138082, /*  358 */
128'h0513000095178287879300c74963fee6, /*  359 */
128'h580505130000951783878713bfe956e5, /*  360 */
128'h580505130000951784078793fce608e3, /*  361 */
128'hf022717980825365051300009517bf75, /*  362 */
128'h07bb00a5893b440184aaf406e84aec26, /*  363 */
128'h942a904114420104551302f044634099, /*  364 */
128'h1542fff54513740270a2952201045513, /*  365 */
128'h0068460985a6808261459141694264e2, /*  366 */
128'h979b0087d71b048900c15783753050ef, /*  367 */
128'hbf45943e93c117c200f117238fd90087, /*  368 */
128'h8793f44ef84afc26e486e0a26785715d, /*  369 */
128'h0e636dd7879367a13cf50463842e8067, /*  370 */
128'h082884b205e9440799638005079b0af5, /*  371 */
128'ha517461985ca00640913701050ef4611, /*  372 */
128'h0793017445836ed050ef5d2505130000, /*  373 */
128'h1cf5816347b108b7e76332f5886302e0, /*  374 */
128'h478502b7e3631af58263479104b7e563, /*  375 */
128'h83634ba5051300009517478910f58463, /*  376 */
128'ha41503a040ef656505130000951702f5, /*  377 */
128'h4c0505130000951747a118f581634799, /*  378 */
128'h2cf5816347f5a429020040effef591e3, /*  379 */
128'h0000951747d916f5896347c500b7ed63, /*  380 */
128'h856302100793bf6dfef580e34dc50513, /*  381 */
128'h051300009517faf596e3029007932af5, /*  382 */
128'h04b7e2632cf5816306200793b7c94f65, /*  383 */
128'h02f0079300b7ef632af5816303300793, /*  384 */
128'h4f850513000095170320079328f58663, /*  385 */
128'h079328f5836305c00793b7bdf8f58ae3, /*  386 */
128'hbf91f6f58de350e505130000951705e0, /*  387 */
128'h0670079300b7ef6328f5856308400793, /*  388 */
128'h520505130000951706c0079326f58a63, /*  389 */
128'h079326f5876308900793b73df4f58ae3, /*  390 */
128'h9517f0f59ce30880079326f588630ff0, /*  391 */
128'h0000a79701e45703b73d52a505130000, /*  392 */
128'h12f713634dc989930000a9974e47d783, /*  393 */
128'h10f71b634ce7d7830000a79702045703, /*  394 */
128'h0000a597461958d050ef852285ca4619, /*  395 */
128'h012301a4578357d050ef854a49c58593, /*  396 */
128'h859b01c4578300f41f23020412230204, /*  397 */
128'h1d230009d78302f4102302240513fde4, /*  398 */
128'h579bdb3ff0ef00f41e230029d78300f4, /*  399 */
128'h862602a4122300a11e238d5d05220085, /*  400 */
128'h051300009517a06ddcdfe0ef450185a2, /*  401 */
128'h9517b56133c5051300009517bd4932e5, /*  402 */
128'h0264470302444783bdbd34a505130000, /*  403 */
128'h01c1178300f10e230254478300f10ea3, /*  404 */
128'h470300e10e2327810274470300e10ea3, /*  405 */
128'h0e230234470300e10ea301c119030224, /*  406 */
128'ha79704e79b6301c156830450071300e1, /*  407 */
128'h85930000a597461947e23ad79f230000, /*  408 */
128'h2f230000a71739e505130000a5173965, /*  409 */
128'h0000a79766a2476249f050efe43638f7, /*  410 */
128'h60ef450102a40593ff89061b37478793, /*  411 */
128'h8082616179a2794274e2640660a65900, /*  412 */
128'h2f230000a71747e204e6946304300713, /*  413 */
128'ha797c799439c362787930000a79734f7, /*  414 */
128'h86930000a697f7e9439c352787930000, /*  415 */
128'h85930000a597342606130000a6173466, /*  416 */
128'h4d200713b765d73fe0ef02a405133465, /*  417 */
128'h5a9030ef264505130000951702e79863, /*  418 */
128'h2605051300009517ccaff0ef852285a6, /*  419 */
128'hbf95cb4ff0ef02a4051385ca595030ef, /*  420 */
128'h17fd67c101e45703f6e787e35fe00713, /*  421 */
128'ha5974611f4f70de302045703f6f701e3, /*  422 */
128'h9517b7993cb050ef0868302585930000, /*  423 */
128'h2405051300009517b33d23a505130000, /*  424 */
128'h00009517bb292565051300009517b315, /*  425 */
128'hb31927a5051300009517bb0126450513, /*  426 */
128'h051300009517b9f52805051300009517, /*  427 */
128'h9517b1e52ac5051300009517b9cd29e5, /*  428 */
128'h2e85051300009517b9f92c2505130000, /*  429 */
128'h0265d703b1e92f65051300009517b9d1, /*  430 */
128'h278484930000a4972807d7830000a797, /*  431 */
128'h26a7d7830000a7970285d703ecf711e3, /*  432 */
128'h016589930205891320000793eaf719e3, /*  433 */
128'h4619319050ef854a85ce461900f59a23, /*  434 */
128'h4619309050ef854e228585930000a597, /*  435 */
128'h2f7050ef00640513218585930000a597, /*  436 */
128'h061301c457832ed050ef852285ca4619, /*  437 */
128'hd78302f4142301e4578302f4132302a0, /*  438 */
128'h079300f41f230024d78300f41e230004, /*  439 */
128'h05130000951785aab36900f416236080, /*  440 */
128'hb603300017b7bba54601443030ef27e5, /*  441 */
128'h00f674132601608130239f0101138307, /*  442 */
128'h879b0387f5930034179b66858387b703, /*  443 */
128'h5e913c23639c97ae300005b79fad8406, /*  444 */
128'h849b5f200513fee7881b278160113423, /*  445 */
128'h00c5163b101005138a1d09056c63ffc7, /*  446 */
128'h07130000a717c34927018f71fff74713, /*  447 */
128'h871b700776130084171beb3d431814e7, /*  448 */
128'h969b00d100a345d495ba070e9f318006, /*  449 */
128'h550300d100230086d69b0106d69b0106, /*  450 */
128'h1e63806686936685c6918005069b0001, /*  451 */
128'h30000837860a27850077e79337ed02d5, /*  452 */
128'h983a00369813974285b246814037d79b, /*  453 */
128'h0006881bff063c230621068500083803, /*  454 */
128'h300017b70405a9bff0ef8626fef845e3, /*  455 */
128'h3483852660013403608130838287b823, /*  456 */
128'he8220c2007b711018082610101135f81, /*  457 */
128'hb703300014b747812401ec06e42643c0, /*  458 */
128'h00009517e7990206c163033716938304, /*  459 */
128'h60e2c3c00c2007b7311030ef16450513, /*  460 */
128'hbfc14785ec3ff0ef8082610564a26442, /*  461 */
128'h0000a597461184ae8432ec26f0227179, /*  462 */
128'h0000a79714b050eff406006808458593, /*  463 */
128'ha89785a6862247b20007a80303c78793, /*  464 */
128'h0693026757030000a717022888930000, /*  465 */
128'h85228e0ff0ef02e505130000a5170450, /*  466 */
128'h05220085579b8082614564e2740270a2, /*  467 */
128'h0185579b0185171b8082914115428d5d, /*  468 */
128'h8fd98f750085571bf00686938fd966c1, /*  469 */
128'h808225018d5d8d7900ff07370085151b, /*  470 */
128'h4585460100740207879b070007b7715d, /*  471 */
128'hf052f44ef84afc26e0a2e48604b00513, /*  472 */
128'h0513000095178a2a071070efc63eec56, /*  473 */
128'h89930000a9975ae14401233030ef09e5, /*  474 */
128'h028a863b44990969091300009917fa69, /*  475 */
128'h0286061b0405854a0004059b013407b3, /*  476 */
128'h1f9030ef00c780230ff6761300ca5633, /*  477 */
128'h0048f6c585930000a5974611fc941ee3, /*  478 */
128'h0028f5a585930000a5974609053050ef, /*  479 */
128'h010006374722f43ff0ef4512043050ef, /*  480 */
128'h0ff777138ff183210087179bf0060613, /*  481 */
128'h80a6b02317c29101300016b78fd91502, /*  482 */
128'h60a68086b7838006b78380f6b42393c1, /*  483 */
128'h7a0279a2794274e282f6b42347a16406, /*  484 */
128'hb5838007b603300017b7808261616ae2, /*  485 */
128'hfc068f4d91c115c20080073771398087, /*  486 */
128'hb423e05ae456e852ec4ef04af426f822, /*  487 */
128'ha71714b030effde505130000951780e7, /*  488 */
128'ha817ebe7c7830000a797ec5747030000, /*  489 */
128'ha617eac6c6830000a697eb7848030000, /*  490 */
128'h9517e9a5c5830000a597ea3646030000, /*  491 */
128'h04130000a41710f030effb2505130000, /*  492 */
128'he60989930000a997448100044783e864, /*  493 */
128'h0000aa1700144783e6f70c230000a717, /*  494 */
128'h4783e6f701a30000a7176a89e54a0a13, /*  495 */
128'h08230000a7173000193700262b370024, /*  496 */
128'h4783e4f702a30000a71700344783e4f7, /*  497 */
128'ha71700544783e2f70d230000a7170044, /*  498 */
128'ha797e00793230000a797e2f707a30000, /*  499 */
128'ha797e007a1230000a797de07ad230000, /*  500 */
128'he4a9de07a5230000a797de07ab230000, /*  501 */
128'h5a0b0493f23fe0ef8522e78d0009a783, /*  502 */
128'h83093783020745630337971383093783, /*  503 */
128'h2783bfc5c13ff0effc075de303379713, /*  504 */
128'h710a849300a060ef4501dff154fd000a, /*  505 */
128'h300017b7b7d914fdb7e9bf9ff0efbfc1, /*  506 */
128'h8f75e40616fd1141ff8006b78087b703, /*  507 */
128'hb58382e7b823f0070713670580e7b423, /*  508 */
128'h95177fa030efece50513000095178307, /*  509 */
128'h6709300027f37ee030efeea505130000, /*  510 */
128'h907307fe4785300790738fd988070713, /*  511 */
128'h100f7ca030efee650513000095173417, /*  512 */
128'h8082014160a2302000730ff0000f0000, /*  513 */
128'h002547838f5d07a20005470300154783, /*  514 */
128'h808225018d5d05628fd907c200354503, /*  515 */
128'h00f58733808200e613630007871b4781, /*  516 */
128'hb7d500d70023078500f5073300074683, /*  517 */
128'h0fa30505808200f613630005079b9e29, /*  518 */
128'he04ae426ec06e8221101495cbfc5feb5, /*  519 */
128'h02000613478101853903cfb500958413, /*  520 */
128'h470300f9073346ad02e0089348214515, /*  521 */
128'h831b0e50071300a7146302c700630007, /*  522 */
128'h00e40023040501140023010315630007, /*  523 */
128'h01c9051300b94783fcd79be307850405, /*  524 */
128'h01994783c088f4bff0ef00f5842384ae, /*  525 */
128'h478300f492238fd90087979b01894703, /*  526 */
128'h00f493238fd90087979b016947030179, /*  527 */
128'h80826105690264a2644260e200040023, /*  528 */
128'h468303a0061302000593cf99873e611c, /*  529 */
128'h06630017869300c6986302d5fc630007, /*  530 */
128'h46050007c683b7dd0705a00d577d00d7, /*  531 */
128'h078900b666630ff6f593fd06869b577d, /*  532 */
128'h47030000a7178082853ae11c0006871b, /*  533 */
128'hc70d0007c703cb85611cc915bfd5c2e7, /*  534 */
128'he406114102e69063008557030067d683, /*  535 */
128'hc3914501001577933b8060ef0017c503, /*  536 */
128'h01b5c783808245258082014160a24525, /*  537 */
128'h0006879b8edd0087979b470d01a5c683, /*  538 */
128'h0087179b0145c6030155c70300e51d63, /*  539 */
128'h71798082853e27818fd50107979b8fd1, /*  540 */
128'h0993e052e84af4065904e44eec26f022, /*  541 */
128'h60ef85ce8626468500154503842a0345, /*  542 */
128'h87bb000402234c58505ce13125013460, /*  543 */
128'h694264e2740270a2450100e7eb6340f4, /*  544 */
128'h74e34a0500344903808261456a0269a2, /*  545 */
128'h85ce86269cbd4685001445034c5cff2a, /*  546 */
128'h00454783b7f94505b7e5397d304060ef, /*  547 */
128'he8221101591c80824501f8dff06fc399, /*  548 */
128'h892e84aa02b787634401e04ae426ec06, /*  549 */
128'h46850014c503ec190005041bfddff0ef, /*  550 */
128'h4405c119250128c060ef03448593864a, /*  551 */
128'h690264a2644260e285220324a823597d, /*  552 */
128'h57fde04ae426ec06e822110180826105, /*  553 */
128'he52d2501fa3ff0ef842ad91c00050223, /*  554 */
128'h8fd90087979b45092324470323344783, /*  555 */
128'h9f63a55707134107d79b776d0107979b, /*  556 */
128'h05370005079bd4bff0ef06a4051302e7, /*  557 */
128'hf7b31465049300544537fff509130100, /*  558 */
128'hd25ff0ef0864051300978c6345010127, /*  559 */
128'h644260e200a035338d05012575332501, /*  560 */
128'hf84a715dbfcd450d80826105690264a2, /*  561 */
128'h00053023ec56f052fc26e0a2e486f44e, /*  562 */
128'h02054e6347adddbff0ef8932852e89aa, /*  563 */
128'h638097baa34787930000a79700351713, /*  564 */
128'hc79d000447830089b023c01547b184aa, /*  565 */
128'h0563e385001577931d8060ef00144503, /*  566 */
128'h794274e2640660a647a9c11189110009, /*  567 */
128'h0ff4f51380826161853e6ae27a0279a2, /*  568 */
128'h001577130ec060ef00a400a300040023, /*  569 */
128'h85224581f571891100090463fb79478d, /*  570 */
128'h1fa40913848a04f51a634785ee5ff0ef, /*  571 */
128'h854ac7894501ffc9478389a623a40a13, /*  572 */
128'h14e30991094100a9a0232501c51ff0ef, /*  573 */
128'h000a076345090004aa0301048913ff2a, /*  574 */
128'hfe9915e30491c10dea1ff0ef852285d2, /*  575 */
128'h05e34785470dbf8500e519634785470d, /*  576 */
128'h470304044783b78547b5c1194a01f6e5, /*  577 */
128'h4107d79b0107979b8fd90087979b03f4, /*  578 */
128'h04a4478304b44983fee791e320000713, /*  579 */
128'h448329811a09876300f9e9b30089999b, /*  580 */
128'h009401a3fff4879b470501342e230444, /*  581 */
128'h0124012304144903faf769e30ff7f793, /*  582 */
128'hffc100f977b3fff9079b2901fa0903e3, /*  583 */
128'h00faeab3008a9a9b0454478304644a83, /*  584 */
128'h478304844503ffbd00faf79301541423, /*  585 */
128'h0434478314050e638d5d0085151b0474, /*  586 */
128'h86bbdfa98fd90087979b250104244703, /*  587 */
128'h873200d7063b9f3d004ad71b27810334, /*  588 */
128'h6ce384ae032655bb40c5063bf4c563e3, /*  589 */
128'h1955694100b67763490516556605f326, /*  590 */
128'h014787bb24890147073b090900b93933, /*  591 */
128'h10e91163470dd05c03442023cc04d458, /*  592 */
128'h949bd408b09ff0ef06040513f00a93e3, /*  593 */
128'h57fdee99e6e30094d49b1ff4849b0024, /*  594 */
128'h1963478d00f402a3f8000793c45cc81c, /*  595 */
128'h8fd90087979b064447030654478308f9, /*  596 */
128'h059b06e79b6347054107d79b0107979b, /*  597 */
128'h23344783e13d2501ce7ff0ef8522001a, /*  598 */
128'h979b8fd90087979b000402a323244703, /*  599 */
128'h04e79263a55707134107d79b776d0107, /*  600 */
128'h87932501416157b7a8dff0ef03440513, /*  601 */
128'h77b7a77ff0ef2184051302f517632527, /*  602 */
128'h21c4051300f51c632727879325016141, /*  603 */
128'hc448a57ff0ef22040513c808a61ff0ef, /*  604 */
128'h971793c117c227857ba7d78300009797, /*  605 */
128'h2a230124002300f413237af716230000, /*  606 */
128'h099ba27ff0ef05840513b35147810004, /*  607 */
128'h84e3b545a19ff0ef05440513b5b10005, /*  608 */
128'h0014949b00f915634789d41c9fb5e00a, /*  609 */
128'h9cbd0017d79b8885029787bb478db709, /*  610 */
128'hc01ff0ef842ae426ec06e8221101bdcd, /*  611 */
128'h47030cf71063478d00044703ed692501, /*  612 */
128'h20000613034404930af71b6347850054, /*  613 */
128'h22f40923055007939fdff0ef85264581, /*  614 */
128'h02f40a230520079322f409a3faa00793, /*  615 */
128'h20f40da302f40b230610079302f40aa3, /*  616 */
128'h971b20e40d2302e40ba304100713481c, /*  617 */
128'h0ea320f40e230087571b0107571b0107, /*  618 */
128'h445c20f40fa30187d79b0107d71b20e4, /*  619 */
128'h571b0107571b0107971b501020e40f23, /*  620 */
128'h00a322f4002307200693001445030087, /*  621 */
128'h20d40c230187d79b0107d71b260522e4, /*  622 */
128'h4685d81022f401a322e4012320d40ca3, /*  623 */
128'h460100144503000402a3633050ef85a6, /*  624 */
128'h644260e200a035332501627050ef4581, /*  625 */
128'h377985beffe5879b4d188082610564a2, /*  626 */
128'h9d3d02b787bb55480025478300e7f963, /*  627 */
128'h71794d180eb7f5634785808245018082, /*  628 */
128'h02e5f963892ae44eec26f022f406e84a, /*  629 */
128'h0d63468d06d70b63842e468900054703, /*  630 */
128'hd59b9cad515c0015d49b00f71e6308d7, /*  631 */
128'h70a257fdc9112501ac7ff0ef9dbd0094, /*  632 */
128'h278380826145853e69a2694264e27402, /*  633 */
128'h94ca1ff4f4930099d59b0014899b0249, /*  634 */
128'hf5792501a93ff0ef0344c483854a9dbd, /*  635 */
128'h0087979b880503494783994e1ff9f993, /*  636 */
128'h515cbf4d93d117d2bf658391c0198fc5, /*  637 */
128'h141bf1452501a65ff0ef9dbd0085d59b, /*  638 */
128'h034945030359478399221fe474130014, /*  639 */
128'h9dbd0075d59b515cb7618fc90087979b, /*  640 */
128'h1fc575130024151bf93d2501a3bff0ef, /*  641 */
128'h024557931512ffaff0ef954a03450513, /*  642 */
128'hf04a4544f42671398082853e4785bfb9, /*  643 */
128'h478500b51523e456e852ec4ef822fc06, /*  644 */
128'h790274a2744270e2450900f49c63892a, /*  645 */
128'hf4e34f98611c808261216aa26a4269e2, /*  646 */
128'h00e69463470d0007c683e0a9842efee4, /*  647 */
128'h28235788fce477e30087d703eb0d5798, /*  648 */
128'h378300f92a239fa90044579bd1710099, /*  649 */
128'h00893c23943e034787930416883d0009, /*  650 */
128'h09924a855a7d0027c98384bab75d4501, /*  651 */
128'h2501e5dff0ef0134766385a600093503, /*  652 */
128'hfce301448c630005049be75ff0efbf7d, /*  653 */
128'h4134043bf6f4f7e34f9c00093783f69a, /*  654 */
128'he426e822110100a55583b7954505bfc1, /*  655 */
128'h484ce4950005049bf35ff0ef842aec06, /*  656 */
128'h06136c08ec990005049b939ff0ef6008, /*  657 */
128'h00e7802357156c1cf3cff0ef45810200, /*  658 */
128'h64a28526644260e200e782234705601c, /*  659 */
128'hf426f822fc06e852ec4e713980826105, /*  660 */
128'h84aa4d1c0ab9f5634a094985e456f04a, /*  661 */
128'h842e89324709000547830af5f0634a09, /*  662 */
128'hd99b093794630ee78863470d0ae78f63, /*  663 */
128'hf0ef9dbd0099d59b00b989bb515c0015, /*  664 */
128'h00198a9b8805060a166300050a1b8bdf, /*  665 */
128'hc783013487b3cc191ff9f9930ff97793, /*  666 */
128'h8ff50049179b00f7f71316c166850347, /*  667 */
128'h8223478502f98a2399a60ff7f7938fd9, /*  668 */
128'h86fff0ef9dbd8526009ad59b50dc00f4, /*  669 */
128'h591bc40d1ffafa93000a1f6300050a1b, /*  670 */
128'h82234785032a8a239aa60ff979130049, /*  671 */
128'h6a4269e2790274a28552744270e200f4, /*  672 */
128'h591b0347c783015487b3808261216aa2, /*  673 */
128'h515cb7e90127e9339bc100f979130089, /*  674 */
128'h12e300050a1b815ff0ef9dbd0085d59b, /*  675 */
128'h03240a2394261fe474130014141bfc0a, /*  676 */
128'h03240aa30089591b0109591b0109191b, /*  677 */
128'hf0ef9dbd0075d59b515cbf7901348223, /*  678 */
128'h74130024141bf80a16e300050a1bfdcf, /*  679 */
128'h2501d96ff0ef85569aa603440a931fc4, /*  680 */
128'h0109179b2901012569338d71f0000637, /*  681 */
128'h80a30087d79b03240a230107d79b9426, /*  682 */
128'h81a300fa81230189591b0109579b00fa, /*  683 */
128'hf04af822fc06ec4ef4267139bf79012a, /*  684 */
128'h056300c52903e99189ae84aae456e852, /*  685 */
128'hc5bff0efa815490502f96d634d1c0009, /*  686 */
128'h70e2852244050087ed6347850005041b, /*  687 */
128'h808261216aa26a4269e2790274a27442, /*  688 */
128'h844afef461e3894e4c9c08f4026357fd, /*  689 */
128'h012a646300f4676324054c9c5afd4a05, /*  690 */
128'h2501c0dff0ef852685a24409b7e94401, /*  691 */
128'hb7cdfd241de3fb450ae305550a63c901, /*  692 */
128'h2501debff0ef852685a2167d10000637, /*  693 */
128'hf8e788e3577dc4c0489c02099063e905, /*  694 */
128'h00f482a30017e7930054c783c89c37fd, /*  695 */
128'hdd612501dbdff0ef852685ce8622bfb5, /*  696 */
128'h5903f04a7139b795547df6f514e34785, /*  697 */
128'hec4ef426030917932905f822fc0600a5, /*  698 */
128'h74a2744270e24511eb9993c1e456e852, /*  699 */
128'hd7ed495c808261216aa26a4269e27902, /*  700 */
128'h2785480c00099d63842a8a2e00f97993, /*  701 */
128'h75e30009071b00855783e18dc85c6108, /*  702 */
128'h97ce03478793012415230996601cfcf7, /*  703 */
128'h37fd00495a9b00254783bf5d4501ec1c, /*  704 */
128'h0005049bb2fff0effc0a9fe30157fab3, /*  705 */
128'h00f4946357fdbf4945090097e4634785, /*  706 */
128'hf60a0ee306f4e0634d1c6008b7614505, /*  707 */
128'h4785d4bd451d0005049be83ff0ef480c, /*  708 */
128'hde0ff0ef6008fcf48de357fdfcf48be3, /*  709 */
128'h034505134581200006136008f5792501, /*  710 */
128'haabff0ef855285a600043a03bf0ff0ef, /*  711 */
128'h00faed630025478360084a0502aa2823, /*  712 */
128'hf0ef85a6c8046008d91c415787bb591c, /*  713 */
128'h2501d24ff0ef01450223b7b9c848a89f, /*  714 */
128'h7139b7e9db1c27855b1c2a856018f141, /*  715 */
128'he05ae456e852ec4ef04afc06f426f822, /*  716 */
128'h00e78663842e84aa02f007130005c783, /*  717 */
128'h47030004a62304050ce7946305c00713, /*  718 */
128'h05c00a9302f00a130ce7f06347fd0004, /*  719 */
128'h84630d478663000447834b2102e00993, /*  720 */
128'hf0ef854a02000593462d0204b9030d57, /*  721 */
128'h4783013900230d37966300044783b42f, /*  722 */
128'h478300f900a302e007930b3794630014, /*  723 */
128'h0793943a09479b63470d1d3789630024, /*  724 */
128'h2501adfff0ef8526458100f905a30200, /*  725 */
128'h2501ce0ff0ef608848cc492d10051963, /*  726 */
128'h478312078063000747836c9810051163, /*  727 */
128'h8633078500f706b3708cef898ba100b7, /*  728 */
128'h45810cd60a63fff646030006c68300f5, /*  729 */
128'h4bdc611ca0e1dd5d2501df9ff0ef8526, /*  730 */
128'hbc232501a81ff0ef85264581bf35c55c, /*  731 */
128'h6aa26a4269e2790274a2744270e20004, /*  732 */
128'h87e3b7b54709b73d0405808261216b02, /*  733 */
128'h02400793943a12f6e76302000693f757, /*  734 */
128'h48e502000313478145a147014681b78d, /*  735 */
128'h9101020695130027e793a2110505a8c9, /*  736 */
128'h051392011602a865268500e50023954a, /*  737 */
128'h4683c6e5460100e57363461194320200, /*  738 */
128'h00e90023471500e695630e5007130009, /*  739 */
128'h47118bb10ff7f7930027979b01659f63, /*  740 */
128'hf713bded00c905a30086661300e79463, /*  741 */
128'h9de3b7c501066613fed714e346850037, /*  742 */
128'hf4e513e34711c51500b7c783709cf127, /*  743 */
128'hbc230004a623cb990207f7930047f713, /*  744 */
128'hf315bfd94511b72d4501e6070ae30004, /*  745 */
128'h8bc100b5c7836c8cfbe58b91b7054515, /*  746 */
128'hb5a1c4c8ae4ff0ef0007c503609cdbe5, /*  747 */
128'h45ad46a10ff7f7930027979b05659a63, /*  748 */
128'h000747039722930117020017061b8732, /*  749 */
128'hfd370ae3f35709e3f3470be3f2e37de3, /*  750 */
128'h00054c634185551b0187151b02b6f263, /*  751 */
128'h00080663000548030005051300008517, /*  752 */
128'h0ff57513fbf7051bb5754519ef0719e3, /*  753 */
128'heca8efe30ff57513f9f7051beea8f3e3, /*  754 */
128'hf0227179bdc10ff777130017e7933701, /*  755 */
128'h0913451184aef406842ae44ee84aec26, /*  756 */
128'hf0ef6008a0b1c90de199484c49bd0e50, /*  757 */
128'hc783c3210007c7036c1ce1292501aecf, /*  758 */
128'h8bfd033780630327026303f7f79300b7, /*  759 */
128'h740270a2450100979a630017b79317e1, /*  760 */
128'hf0ef852245818082614569a2694264e2, /*  761 */
128'hbfe54511b7cd00042a23d9452501bfdf, /*  762 */
128'h87dff0ef842ae426ec06e82245811101, /*  763 */
128'ha7eff0ef6008484c0e500493e50d2501, /*  764 */
128'hcb9900978d630007c7836c1ced092501, /*  765 */
128'h13634791dd792501bb7ff0ef85224585, /*  766 */
128'h11018082610564a2644260e2451d00f5, /*  767 */
128'h0005049bfa9ff0ef842aec06e426e822, /*  768 */
128'he0850005049ba34ff0ef6008484ce49d, /*  769 */
128'h6c08700c838ff0ef4581020006136c08, /*  770 */
128'h60e200e782234705601c80eff0ef462d, /*  771 */
128'h08b7f06347858082610564a285266442, /*  772 */
128'he052e44eec26f406e84af02271794d1c, /*  773 */
128'h852285ca59fd4a0506f5f063892e842a, /*  774 */
128'h740270a24501e8910005049bed6ff0ef, /*  775 */
128'h03448c63808261456a0269a2694264e2, /*  776 */
128'h25018abff0ef852285ca460103348c63, /*  777 */
128'h00544783c81c278501378a63481cfd71, /*  778 */
128'he7e30004891b4c1c00f402a30017e793, /*  779 */
128'h80824509bf4d4505bf5d4509bf65faf4, /*  780 */
128'hf0eff42ee432e82efc061028ec2a7139, /*  781 */
128'h050ec92787930000979704054263832f, /*  782 */
128'h676200070023c3196622631800a78733, /*  783 */
128'h4785cb114501e39897aa00070023c319, /*  784 */
128'h2501a02ff0ef0828080c460100f61863, /*  785 */
128'he122e5067175bfe5452d8082612170e2, /*  786 */
128'h16050c63e42eecd6f0d2f4cef8cafca6, /*  787 */
128'hf0ef1028002c8a7984aa893200053023, /*  788 */
128'hf0efe4be1028083c65a2e91d25019cef, /*  789 */
128'h01c977934519e011e11964062501b61f, /*  790 */
128'h00f517634791c11510078e6301f97993, /*  791 */
128'h74e6640a60aac9052501e7dff0ef1028, /*  792 */
128'h00b44783808261496ae67a0679a67946, /*  793 */
128'h7913fff9452100497793f3fd8bc5451d, /*  794 */
128'h7a220089e9936406a02108090a630089, /*  795 */
128'h00f40ca300f408a30210071304600793, /*  796 */
128'h00040b2300e40823000407a300040723, /*  797 */
128'h00040e23000405a300e40c2300040ba3, /*  798 */
128'h000a450300040fa300040f2300040ea3, /*  799 */
128'h00040da300040d234785f9bfe0ef85a2, /*  800 */
128'h00fa02230005091b00040aa300040a23, /*  801 */
128'he1fff0ef030a2a83855285ca02090363, /*  802 */
128'hf0ef0125262385d6397d7522fd212501, /*  803 */
128'h0209e993c3990089f793f139250180cf, /*  804 */
128'hd09c01348523f4800309278385a27922, /*  805 */
128'h0513c8c8f35fe0ef00094503000485a3, /*  806 */
128'h0004a623c88800695783daffe0ef01c4, /*  807 */
128'hbdf5450100f494230124b0230004ae23, /*  808 */
128'h16e30107f713451100b44783ee051de3, /*  809 */
128'h9ee3451d8b85fa0900e300297913ee07, /*  810 */
128'he8d2eccef8a27119bdd14525bf51ec07, /*  811 */
128'hf466f862fc5ee0daf0caf4a6fc86e4d6, /*  812 */
128'h8ab6e4328a2e842a0006a023ec6ef06a, /*  813 */
128'h00b44783000998630005099be85fe0ef, /*  814 */
128'h74a6854e744670e60007899bc39d6622, /*  815 */
128'h7ca27c427be26b066aa66a4669e67906, /*  816 */
128'h8c638b8500a44783808261096de27d02, /*  817 */
128'h7463893e40f907bb445c010429031607, /*  818 */
128'h0b131ff00c1320000b930006091b00f6, /*  819 */
128'h91631ff777934458fa090ae35cfd0304, /*  820 */
128'hfd3337fd0025478300975d1b60081207, /*  821 */
128'h47854848eb11020d19630ffd7d1301a7, /*  822 */
128'h4c0cbfb5498900f405a3478900a7ec63, /*  823 */
128'h05a3478501951763b7e52501bc6ff0ef, /*  824 */
128'he43e853e4c0c601ccc08b795498500f4, /*  825 */
128'h00a6083b000d061bd5792501b86ff0ef, /*  826 */
128'h0099549b0027c683072c7a6367a28dc2, /*  827 */
128'h0017c50341a684bb00e6f46300c4873b, /*  828 */
128'h4783f945250112c050ef85d2864286a6, /*  829 */
128'hfc6341b507bb4c48c3850407f79300a4, /*  830 */
128'h85da20000613910115020097951b0097, /*  831 */
128'h9381020497930094949bc3ffe0ef9552, /*  832 */
128'h000aa783c45c9fa54099093b445c9a3e, /*  833 */
128'h4703050601634c50bf3900faa0239fa5, /*  834 */
128'h85da46850017c503c30d0407771300a4, /*  835 */
128'h682200a44783f13125010f2050efe442, /*  836 */
128'hc50386424685601c00f40523fbf7f793, /*  837 */
128'h01b42e23f10d250109e050ef85da0017, /*  838 */
128'h746340bb873b1ff5f5930009049b444c, /*  839 */
128'h855295a28626030585930007049b0127, /*  840 */
128'hf0caf8a27119b585499dbf9dbb1fe0ef, /*  841 */
128'hf862fc5ee0daf4a6fc86e4d6e8d2ecce, /*  842 */
128'h89328a2e842a0006a023ec6ef06af466, /*  843 */
128'h4783000997630005099bca3fe0ef8ab6, /*  844 */
128'h74a6854e744670e60007899bc39d00b4, /*  845 */
128'h7ca27c427be26b066aa66a4669e67906, /*  846 */
128'h82638b8900a44783808261096de27d02, /*  847 */
128'h20000b9304f76e630127873b445c1a07, /*  848 */
128'h0409046344585cfd03040b131ff00c13, /*  849 */
128'h478300975d1b6008140794631ff77793, /*  850 */
128'h040d1a630ffd7d1301a7fd3337fd0025, /*  851 */
128'h478902e798634705cb914581485cef01, /*  852 */
128'h079bd6aff0ef4c0cb749498900f405a3, /*  853 */
128'h00a4478312f76b634818445cf3fd0005, /*  854 */
128'h478501979763b78500f405230207e793, /*  855 */
128'hc85ce311cc1c4858bf89498500f405a3, /*  856 */
128'h46854c50601cc38d0407f79300a44783, /*  857 */
128'h4783f969250178f040ef85da0017c503, /*  858 */
128'h853e4c0c601c00f40523fbf7f79300a4, /*  859 */
128'h063b000d081bd1592501964ff0efe43e, /*  860 */
128'h549b0027c683072c7a6367a28db200a8, /*  861 */
128'hc50341a684bb00e6f4630104873b0099, /*  862 */
128'h4c4cf149250173f040ef85d286a60017, /*  863 */
128'h918115820097959b0297f26341b587bb, /*  864 */
128'h00a44783a29fe0ef855a95d220000613, /*  865 */
128'h020497930094949b00f40523fbf7f793, /*  866 */
128'ha783c45c9fa54099093b445c9a3e9381, /*  867 */
128'h00c70e634c58bdc900faa0239fa5000a, /*  868 */
128'h85da46850017c50300d77a6344584814, /*  869 */
128'h049b444801b42e23fd0125016a3040ef, /*  870 */
128'h049b0127746340ab873b1ff575130009, /*  871 */
128'h9b5fe0ef952285d28626030505130007, /*  872 */
128'hc81cbf4100f405230407e79300a44783, /*  873 */
128'he0ef842ae406e0221141bd15499db5f1, /*  874 */
128'hcf610207f71300a44783e16d2501ab7f, /*  875 */
128'h0017c50346854c50601cc3950407f793, /*  876 */
128'h00a44783ed4d2501661040ef03040593, /*  877 */
128'hb5ffe0ef6008500c00f40523fbf7f793, /*  878 */
128'h85a30207671300b7c703741ce1552501, /*  879 */
128'h0086d69b0106d69b0107169b481800e7, /*  880 */
128'h0187571b0107569b00d78ea300e78e23, /*  881 */
128'h8ba300078b23485800e78fa300d78f23, /*  882 */
128'h8a230107571b0107169b00e78d230007, /*  883 */
128'h8aa30087571b0107571b0107171b00e7, /*  884 */
128'hd69b00e78c23021007130106d69b00e7, /*  885 */
128'h892300e78ca300d78da3046007130086, /*  886 */
128'hfdf7f793600800a44783000789a30007, /*  887 */
128'h014160a2640200f50223478500f40523, /*  888 */
128'h114180820141640260a24505ea3fe06f, /*  889 */
128'h8522e9012501f01ff0ef842ae406e022, /*  890 */
128'h640260a200043023e11925019b5fe0ef, /*  891 */
128'h945fe0efec060028e42a110180820141, /*  892 */
128'h60e245015aa78a230000879700054a63, /*  893 */
128'h002c4601e42a7159bfe5452d80826105, /*  894 */
128'h0005041bb25fe0efeca6f486f0a21028, /*  895 */
128'h041bcb4ff0efe4be1028083c65a2ec19, /*  896 */
128'h8522cbd8575277a2e9916586e41d0005, /*  897 */
128'h8bc100b5c7838082616564e6740670a6, /*  898 */
128'hb7c5c8c8965fe0ef0004c50374a2cb99, /*  899 */
128'he42afca67175bfd94415fcf41ee34791, /*  900 */
128'h460184ae00050023f4cef8cae122e506, /*  901 */
128'hecbe081ce5212501ab9fe0ef1828002c, /*  902 */
128'h91634996c2be4bdc02f00913842677e2, /*  903 */
128'h5007470300008717e50567a245010409, /*  904 */
128'h00e780a303a0071300e780230307071b, /*  905 */
128'h8023078d00e7812302f007130e941563, /*  906 */
128'h8082614979a6794674e6640a60aa0007, /*  907 */
128'h18284581fd4d2501f75fe0ef18284585, /*  908 */
128'h0007c50365c677e2f55d2501e6cff0ef, /*  909 */
128'h2501f4ffe0ef18284581c2aa8bdfe0ef, /*  910 */
128'h77e2e1052501e46ff0ef18284581f951, /*  911 */
128'h01350e632501897fe0ef0007c50365c6, /*  912 */
128'h67a24711dd612501a86ff0ef18284581, /*  913 */
128'hf48fe0ef1828100cb7614509f6e512e3, /*  914 */
128'hfc974703973610949301020797134781, /*  915 */
128'h36fd86a285be04e460630037871be705, /*  916 */
128'hfff7c793e989963a9301020697136622, /*  917 */
128'hfff5871bb7e12785bf199c3d01260023, /*  918 */
128'hfc974703972a1088930117020007059b, /*  919 */
128'h169367220789bdf54545b7e900e60023, /*  920 */
128'h8fa32405078500074703973692810204, /*  921 */
128'hf04af426f8227139b721fe9465e3fee7, /*  922 */
128'hfa8fe0ef84ae842ae456e852ec4efc06, /*  923 */
128'h891bcf8900b44783000917630005091b, /*  924 */
128'h6a4269e2790274a2854a744270e20007, /*  925 */
128'h00a44783009777634818808261216aa2, /*  926 */
128'h445ce4bd00042623445884bae3918b89, /*  927 */
128'h0207e79300a44783c81cfcf778e34818, /*  928 */
128'hd3e51ff7f793445c4481bf7d00f40523, /*  929 */
128'hf7930304099300a44783fc960ee34c50, /*  930 */
128'h40ef0017c50385ce4685601cc3850407, /*  931 */
128'h0523fbf7f79300a44783ed5125012f70, /*  932 */
128'h40ef85ce0017c50386264685601c00f4, /*  933 */
128'h002547836008bf59cc44ed3525012a50, /*  934 */
128'h0336d6bbfff4869b377dc7290097999b, /*  935 */
128'h4c0c8ff9413007bb02c6ed630337563b, /*  936 */
128'h0499ea634a855a7dd1c19c9dc45c2781, /*  937 */
128'he0ef6008d7b51ff4f793c45c9fa5445c, /*  938 */
128'h484cbfb19ca90094d49bcd112501c79f, /*  939 */
128'h00f5976347850005059b802ff0efe595, /*  940 */
128'h00f5976357fdbded490900f405a34789, /*  941 */
128'hb765cc0cc84cb5ed490500f405a34785, /*  942 */
128'h059bfcbfe0efcb818b89600800a44783, /*  943 */
128'h0005059bc3ffe0efbf6984cee5990005, /*  944 */
128'hfaf5fae34f9c601cfabafee3fd4588e3, /*  945 */
128'hb7bdc45c013787bb413484bbcc0c445c, /*  946 */
128'h002c4601842ac52de42ef822fc067139, /*  947 */
128'h852265a267e2e1152501fdafe0ef0828, /*  948 */
128'h6c0ce5292501968ff0eff01c101ce01c, /*  949 */
128'h000430234515e7898bc100b5c783cd99, /*  950 */
128'h67e2c448e24fe0ef0007c50367e2a02d, /*  951 */
128'hcadfe0ef00f414230067d78385224581, /*  952 */
128'h6121744270e2f971fcf50be347912501, /*  953 */
128'h1141b7c1fcf501e34791bfdd45258082, /*  954 */
128'h3023e1192501daefe0ef842ae406e022, /*  955 */
128'hec26f022717980820141640260a20004, /*  956 */
128'h0005049bd8cfe0ef892e842af406e84a, /*  957 */
128'h049bc4ffe0ef8522458100091f63e889, /*  958 */
128'h8082614564e269428526740270a20005, /*  959 */
128'h47912501b34ff0ef8522458102243023, /*  960 */
128'hc58fe0ef852285ca00042a2302f51363, /*  961 */
128'h00f5166347912501f77fe0ef85224581, /*  962 */
128'heca67159bf6584aad16dbf7d00042a23, /*  963 */
128'he0eff486f0a21028002c460184aee42a, /*  964 */
128'he4be1028083c65a2e00d0005041becef, /*  965 */
128'hc489cf816786e8010005041b85eff0ef, /*  966 */
128'h64e6740670a68522c00fe0ef102885a6, /*  967 */
128'hf85a8432f0a27159bfcd441980826165, /*  968 */
128'heca6f486e0d28522002c46018b2ee42a, /*  969 */
128'he70fe0efec66f062f45efc56e4cee8ca, /*  970 */
128'h481c01842c836000000a1c6300050a1b, /*  971 */
128'h740670a600fb202302f76263ffec871b, /*  972 */
128'h7ba27b427ae26a0669a6694664e68552, /*  973 */
128'h9f63478500044b83808261656ce27c02, /*  974 */
128'he0ef852285ca4a8559fd4481490902fb, /*  975 */
128'h2485e11109550863093508632501a49f, /*  976 */
128'he793c80400544783fef963e329054c1c, /*  977 */
128'h0ab7504cb74d009b202300f402a30017, /*  978 */
128'h00099e631afd4c094481498149011000, /*  979 */
128'h85cee9212501d04fe0ef0015899b8522, /*  980 */
128'h00194783038b91632000099303440913, /*  981 */
128'h09092485e3918fd90087979b00094703, /*  982 */
128'he0efe02e854ab745fc0c94e33cfd39f9, /*  983 */
128'h09112485e1116582015575332501aa2f, /*  984 */
128'hbfad8a2abfbd4a09b7494a05b7c539f1, /*  985 */
128'hbb8fe0ef842ae04aec06e426e8221101, /*  986 */
128'h0007849bcb9100b44783e4910005049b, /*  987 */
128'h47838082610564a269028526644260e2, /*  988 */
128'hfed772e348144458cf390027f71300a4, /*  989 */
128'h484cef01600800f40523c8180207e793, /*  990 */
128'h00a405a3c53900042a232501a5aff0ef, /*  991 */
128'h57fd0005091b941fe0ef4c0cbf7d84aa, /*  992 */
128'h167d100006374c0cb7dd450502f91463, /*  993 */
128'ha1eff0ef85ca6008f9792501b25fe0ef, /*  994 */
128'hfcf900e345094785b769449db7e12501, /*  995 */
128'h0407f79300a44783fcf96ae34d1c6008, /*  996 */
128'h030405930017c50346854c50601cdba5, /*  997 */
128'hfbf7f79300a44783f55d25016d4040ef, /*  998 */
128'h1008002c4605e42a7175b7b100f40523, /*  999 */
128'he9052501c94fe0eff8cafca6e122e506, /* 1000 */
128'he1052501e27fe0efe0be1008081c65a2, /* 1001 */
128'h75e2eb890207f79300b7c78345196786, /* 1002 */
128'h60aa451dcb810014f79300b5c483c599, /* 1003 */
128'h00094503790280826149794674e6640a, /* 1004 */
128'h2783c89d88c1cc0d0005041baccfe0ef, /* 1005 */
128'he0ef00a8100c02800613fc878de30149, /* 1006 */
128'hf1612501941fe0efcaa200a84589952f, /* 1007 */
128'h18e34791d94d2501838ff0ef00a84581, /* 1008 */
128'h7502e411f15525019e3fe0ef1008faf5, /* 1009 */
128'h91eff0ef85a27502bf612501f12fe0ef, /* 1010 */
128'h1028002c4605e42a7171b7edf5512501, /* 1011 */
128'hf8dafcd6e152e54ee94aed26f506f122, /* 1012 */
128'h0005041bbc4fe0efe8eaece6f0e2f4de, /* 1013 */
128'hd53fe0efe4be1028083c65a21c041263, /* 1014 */
128'h67a61af4156347911c0407630005041b, /* 1015 */
128'h752218079d630207f79300b7c7834419, /* 1016 */
128'h4785180480630005049bb33fe0ef4581, /* 1017 */
128'h16f48863440557fd16f48c6344097522, /* 1018 */
128'h85a67422160412630005041ba8cfe0ef, /* 1019 */
128'h061303440b13f60fe0ef85220104d91b, /* 1020 */
128'h462d886fe0ef855a00050c1b45812000, /* 1021 */
128'h0ff97a9347c187afe0ef855a02000593, /* 1022 */
128'h0109d99b02f40fa30109191b0104999b, /* 1023 */
128'h04f4062302e00b930109591b02100793, /* 1024 */
128'h0089591b0089d99b046007930ff4fa13, /* 1025 */
128'h0404052303740a230200061304f406a3, /* 1026 */
128'h05540423053407a305440723040405a3, /* 1027 */
128'h7722ff7fd0ef0544051385da052404a3, /* 1028 */
128'h00d6166357d200074603468d05740aa3, /* 1029 */
128'h0107969b06f40723478100f693635714, /* 1030 */
128'h0106d69b0107979b06f404230107d79b, /* 1031 */
128'h06d407a30087d79b0086d69b0107d79b, /* 1032 */
128'h1028040b99634c8500274b8306f404a3, /* 1033 */
128'h752247416786e8350005041bf5ffe0ef, /* 1034 */
128'h0460071300e78c230210071300e785a3, /* 1035 */
128'h01478d2300e78ca300078ba300078b23, /* 1036 */
128'h0223478501278aa301578a2301378da3, /* 1037 */
128'h0d1b7522a82d0005041bd50fe0ef00f5, /* 1038 */
128'h041b8d4fe0ef0195022303852823001c, /* 1039 */
128'hd0ef3bfd855a458120000613ec090005, /* 1040 */
128'h85a67522441db7498c6a0ffbfb93f53f, /* 1041 */
128'h69aa694a64ea740a70aa8522f2bfe0ef, /* 1042 */
128'h614d6d466ce67c067ba67b467ae66a0a, /* 1043 */
128'h84aee42aeca6f0a27159b7c544218082, /* 1044 */
128'h25019c2fe0eff48610284605002c8432, /* 1045 */
128'h2501b55fe0efe4be1028083c65a2e131, /* 1046 */
128'he39d0207f79300b7c783451967a6e915, /* 1047 */
128'h74138c658cbd752200b74783c30d6706, /* 1048 */
128'he0ef00f502234785008705a38c3d0274, /* 1049 */
128'h71718082616564e6740670a62501c94f, /* 1050 */
128'hed26f122f5060088002c4605e02ee42a, /* 1051 */
128'h65a26786120795630005079b95cfe0ef, /* 1052 */
128'h0005079bae7fe0eff0be083cf4be0088, /* 1053 */
128'h02077713479900b7c703778610079963, /* 1054 */
128'h05ad46550e058d63479165e610071163, /* 1055 */
128'hd0ef10a8008c02800613e3ffd0ef1028, /* 1056 */
128'h65820c054c6347adefdfd0ef850ae33f, /* 1057 */
128'h92634711cbf10005079ba9dfe0ef10a8, /* 1058 */
128'h648aebdd0005079bdcbfe0ef10a80ce7, /* 1059 */
128'h4783df7fd0ef00d4851302a10593464d, /* 1060 */
128'h0223478500f485a30207e79364060281, /* 1061 */
128'h076357d64736cbb58bc100b4c78300f4, /* 1062 */
128'h0005059bf25fd0ef85a60004450306f7, /* 1063 */
128'h8522c1bd47890005059bca4fe0ef8522, /* 1064 */
128'h02e007936706efa90005079bfbbfd0ef, /* 1065 */
128'h07230107969b57d602f69c6305574683, /* 1066 */
128'hd79b0107979b06f704230107d79b06f7, /* 1067 */
128'h04a30086d69b0106d69b0087d79b0107, /* 1068 */
128'he0ef008800f7022306d707a3478506f7, /* 1069 */
128'h079bb48fe0ef6506e7910005079be18f, /* 1070 */
128'h47a18082614d853e64ea740a70aa0005, /* 1071 */
128'h1028002c4605842ee42ae8a2711dbfcd, /* 1072 */
128'h1028083c65a2e929250180afe0efec86, /* 1073 */
128'hc783451967a6e129250199dfe0efe4be, /* 1074 */
128'h00645703cb856786eb950207f79300b7, /* 1075 */
128'h570300e78ba30087571b00e78b237522, /* 1076 */
128'h478500e78ca30087571b00e78c230044, /* 1077 */
128'h6125644660e62501acefe0ef00f50223, /* 1078 */
128'h002c893284aee42ae0cae4a6711d8082, /* 1079 */
128'h0005041bf95fd0efec86e8a208284601, /* 1080 */
128'h2501c9efe0efd20208284581c4b9e051, /* 1081 */
128'h75c2e93d2501b97fe0ef08284585e559, /* 1082 */
128'h061346ad00b48713c8dfd0ef8526462d, /* 1083 */
128'h0007869bfff6879bce89000700230200, /* 1084 */
128'hfec783e3177d0007c78397a693811782, /* 1085 */
128'h0005041be63fd0ef510c656202090a63, /* 1086 */
128'h84630005468304300793470d6562e015, /* 1087 */
128'hc15fd0ef953e034787930270079300e6, /* 1088 */
128'h6125690664a6644660e6852200a92023, /* 1089 */
128'h842abf550004802300f5156347918082, /* 1090 */
128'hec86e8a21028002c4605e42a711db7d5, /* 1091 */
128'h00010c236522e4710005041beddfd0ef, /* 1092 */
128'heb2900074703972a9301020797134781, /* 1093 */
128'hbccfe0efda0210284581ebb102000613, /* 1094 */
128'h2501ac3fe0ef10284585e0450005041b, /* 1095 */
128'h082c462dc7e565060181478310051563, /* 1096 */
128'h071300e78c23021007136786bb1fd0ef, /* 1097 */
128'ha0e900e78ca300078ba300078b230460, /* 1098 */
128'h02071693fff7871bb77d87bab7452785, /* 1099 */
128'h48e54701fec686e30006c68396aa9281, /* 1100 */
128'h96930017061b0006c58300e506b3432d, /* 1101 */
128'hec63030858131842f9f6881b92c10305, /* 1102 */
128'ha18585930000759792c116c236810108, /* 1103 */
128'h45e34185d59b0185959ba83100068e1b, /* 1104 */
128'h058580826125644660e685224419feb0, /* 1105 */
128'h02e3b7ddffc81be3000805630005c803, /* 1106 */
128'h0007069b00d58023070595ba082cfe67, /* 1107 */
128'h020006134729938102061793f8f6e9e3, /* 1108 */
128'h0e5007930181470300d779630007869b, /* 1109 */
128'h078500c6802396be0834b77df0f713e3, /* 1110 */
128'h00f502234785752200f500235795b7c5, /* 1111 */
128'h02f51b634791b7710005041b8b2fe0ef, /* 1112 */
128'h0005041ba19fe0ef1028d3c101814783, /* 1113 */
128'h6506ab7fd0ef4581020006136506f835, /* 1114 */
128'h00e785a347216786a8dfd0ef082c462d, /* 1115 */
128'h230305452e0305052e83bf81842abdd1, /* 1116 */
128'h8f2ae44ae826ec22110105c528830585, /* 1117 */
128'h00005f97887687f2869a864604050293, /* 1118 */
128'ha38300b647338dfd00c6c5b3514f8f93, /* 1119 */
128'h007585bb0fc1008fa403000f2583000f, /* 1120 */
128'h159b0105883b004f2703ff4fa3839db9, /* 1121 */
128'h05bb0077073b0105e8330198581b0078, /* 1122 */
128'h008f23838e358e6d00f6c6339f3100f8, /* 1123 */
128'h008383bb8e590146561b00c6171b9e39, /* 1124 */
128'h24038ef900b7c6b300d383bb00c5873b, /* 1125 */
128'h0116969b00f6d39b007686bb8ebd00cf, /* 1126 */
128'h061b00d703bbffcfa4039fa100d3e6b3, /* 1127 */
128'h579b9f3d8f2d9fa1007777338f2d0007, /* 1128 */
128'h869b0005881b0f418f5d0167171b00a7, /* 1129 */
128'h0f1300005f17f45f17e300e387bb0003, /* 1130 */
128'h82930000529748ef8f9300005f97556f, /* 1131 */
128'h000fa58300b6c7338df100d7c5b35562, /* 1132 */
128'h038a000f47039db9002f4403001f4383, /* 1133 */
128'ha7039db9942a040a4318972a070a93aa, /* 1134 */
128'h01b8581b9e390058159b0105883b004f, /* 1135 */
128'hc6339f3100f805bb0105e8330003a703, /* 1136 */
128'h0096139b008fa7039e398e3d8e7500b7, /* 1137 */
128'h00c583bb00c3e63340189eb90176561b, /* 1138 */
128'h8eadffff44838efd0075c6b30f119f35, /* 1139 */
128'h00e6941b94aa048affcfa7039eb90fc1, /* 1140 */
128'h9fb900d3843b8ec140980126d69b9fb9, /* 1141 */
128'h00c7579b9f3d007747338f6d0083c733, /* 1142 */
128'h069b0003861b0005881b8f5d0147171b, /* 1143 */
128'h8f9300005f97f25f1ee300e407bb0004, /* 1144 */
128'h0102c4033ec383930000539782fe476f, /* 1145 */
128'h00c5c4b3942a040a00d7c5b30003a703, /* 1146 */
128'h048a0043a4039f210112c4839f254000, /* 1147 */
128'h171b0122c4830107083b40809e2194aa, /* 1148 */
128'h0083a4039e210107683301c8581b0048, /* 1149 */
128'h40809e2d9ea194aa8db9048a00f8073b, /* 1150 */
128'h03c18e4d0156561b0132c90300b6159b, /* 1151 */
128'h8ead00e7c6b3ffc3a4839c3500c705bb, /* 1152 */
128'h0106d69b9fa50106941b992a9ea1090a, /* 1153 */
128'h8f2d0007081b00d5843b8ec100092483, /* 1154 */
128'h8f5d0177171b0097579b9f3d8f219fa5, /* 1155 */
128'h17e300e407bb0004069b0005861b0291, /* 1156 */
128'h8f5dfff6471336e2829300005297f45f, /* 1157 */
128'h022fc403021fc3830002a70300d745b3, /* 1158 */
128'h418c95aa058a93aa038a020fc5839f2d, /* 1159 */
128'h171b0107083b0042a5839f2d942a040a, /* 1160 */
128'h0107683301a8581b0003a5839e2d0068, /* 1161 */
128'h9e2d8e3d8e59fff6c6139db100f8073b, /* 1162 */
128'h400c9ead0166561b00a6139b0082a583, /* 1163 */
128'hc593023fc4839ead00c703bb00c3e633, /* 1164 */
128'h9db5ffc2a4038db902c10075e5b3fff7, /* 1165 */
128'h9fa18dd50115d59b94aa00f5969b048a, /* 1166 */
128'h8f4dfff747130007081b00b385bb4080, /* 1167 */
128'h0157171b00b7579b9f3d007747339fa1, /* 1168 */
128'h00e587bb0005869b0003861b0f918f5d, /* 1169 */
128'h06bb00fe07bb010e883b6462f3ff1de3, /* 1170 */
128'hcd70cd34c97c0505282300c8863b00d3, /* 1171 */
128'hfc26e0a2715d653c80826105692264c2, /* 1172 */
128'hf413ec56f052e486e45ee85af44ef84a, /* 1173 */
128'h04000b13e53c893289ae84aa97b203f7, /* 1174 */
128'h9381178200078a1b408b07bb04000b93, /* 1175 */
128'h020ada93020a1a9300090a1b00f97463, /* 1176 */
128'h4a7020ef0144043b86560084853385ce, /* 1177 */
128'h4401852660bc0174176399d641590933, /* 1178 */
128'h7a0279a2794274e2640660a6b7c99782, /* 1179 */
128'hf0227179653c808261616ba26b426ae2, /* 1180 */
128'h8513e84af406e44eec26842a03f7f793, /* 1181 */
128'h0400099300e7802397a2f80007130017, /* 1182 */
128'h4581920116020006091b40a9863b449d, /* 1183 */
128'hfc1c078e643c0124f5633f3020ef9522, /* 1184 */
128'h740270a2fd24fde3450197828522603c, /* 1185 */
128'h8793000077978082614569a2694264e2, /* 1186 */
128'h879300007797e93c04053423639c0567, /* 1187 */
128'he13cb807879300000797ed3c639c04e7, /* 1188 */
128'h20efec06850a46410505059311018082, /* 1189 */
128'h0000659732c686930000769747013e50, /* 1190 */
128'h06890007c78300e107b345414b458593, /* 1191 */
128'h97ae000646038bbd962e0047d6130705, /* 1192 */
128'hfca71de3fef68fa3fec68f230007c783, /* 1193 */
128'h7175808261052ee505130000751760e2, /* 1194 */
128'h6622f71ff0efe42ee5060808842ae122, /* 1195 */
128'h0808f01ff0ef0808e85ff0ef080885a2, /* 1196 */
128'h46a1595880826149640a60aaf83ff0ef, /* 1197 */
128'h0200071300d71763469100d70d63711c, /* 1198 */
128'h8082556dbfe50007ac2380824501cf98, /* 1199 */
128'h84ae842a200007b7ec06e426e8221101, /* 1200 */
128'h0880061311c686930000569702f50263, /* 1201 */
128'h42850513000065174185859300006597, /* 1202 */
128'h8082610564a2644260e2fc24189030ef, /* 1203 */
128'h84ae200007b7ec06e4266100e8221101, /* 1204 */
128'h02f006130f4686930000569702f40263, /* 1205 */
128'h3e850513000065173d85859300006597, /* 1206 */
128'h8082610564a2644260e2e004149030ef, /* 1207 */
128'h84ae200007b7ec06e4266100e8221101, /* 1208 */
128'h036006130c4686930000569702f40263, /* 1209 */
128'h3a850513000065173985859300006597, /* 1210 */
128'h8082610564a2644260e2e404109030ef, /* 1211 */
128'h842e200007b7ec06e8226104e4261101, /* 1212 */
128'h03e00613f1c686930000769702f48263, /* 1213 */
128'h36850513000065173585859300006597, /* 1214 */
128'h64a2644260e2e880900114020c9030ef, /* 1215 */
128'h07b7ec06e8226104e426110180826105, /* 1216 */
128'hed0686930000769702f48263842e2000, /* 1217 */
128'h00006517314585930000659704500613, /* 1218 */
128'h60e2ec8090011402085030ef32450513, /* 1219 */
128'he4266100e82211018082610564a26442, /* 1220 */
128'h0000569702f4026384ae200007b7ec06, /* 1221 */
128'h2d0585930000659704c0061300c68693, /* 1222 */
128'h60e2f004041030ef2e05051300006517, /* 1223 */
128'he4266100e82211018082610564a26442, /* 1224 */
128'h0000569702f4026384ae200007b7ec06, /* 1225 */
128'h290585930000659705300613fdc68693, /* 1226 */
128'h60e2f404001030ef2a05051300006517, /* 1227 */
128'h00053983ec4e71398082610564a26442, /* 1228 */
128'h893284ae200007b7fc06f04af426f822, /* 1229 */
128'h0613fa2686930000569702f984638436, /* 1230 */
128'h051300006517246585930000659705a0, /* 1231 */
128'h88090014141b67227b4030efe43a2565, /* 1232 */
128'h0034949b8c59004979130029191b8b05, /* 1233 */
128'h744270e20289b8238c4588a101246433, /* 1234 */
128'h7100e02211418082612169e2790274a2, /* 1235 */
128'hf7dff0efe40645818522460546814705, /* 1236 */
128'h4605468547058522f35ff0ef45818522, /* 1237 */
128'h60a2d97ff0ef45816008f67ff0ef4581, /* 1238 */
128'h4705e022e40611418082014145016402, /* 1239 */
128'h842a45810405302302053c2346054681, /* 1240 */
128'h45818522ef1ff0ef45818522f39ff0ef, /* 1241 */
128'h60a264026008f23ff0ef460546854705, /* 1242 */
128'he8226104e4261101d4dff06f01414581, /* 1243 */
128'h0000569702f48263842e200007b7ec06, /* 1244 */
128'h160585930000659706100613ecc68693, /* 1245 */
128'h904114426d0030ef1705051300006517, /* 1246 */
128'he42611018082610564a2644260e2fc80, /* 1247 */
128'h02f48263842e200007b7ec06e8226104, /* 1248 */
128'h0000659706800613e986869300005697, /* 1249 */
128'h68c030ef12c505130000651711c58593, /* 1250 */
128'h8082610564a2644260e2e0a090511452, /* 1251 */
128'h84ae200007b7ec06e4266100e8221101, /* 1252 */
128'h06f00613e64686930000569702f40263, /* 1253 */
128'h0e850513000065170d85859300006597, /* 1254 */
128'h8082610564a2644260e2e424648030ef, /* 1255 */
128'h07b7ec06e426e82200053903e04a1101, /* 1256 */
128'h86930000569702f9026384ae842a2000, /* 1257 */
128'h6517092585930000659707600613e2e6, /* 1258 */
128'hc84404993c23602030ef0a2505130000, /* 1259 */
128'hf0a2715980826105690264a2644260e2, /* 1260 */
128'hf85afc56e0d2e4cef486e8caeca67100, /* 1261 */
128'h892e0005d783020408a3ec66f062f45e, /* 1262 */
128'h20ef00c9051345814611d01ce03084b2, /* 1263 */
128'h3983bf7ff0ef458560080e049c636f60, /* 1264 */
128'h278316f99a6304043a03200007b70004, /* 1265 */
128'he391448d8b89c7090017f71344810049, /* 1266 */
128'h2783000a09638cdd03243c234c1c4485, /* 1267 */
128'h468147050144e493160786638b85008a, /* 1268 */
128'hf0ef85224581d73ff0ef852245814605, /* 1269 */
128'hc55ff0ef00989a37852200892583be3f, /* 1270 */
128'h85a6c8bff0ef681a0a13852200095583, /* 1271 */
128'h4705cffff0ef85224581cc7ff0ef8522, /* 1272 */
128'h000f45b7d31ff0ef8522458146054685, /* 1273 */
128'hf0ef85224585e9bff0ef852224058593, /* 1274 */
128'hd58c8c9300005c9785220d89b583cdbf, /* 1275 */
128'h8a9300006a97ebbff0ef25810015e593, /* 1276 */
128'h70a6efe9485cf7eb0b1300006b17f6ea, /* 1277 */
128'h7ba27b427ae26a0669a6694664e67406, /* 1278 */
128'he024852244cc8082616545016ce27c02, /* 1279 */
128'h8b85449cdf5ff0ef8522488cdb9ff0ef, /* 1280 */
128'h0107e683654100043883603cee079be3, /* 1281 */
128'h051300ff0e3743114701478145816390, /* 1282 */
128'h00371f1b00064803ec0689e36e89f005, /* 1283 */
128'h16fd060527810107e7b301e8183b0705, /* 1284 */
128'h67330187971b0187d81bf2e500670363, /* 1285 */
128'h67330087d79b01c878330087981b0107, /* 1286 */
128'h83751782170200be873b8fd98fe90107, /* 1287 */
128'h5697b765470147812585e31c97469381, /* 1288 */
128'h85930000659714900613c4a686930000, /* 1289 */
128'hbd8540e030efeae5051300006517e9e5, /* 1290 */
128'h9d633bfd20000c378bd2bd6100c4e493, /* 1291 */
128'h051300006517c2e5859300005597000b, /* 1292 */
128'h0189096300043903b711702000efe9e5, /* 1293 */
128'h34833ce030ef855a85d60f20061386e6, /* 1294 */
128'h37031404806324818cfd4981485c0709, /* 1295 */
128'h0793c7817c1c00f76f630c8937830209, /* 1296 */
128'h85224581b71ff0ef85224581cc5cf920, /* 1297 */
128'h852201442903c39d0044f793b29ff0ef, /* 1298 */
128'hd45ff0ef85ca290100896913ff397913, /* 1299 */
128'hf79368a000efe3e505130000651785ca, /* 1300 */
128'h6913ff397913852201442903c39d0084, /* 1301 */
128'h0000651785cad1bff0ef85ca29010049, /* 1302 */
128'h3983cfb50014f793660000efe3c50513, /* 1303 */
128'h86930000569701898c63038439030004, /* 1304 */
128'h7c1c31e030ef855a85d609c00613b966, /* 1305 */
128'h0037f693470d02043c2300492783cba9, /* 1306 */
128'h480d468100c907930189871308e69f63, /* 1307 */
128'h8763c3900086161bff87051363104591, /* 1308 */
128'h872a2685c3988f518361ff8737030106, /* 1309 */
128'h0027e793485ccbb5603cfeb690e30791, /* 1310 */
128'h6004cc9d49858889c85c9bf9485cc85c, /* 1311 */
128'hb30686930000569701848c6304043903, /* 1312 */
128'h040430232a0030ef855a85d60ca00613, /* 1313 */
128'hf0ef8522ef8d8b850089278300090963, /* 1314 */
128'hf0ef8522484cc85c9bf54985485cb4bf, /* 1315 */
128'h8b85bd85645020ef4505d8098ce3c43f, /* 1316 */
128'hf0ef8522b77100f926230009b783dbd9, /* 1317 */
128'h010964830009398397a667a1bf41b1bf, /* 1318 */
128'he43e002c4621854e639c00878913dcd5, /* 1319 */
128'h41635535b7dd87ca14e109a13c2020ef, /* 1320 */
128'hf406e84aec26f02204800513717908b0, /* 1321 */
128'hc41d5551842a192030ef892e84b2e44e, /* 1322 */
128'h89aa7b3010efa9e505130000551785a2, /* 1323 */
128'h508000efd0c5051300006517862285aa, /* 1324 */
128'h740270a2557d1ac030ef852200099d63, /* 1325 */
128'he01c200007b78082614569a2694264e2, /* 1326 */
128'hc45c4789c7890024f793f40401242423, /* 1327 */
128'hb7f9c45c4785d8f145018885bfe94501, /* 1328 */
128'h050ef73ff06f20000537458146098082, /* 1329 */
128'h1141711c80822501638897aa200007b7, /* 1330 */
128'h569702f40263200007b7e4066380e022, /* 1331 */
128'h85930000659734c00613a3a686930000, /* 1332 */
128'h703c15e030efbfe5051300006517bee5, /* 1333 */
128'h110180820141640260a2557de3914505, /* 1334 */
128'h85a2501010efe42eec064501842ae822, /* 1335 */
128'h71797a00006f6105468560e266226442, /* 1336 */
128'he052e44ee84aec26f022f40620000513, /* 1337 */
128'h30efc62505130000651784aa098030ef, /* 1338 */
128'h4bf010ef4501479010ef0001b5031a00, /* 1339 */
128'hc485051300006517681c224010ef842a, /* 1340 */
128'h05130000651706f44583402000ef638c, /* 1341 */
128'hc505051300006517546c3f2000efc465, /* 1342 */
128'h458358303dc000ef91c115c20085d59b, /* 1343 */
128'h569b0086571bc46505130000651706c4, /* 1344 */
128'h561b0ff6f6930ff777130ff677930106, /* 1345 */
128'hc3850513000065175c0c3b2000ef0186, /* 1346 */
128'hc789bc25859300006597545c3a4000ef, /* 1347 */
128'hc285051300006517bb05859300006597, /* 1348 */
128'h0f2030efc345051300006517384000ef, /* 1349 */
128'h2783d8dfb0ef1ce58593000065977448, /* 1350 */
128'h6617e789b8c6061300006617584c19c4, /* 1351 */
128'h00efc125051300006517eea606130000, /* 1352 */
128'h00006a174401ed9ff0ef852645813460, /* 1353 */
128'h20000913c149899300006997c14a0a13, /* 1354 */
128'h318000ef8552e7810004059b01f47793, /* 1355 */
128'h00f5f6130405854e0007c583008487b3, /* 1356 */
128'h051300006517fd241de3302000ef8191, /* 1357 */
128'h69a2694264e2740270a22f2000ef1565, /* 1358 */
128'h0083b7830103b7038082614545016a02, /* 1359 */
128'hfe6393811782278540f707b30003b683, /* 1360 */
128'hb78300a7002300f3b8230017079300d7, /* 1361 */
128'hb7038082450180820007802345050103, /* 1362 */
128'hb7038f999201020596130103b7830083, /* 1363 */
128'hfff7059b00c6f5638e9dfff706930003, /* 1364 */
128'h00b6e6630103b7030007869b47819d9d, /* 1365 */
128'h00d3b823001706938082852e00070023, /* 1366 */
128'hbfd900d7002307850006c68300f506b3, /* 1367 */
128'h0693430540a0053be681000556634301, /* 1368 */
128'h86ba4e250ff6f81304100693c2190610, /* 1369 */
128'h6a630ff5761302b8f53b0005089b3859, /* 1370 */
128'hfec68fa306850ff676130306061b04ae, /* 1371 */
128'h059340e0063b8536fcb8ffe302b8d53b, /* 1372 */
128'h07930003076302f6e96300a606bb0300, /* 1373 */
128'h559b9d1900050023050500f5002302d0, /* 1374 */
128'h00b7ea630006879bfff5081b46810015, /* 1375 */
128'hb7d1feb50fa30505bf4500c8063b8082, /* 1376 */
128'hc30300d7063397ba9381178240f807bb, /* 1377 */
128'h01178023006600230685000648830007, /* 1378 */
128'heccef4a6f8a2597d011cf0ca7119b7e1, /* 1379 */
128'hf42afc3e843684b2e0dafc86e4d6e8d2, /* 1380 */
128'h03000a9306c00a1302500993f82af02e, /* 1381 */
128'hc52d8f1d0004c50377a2774202095913, /* 1382 */
128'h086304d7ff639381178276820017079b, /* 1383 */
128'hc503bfe1e71ff0ef0201039304850135, /* 1384 */
128'hc783035510634781048905450f630014, /* 1385 */
128'hf36346a50ff7f793fd07879bcb9d0004, /* 1386 */
128'h0f630640069304890014c503478100f6, /* 1387 */
128'h079304d50f630580069302a6eb6306d5, /* 1388 */
128'h790674a6744670e6f55d08f509630630, /* 1389 */
128'h808261090007051b6b066aa66a4669e6, /* 1390 */
128'h06e50e6307300713b74d048d0024c503, /* 1391 */
128'h00840b13f6e51ee30700071300a76c63, /* 1392 */
128'h02e5006307500713a00d460146850038, /* 1393 */
128'h00840b13fa850613f6e510e307800713, /* 1394 */
128'hf8b50693a81145c10016361346850038, /* 1395 */
128'h400845a946010016b693003800840b13, /* 1396 */
128'hf0ef0028020103930005059be31ff0ef, /* 1397 */
128'h00840b130201039300044503a809dd1f, /* 1398 */
128'h7433600000840b13b5fd845ad89ff0ef, /* 1399 */
128'h020103930005059b501010ef85220124, /* 1400 */
128'hfc3ef83aec061034f436715db7f18522, /* 1401 */
128'h8082616160e2e8dff0efe436e4c6e0c2, /* 1402 */
128'hec06100005931014862ef436f032715d, /* 1403 */
128'h60e2e69ff0efe436e4c6e0c2fc3ef83a, /* 1404 */
128'h1234862afe36fa32f62e710d80826161, /* 1405 */
128'heac2e6bee2baea22ee06080810000593, /* 1406 */
128'h125020ef0808842ae3fff0efe436eec6, /* 1407 */
128'hb303679c691c80826135645260f28522, /* 1408 */
128'hec63479d808245018302000303630087, /* 1409 */
128'h97360025971358e686930000469704b7, /* 1410 */
128'h795c878297b6e426e822ec061101431c, /* 1411 */
128'h0e7010ef908114827540f55c08c52483, /* 1412 */
128'h610545016442e90064a260e202945433, /* 1413 */
128'h058e05e135f1bfe1617cbff17d5c8082, /* 1414 */
128'h11418082557d8082557db7f1659c95aa, /* 1415 */
128'h681c00055e63ff5ff0ef842ae406e022, /* 1416 */
128'h60a264028522000307630207b303679c, /* 1417 */
128'h557d80820141640260a2450183020141, /* 1418 */
128'h879300004797150200a7eb6347ad8082, /* 1419 */
128'h05130000651780826108953e81755267, /* 1420 */
128'h715d83020007b303679c691c80828065, /* 1421 */
128'h078517824785d23e47d502f1102347a1, /* 1422 */
128'hd402e486100c200007930030e83ee42e, /* 1423 */
128'h07374d148082616160a6fd3ff0efcc3e, /* 1424 */
128'h041322813823dc01011308e6e0634004, /* 1425 */
128'h348322113c232291342385a2980101f1, /* 1426 */
128'h0a0447830a04c703e909fadff0ef1a05, /* 1427 */
128'h2301340323813083fb60051300f70d63, /* 1428 */
128'h47830dd4c70380822401011322813483, /* 1429 */
128'h1be30c0447830c04c703fef711e30dd4, /* 1430 */
128'h4611fcf715e30e0447830e04c703fcf7, /* 1431 */
128'h4501fd4559b010ef0d4485130d440593, /* 1432 */
128'h3e800513842af022717980824501bf65, /* 1433 */
128'h00011023858a460185226ea020eff406, /* 1434 */
128'h7d000513e509842af21ff0efc202c402, /* 1435 */
128'h717980826145740270a285226cc020ef, /* 1436 */
128'hc402c23ef406f022478500f110234785, /* 1437 */
128'h86934bdc008006b74538691cc195842a, /* 1438 */
128'h07378fd98f75600006b78ff58ff9f806, /* 1439 */
128'hec9ff0ef8522858a4601c43e8fd94000, /* 1440 */
128'h711d80826145740270a2c43c47b2e119, /* 1441 */
128'he0ca07c55783c23e47d500f1102347b5, /* 1442 */
128'h6a056989fdf949370107979bf852fc4e, /* 1443 */
128'hc43e842e8b2af456ec86f05ae4a6e8a2, /* 1444 */
128'h4601e00a0a13e0098993080909134495, /* 1445 */
128'h1005f79345b2ed15e71ff0ef855a858a, /* 1446 */
128'hc7950125f7b3054795630135f7b3c789, /* 1447 */
128'hfba00513d4dff0ef6605051300005517, /* 1448 */
128'h7b027aa27a4279e2690664a6644660e6, /* 1449 */
128'h5863fff40a9bfe04c5e334fd80826125, /* 1450 */
128'h8456b74d84565d6020ef3e8005130080, /* 1451 */
128'hf0ef6325051300005517fc8047e34501, /* 1452 */
128'h7139e7a919c52783bf6df9200513d07f, /* 1453 */
128'hf822858a460147d5c42e00f1102347c1, /* 1454 */
128'h2783c11ddddff0efc23e842af426fc06, /* 1455 */
128'hf0ef8522858a46014495cb918b891b84, /* 1456 */
128'h612174a2744270e2f8ed34fdc901dc7f, /* 1457 */
128'he0cae4a6711d80824501bfd545018082, /* 1458 */
128'h47c906d7f66384b6892a4785e8a2ec86, /* 1459 */
128'hcf3108c92783260102f1102302c92703, /* 1460 */
128'h854a100c47850030cc3ee42e4755d432, /* 1461 */
128'h4785e529842ad6fff0efc83eca26d23a, /* 1462 */
128'h100c47f5460102f1102347b10497f063, /* 1463 */
128'h00005517c11dd4fff0efd23ed402854a, /* 1464 */
128'h64a6644660e68522c41ff0ef58c50513, /* 1465 */
128'hb74d02f6063bbf6147c5808261256906, /* 1466 */
128'hf822fc067139b7c54401b7d50004841b, /* 1467 */
128'h4148842ace05e456e852ec4ef04af426, /* 1468 */
128'h4583c11d892a4a4010ef8ab684b28a2e, /* 1469 */
128'h85b3681000054d63891fa0ef852200b4, /* 1470 */
128'hf0ef542505130000551700b67a630144, /* 1471 */
128'hecdff0ef854a08c92583a0894481bd7f, /* 1472 */
128'h0089f3630207e4030109378389a6f96d, /* 1473 */
128'h1ae3f01ff0ef854a85d6865286a2844e, /* 1474 */
128'h028784339a22408989b308c96783fc85, /* 1475 */
128'h74a279028526744270e2fc0999e39aa2, /* 1476 */
128'h161b0086969b808261216aa26a4269e2, /* 1477 */
128'h00f11023030006b78e55479971390106, /* 1478 */
128'hc432c23e84aafc06f426f82247f58e55, /* 1479 */
128'h0593e919c4dff0ef8526858a4601440d, /* 1480 */
128'h612174a2744270e2d8bff0ef85263e80, /* 1481 */
128'h07b7db0101134d18bfcdfc79347d8082, /* 1482 */
128'h24813023241134239fb923213823bffc, /* 1483 */
128'hf36349013ffc07372331342322913c23, /* 1484 */
128'hc03ff0ef84aa85a2980101f104131ce7, /* 1485 */
128'h20000513e7991a04b7831e051a63892a, /* 1486 */
128'h1e0505631a04b5031aa4b023748020ef, /* 1487 */
128'h47210c04478313d010ef85a220000613, /* 1488 */
128'h97ba078a0cc70713000047171cf76d63, /* 1489 */
128'h00e7fd63cc981ff78793400407b753b8, /* 1490 */
128'h0147d69307a68007071367050d442783, /* 1491 */
128'h8f2309b449830a044783f8dc00d77363, /* 1492 */
128'hc7890e244783e7810019f9938b8506f4, /* 1493 */
128'h0a04478300098a6308f480a30b344783, /* 1494 */
128'h0e24478306f48fa309c44783c7898b89, /* 1495 */
128'h0a844783fcdc07c60c84861309140713, /* 1496 */
128'h4583fff74783e0fc07c6468109d40513, /* 1497 */
128'hffe745839fad0105959b0087979b0007, /* 1498 */
128'h85b30e04458300098c634685c39197ae, /* 1499 */
128'h070de21c07ce02b787b30dd4478302f5, /* 1500 */
128'h470308e4478304098f63fce514e30621, /* 1501 */
128'h47039fb90087171b0107979b468508d4, /* 1502 */
128'h0dd4478302f707330e04470397ba08c4, /* 1503 */
128'h08a4470308b44783f8fc07ce02e787b3, /* 1504 */
128'h171b089447039fb90107171b0187979b, /* 1505 */
128'hc319f4fc54d89fb9088447039fb90087, /* 1506 */
128'h09c44783c7898b850a044783f4fc07a6, /* 1507 */
128'h852645850af006134685c6b5e3918bfd, /* 1508 */
128'h0e0447830af407a34785e141e0bff0ef, /* 1509 */
128'h00098663c79954dc08f4aa2300a7979b, /* 1510 */
128'h0dd447030e044783f8dc07a60d442783, /* 1511 */
128'h0a74478308f4ac2300a7979b02e787bb, /* 1512 */
128'h3483854a240134032481308308f48023, /* 1513 */
128'h80822501011322813983230139032381, /* 1514 */
128'hd79b00a7d71b50fcf3dd8b850af44783, /* 1515 */
128'haa2302f707bb278527058bfd8b7d0057, /* 1516 */
128'h5a6020efdd4d1a04b503892ab75d08f4, /* 1517 */
128'h0113b7655929b7755951bf451a04b023, /* 1518 */
128'h3023229134232281382322113c23dc01, /* 1519 */
128'h54a9468104b7ec6306f5846347892321, /* 1520 */
128'hd3fff0ef892a45850b900613842eed85, /* 1521 */
128'h0413ed91258199f5ffe4059be11d84aa, /* 1522 */
128'h4783e9159a7ff0ef854a85a2980101f1, /* 1523 */
128'h2301340323813083df400493e3990b94, /* 1524 */
128'h80822401011322813483220139038526, /* 1525 */
128'hb7554685fef760e354a94705ffc5879b, /* 1526 */
128'hf022f406e44ee84aec267179bfd984aa, /* 1527 */
128'h892e9be10079f6930ff5f99308154783, /* 1528 */
128'hc519cc1ff0ef84aa45850b3006138edd, /* 1529 */
128'h852685ca00091c6300f51e63842a57b5, /* 1530 */
128'h013505a317a010ef8526842a86dff0ef, /* 1531 */
128'h8082614569a2694264e2740270a28522, /* 1532 */
128'h289134232881382328113c23d6010113, /* 1533 */
128'h275134232741382327313c2329213023, /* 1534 */
128'h259134232581382325713c2327613023, /* 1535 */
128'h4d180ac7ed63478923b13c2325a13023, /* 1536 */
128'h87933ffc07b79f3dbff7879bbffc07b7, /* 1537 */
128'h14050513000055178a2e8b3284aabfe7, /* 1538 */
128'h5517e7b90016f79307e4c68300e7eb63, /* 1539 */
128'h8522f8400413f8eff0ef162505130000, /* 1540 */
128'h28013903288134832901340329813083, /* 1541 */
128'h26013b0326813a8327013a0327813983, /* 1542 */
128'h24013d0324813c8325013c0325813b83, /* 1543 */
128'h55170984a70380822a01011323813d83, /* 1544 */
128'h02f109930045aa83db4513a505130000, /* 1545 */
128'hac83e79102eaf7bb060a8063fe09f993, /* 1546 */
128'h1385051300005517cb8902ecf7bb0005, /* 1547 */
128'h4b8502eadabb54dcb7615429f14ff0ef, /* 1548 */
128'h8956866200ca05138c0a009c9c9be399, /* 1549 */
128'h78bb0017859b0005280343114e054781, /* 1550 */
128'hf0ef132505130000551700088d6302e8, /* 1551 */
128'h02e858bbb7f14b814a814c81b7c9ed6f, /* 1552 */
128'h0107c78397d2078e0208006301162023, /* 1553 */
128'h0ffbfb9300fbebb300be17bbcb898b85, /* 1554 */
128'h8963fa6596e387ae061105210128893b, /* 1555 */
128'hee068de311450513000055178a89000b, /* 1556 */
128'hc603ee051ae3842af8aff0ef852685ce, /* 1557 */
128'h9e3d0087979b0106161b09e9c78309f9, /* 1558 */
128'h0000551785ca01267a63963e09d9c783, /* 1559 */
128'hc683008a4783b5c9e50ff0ef10c50513, /* 1560 */
128'h0fe6f9138b89c71989360017f7130a79, /* 1561 */
128'h0017861b4591450547810016e913c399, /* 1562 */
128'h17bbc39d8b850017579b4b9897d2078e, /* 1563 */
128'h8b050189191b0187979b0027571b00c5, /* 1564 */
128'h79130127e933c70d4189591b4187d79b, /* 1565 */
128'h0a69c78302d90263fcb614e387b20ff9, /* 1566 */
128'h352020ef0c45051300005517ef898b85, /* 1567 */
128'h09b9c783bfd100f97933fff7c793b5a9, /* 1568 */
128'hdb8ff0ef0f45051300005517cb898b85, /* 1569 */
128'he3958b850af9c783e20b05e3b535547d, /* 1570 */
128'he579a21ff0ef852645850af006134685, /* 1571 */
128'haa2300a7979b0e09c7830af987a34785, /* 1572 */
128'h061b00dcd6bb003d169b4d914d0108f4, /* 1573 */
128'hf0ef852645850ff676130ff6f693f88d, /* 1574 */
128'h169b4c8dfdbd1fe32d05e9458a2a9edf, /* 1575 */
128'h76130ff6f693f8ca061b00dad6bb003a, /* 1576 */
128'h10e32a05e92d9c5ff0ef852645850ff6, /* 1577 */
128'h4c818ad209b00d934d6108f00a13ff9a, /* 1578 */
128'h0ff6f6930196d6bb45858656000c2683, /* 1579 */
128'h0ffafa932ca12a85e139999ff0ef8526, /* 1580 */
128'hfdba18e30c110ffa7a132a0dffac90e3, /* 1581 */
128'hed19971ff0ef8526458509c0061386de, /* 1582 */
128'h468501279b630a79c783d4fb0ee34785, /* 1583 */
128'hb381842a953ff0ef8526458509b00613, /* 1584 */
128'h842a941ff0ef852645850a70061386ca, /* 1585 */
128'h842ae406e0221141b325842ab335dd79, /* 1586 */
128'h0187b303679c681c00055e63ffdfe0ef, /* 1587 */
128'h45058302014160a26402852200030763, /* 1588 */
128'hf822fc06f426713980820141640260a2, /* 1589 */
128'h92635529478500f5866384aa4791f04a, /* 1590 */
128'h842e07c4d78300f110230370079304f5, /* 1591 */
128'hc43ec24a8526858a46010107979b4955, /* 1592 */
128'h4791c24a00f110234799ed19d44ff0ef, /* 1593 */
128'hf0ef8526858a4601c43e478900f41f63, /* 1594 */
128'h478580826121790274a2744270e2d26f, /* 1595 */
128'h869b4f5c6918e215b7cdc402fef414e3, /* 1596 */
128'h069b0007859b4f1887ae00d5f3630007, /* 1597 */
128'h0823dd0c0007859b87ba00d5f3630007, /* 1598 */
128'h10000737691c80828082c18ff06f02c5, /* 1599 */
128'heccef0caf4a6fc86f8a2070d4b9c7119, /* 1600 */
128'hc17c8fd9f466f862fc5ee0dae4d6e8d2, /* 1601 */
128'heb8d6b9c679c681cc509f07ff0ef842a, /* 1602 */
128'hb98ff0efef4505130000551702042423, /* 1603 */
128'h69e674a679068526744670e6f8500493, /* 1604 */
128'h808261097ca27c427be26b066aa66a46, /* 1605 */
128'h1af42c23478df93ff0eff3e54481541c, /* 1606 */
128'hb8eff0ef852202042c2302f408234785, /* 1607 */
128'h6b9c679c8522681c409010ef7d000513, /* 1608 */
128'h282318042e2308842783f94584aa9782, /* 1609 */
128'hb5eff0ef8522d85c478508f422231a04, /* 1610 */
128'hcdaff0ef8522f13ff0ef852245814601, /* 1611 */
128'h47a1000505a346d000ef8522f14984aa, /* 1612 */
128'h07138ff94bdc00ff8737681c00f11023, /* 1613 */
128'h8522858a460147d50aa00713e3991aa0, /* 1614 */
128'h079300c14703e911be0ff0efc23ec43a, /* 1615 */
128'h3e900913cc1c800207b700f715630aa0, /* 1616 */
128'h00ff8bb74b0502900a934a5503700993, /* 1617 */
128'h10238522858a460140000cb780020c37, /* 1618 */
128'h4c18681ce13db9eff0efc402c2520131, /* 1619 */
128'h1563c43e0177f7b3c25a4bdc01511023, /* 1620 */
128'hf0ef8522858a4601c43e0197e7b30187, /* 1621 */
128'h06090863397d0007ca6347b2ed1db76f, /* 1622 */
128'h800207374c14bf45319010ef3e800513, /* 1623 */
128'h41e7d79bc43ccc188001073700e68563, /* 1624 */
128'hb55d18f40ca3478506041e23d45c8b85, /* 1625 */
128'h4581becff0ef852202f51f63f9200793, /* 1626 */
128'h47850007d663443ced09c1cff0ef8522, /* 1627 */
128'hd965c04ff0ef85224585bfd118f40c23, /* 1628 */
128'hfa1004939fcff0efd705051300005517, /* 1629 */
128'hef26f706f3227161551cb58584aab595, /* 1630 */
128'heee6f2e2f6defadafed6e352e74eeb4a, /* 1631 */
128'h1e7010ef45018baae3b54401e6eeeaea, /* 1632 */
128'he7b5180b8ca3198bc783c7b1199bc783, /* 1633 */
128'hc2be855e008c479d460104f110234789, /* 1634 */
128'h1b8ba78312050ae3842aaa2ff0efc482, /* 1635 */
128'ha88ff0ef855e008c46014495cf818b85, /* 1636 */
128'ha031020ba423f4fd34fd10050de3842a, /* 1637 */
128'h741a70ba8522d55d842ad99ff0ef855e, /* 1638 */
128'h7c167bb67b567af66a1a69ba695a64fa, /* 1639 */
128'h8c23048ba7838082615d6db66d566cf6, /* 1640 */
128'h10ef4501afeff0ef855e0407c163180b, /* 1641 */
128'h855e45853e8009139081020514931550, /* 1642 */
128'h0007cc63048ba783f155842ab1eff0ef, /* 1643 */
128'h10ef0640051308a96fe3131010ef8526, /* 1644 */
128'h048ba78300fbac23400007b7bfe91bf0, /* 1645 */
128'h06fb9e23478502fba6238b8541e7d79b, /* 1646 */
128'h40010737a0292007071b40010737bf05, /* 1647 */
128'h3a178a1d0036571b00ebac234007071b, /* 1648 */
128'h260396529752060a8b3d6d2a0a130000, /* 1649 */
128'h02c7073b018ba88345050f8747031086, /* 1650 */
128'ha823180bae231a0ba8238a0500c7d61b, /* 1651 */
128'h8b3d0107d71b08eba22308eba42304cb, /* 1652 */
128'h090ba8231408dd63090ba62300e5183b, /* 1653 */
128'h003f07370107979b14070f6302cba703, /* 1654 */
128'h97b32689078546a18fd90106d79b8f7d, /* 1655 */
128'hb4230c0bb0230a0bbc23030787b300d7, /* 1656 */
128'hb8230e0bb0230c0bbc230c0bb8230c0b, /* 1657 */
128'ha70308fba6230107d463200007930afb, /* 1658 */
128'hc21508fba82300e7f46320000793090b, /* 1659 */
128'h0107979b471100e78e63577d04cba783, /* 1660 */
128'hf0efc282c4be04e11023855e008c4601, /* 1661 */
128'h4601495507cbd78304f11023479d8f6f, /* 1662 */
128'h8d8ff0efc4bec2ca855e008c0107979b, /* 1663 */
128'h80a357fd08fbaa234785e4051ce3842a, /* 1664 */
128'h855ee40510e3842ac94ff0ef855e08fb, /* 1665 */
128'h842aff3fe0ef855e00b54583113000ef, /* 1666 */
128'h100007b754075963018ba703e20515e3, /* 1667 */
128'hd78306f110230370079304fba0232789, /* 1668 */
128'hd4bed2ca855e0107979b108c460107cb, /* 1669 */
128'h07930bf104934905d2caed05874ff0ef, /* 1670 */
128'h4991d48206f11023988102091a930330, /* 1671 */
128'hd05aec56e826855e108c08104b210a85, /* 1672 */
128'hbb75842afe0996e339fdc529844ff0ef, /* 1673 */
128'h40040737bda940030737bd8940020737, /* 1674 */
128'h08bba82300b515bb89bd0165d59bbd91, /* 1675 */
128'h01e6d71b8ff90027979b17716705b545, /* 1676 */
128'h4098bd798a9d938100f6d69b17828fd9, /* 1677 */
128'h0087161b0187179b0187569b00ff0537, /* 1678 */
128'hf00706138fd167410087569b8e698fd5, /* 1679 */
128'h0187559b40d804fbaa2327818fd58ef1, /* 1680 */
128'h0087571b8de90087159b8ecd0187169b, /* 1681 */
128'h8b3d0187d71b04ebac238f558f718ecd, /* 1682 */
128'h8001073708d70e634689c70109270d63, /* 1683 */
128'h040ba7830007596302d7971300ebac23, /* 1684 */
128'h07b7018ba70304fba0238fd920000737, /* 1685 */
128'h639c12a787930000579708f713638001, /* 1686 */
128'h3497044ba783f0be0ff10c13040ba903, /* 1687 */
128'h478500f97933fe0c7c934ea484930000, /* 1688 */
128'h97bb478540980a8583f9791302079a93, /* 1689 */
128'h0000379704a1ebc5278100f977b300e7, /* 1690 */
128'h9b85051300005517fef493e34cc78793, /* 1691 */
128'h071b80011737b949df400413e15fe0ef, /* 1692 */
128'h800207370007456303079713b7bda007, /* 1693 */
128'h0ab70ff104934905bfa980030737b785, /* 1694 */
128'h886339fd09053ac54995988119020100, /* 1695 */
128'h07931030c33e47d508f1102347990209, /* 1696 */
128'he0efdc3ef84af426c556855e010c0400, /* 1697 */
128'h44dcfbe18b8583a54cdce6051de3eb7f, /* 1698 */
128'h8ff90087d79b0087969bf00707136741, /* 1699 */
128'he793040ba783f20750e302e797138fd5, /* 1700 */
128'h06010993017d8b37bf0104fba0230087, /* 1701 */
128'hf7b300f977b30009ad0340dc840b0b1b, /* 1702 */
128'h0d6345a1400007b712078e63278101a7, /* 1703 */
128'h100005b700fd08634591200007b700fd, /* 1704 */
128'h8daa8bfff0ef855e0015b59340bd05b3, /* 1705 */
128'h073700ed0d6347a1400007370e051963, /* 1706 */
128'h40fd0d33100007b700ed086347912000, /* 1707 */
128'h409cd41fe0ef855e02fbaa23001d3793, /* 1708 */
128'h47994d850ae79d63470d00e786634705, /* 1709 */
128'h17c12d81810007b7d33e47d50af11023, /* 1710 */
128'h855e110c040007930110d53e00fde7b3, /* 1711 */
128'h010cc783e541dcffe0efc93ee556e166, /* 1712 */
128'ha583efd91afba823409c09b790638bbd, /* 1713 */
128'h18fbae2308bba2230017b79317ed088b, /* 1714 */
128'h0af1102303700793895ff0ef855e4601, /* 1715 */
128'h855e110c0107979b4601475507cbd783, /* 1716 */
128'h47b56702ed05d7ffe0efd53ee03ad33a, /* 1717 */
128'h4791d5028dead33a0af11023fe0c7d13, /* 1718 */
128'he556e16ae43e855e110c011004000713, /* 1719 */
128'h37fd670267a2c521d51fe0efe03ac93a, /* 1720 */
128'h096ba2231afba823017d85b74785f3f5, /* 1721 */
128'h81dff0ef855e840585934601180bae23, /* 1722 */
128'h62e34581472db575def98be310bc0991, /* 1723 */
128'hbf91118725839752837902079713f6f7, /* 1724 */
128'h2783f006869300ff0537040d059366c1, /* 1725 */
128'h961b8f510187971b0187d61b0d11000d, /* 1726 */
128'h2e238fd98ff58f510087d79b8e690087, /* 1727 */
128'h00c7579b46a5008da703fda59ee3fefd, /* 1728 */
128'h1c63800306b7018ba60300f6f8638bbd, /* 1729 */
128'ha78397b6078a1be686930000369704d6, /* 1730 */
128'h67c100cda68308fbae230087171b1487, /* 1731 */
128'hd71bc78d27818fd18ff90186d61b17fd, /* 1732 */
128'h02e6073b3e800613c30503f777130126, /* 1733 */
128'ha02302d606bb02f757bb8a8d0106d69b, /* 1734 */
128'ha7831afbaa231b0ba7830adba2230afb, /* 1735 */
128'h08fba82308fba62320000793c79919cb, /* 1736 */
128'ha70300050623000515234a0000ef855e, /* 1737 */
128'h8693aaa78793ccccd6b7aaaab7b708cb, /* 1738 */
128'h37b3068600d036b327818ef98ff9ccc6, /* 1739 */
128'h36b38ef90f068693f0f0f6b79fb500f0, /* 1740 */
128'h8ef9f0068693ff0106b79fb5068a00d0, /* 1741 */
128'h8f750207161376c19fb5068e00d036b3, /* 1742 */
128'h92010a8bb783d11c9fb9071200e03733, /* 1743 */
128'hc603074bd68307abd70302c7d7b3ed10, /* 1744 */
128'h02450513694585930000459784aa06fb, /* 1745 */
128'h077bc883070ba683a8dfe0effef53623, /* 1746 */
128'h0ff6f8130106d71b0086d79b06cbc603, /* 1747 */
128'h000045970186d69b0ff777130ff7f793, /* 1748 */
128'h074ba603a59fe0ef04d4851367458593, /* 1749 */
128'h0106569b062485136705859300004597, /* 1750 */
128'h10ef8526a39fe0ef8a3d8abd0146561b, /* 1751 */
128'h2785100007b7b0cd02fba42347857c20, /* 1752 */
128'h00f778631a0bb603400407b704fba023, /* 1753 */
128'h4517e611b5f1e225ecf769e3400407b7, /* 1754 */
128'h0016879b700006b7b1295e2505130000, /* 1755 */
128'h1abba42303f7f5930c46478304fba023, /* 1756 */
128'h0216869bc58900c7f593cd910027f593, /* 1757 */
128'h04dba0230106e693040ba68304dba023, /* 1758 */
128'h04fba02300c7e793040ba783d7dd8b85, /* 1759 */
128'h044ba783040ba983e6f769e3400407b7, /* 1760 */
128'hf0ef2981855e00f9f9b34601088ba583, /* 1761 */
128'h00003b174a850564849300003497daaf, /* 1762 */
128'h409c09ec8c9300003c974c2d06cb0b13, /* 1763 */
128'h98e304a1eb99278100f9f7b300fa97bb, /* 1764 */
128'hbd2197bfe0ef51e5051300004517ff64, /* 1765 */
128'h10000db720000d370389091300003917, /* 1766 */
128'h04f719630017b79317ed00494703409c, /* 1767 */
128'hc3a127818ff900f9f7b30009270340dc, /* 1768 */
128'h855e0fb6f69345850b70061300894683, /* 1769 */
128'h855e45850b7006134681c90ddbbfe0ef, /* 1770 */
128'h180bae231a0ba823088ba783dabfe0ef, /* 1771 */
128'h0931941fe0ef855e035baa2308fba223, /* 1772 */
128'h4721400006b700092783bfa5fb9910e3, /* 1773 */
128'hb71341b787b301a78663471100d78963, /* 1774 */
128'h855e408c913fe0ef855e02ebaa230017, /* 1775 */
128'he79d0046f79300892683f14dfeffe0ef, /* 1776 */
128'hb79317ed088ba583ef8d1afba823409c, /* 1777 */
128'hf0ef855e460118fbae2308bba2230017, /* 1778 */
128'h0ff6f693bb35f53d9d9fe0ef855ec9af, /* 1779 */
128'hbfa1d171d13fe0ef855e45850b700613, /* 1780 */
128'h25839752837902079713fcfc65e34581, /* 1781 */
128'h00ec4641ef2ff06ffa100413bf6d1187, /* 1782 */
128'hd78304f11023478d6ce000ef06cb8513, /* 1783 */
128'h47d5855ec4be0107979b008c460107cb, /* 1784 */
128'h018ba783ec051163842a943fe0efc2be, /* 1785 */
128'h102347a506fb9e2304e157830007d663, /* 1786 */
128'h979b008c460107cbd783c2be479d04f1, /* 1787 */
128'he8051763842a90ffe0efc4be855e0107, /* 1788 */
128'h04cbae23018ba50345e646d647c64636, /* 1789 */
128'h4000073706bba42306dba22306fba023, /* 1790 */
128'h0007081b377d8b3d01a6571bf0e51c63, /* 1791 */
128'hdc850513000035171702ef056863450d, /* 1792 */
128'h80824501c56c8702972a4318972a8379, /* 1793 */
128'h5797808218b50d238082557d8082557d, /* 1794 */
128'he02247851141ef9d439cd86787930000, /* 1795 */
128'h12a000efd6f7282300005717842ae406, /* 1796 */
128'hfc5ff0ef852200055563ac0fe0ef8522, /* 1797 */
128'h640260a20dc000ef13e000ef02c00513, /* 1798 */
128'h07130000571780824501808201414501, /* 1799 */
128'h451785aa114102e790636394631cd3e7, /* 1800 */
128'h478160a2f3cfe0efe406452505130000, /* 1801 */
128'h87b600a604630fc7a60380820141853e, /* 1802 */
128'hf0efe42eec06110141488082853ebfd1, /* 1803 */
128'h470302b7006365a210354703c105fbdf, /* 1804 */
128'he06f610560e200f70c630ff007930815, /* 1805 */
128'h0513bfe545018082610560e25535e97f, /* 1806 */
128'hf0ef84aee822ec06e4261101bfcdf840, /* 1807 */
128'h0f840413e501ce0ff0ef842acd09f7df, /* 1808 */
128'hbfd555358082610564a2644260e2e080, /* 1809 */
128'hc3980015071b4388ae07879300005797, /* 1810 */
128'hac8787930000579780820f8505138082, /* 1811 */
128'he822c727879300005797110180824388, /* 1812 */
128'h644260e20094176384beec06e4266380, /* 1813 */
128'hf0ef8522c78119a447838082610564a2, /* 1814 */
128'he39cc427879300005797b7d56000a8cf, /* 1815 */
128'h5797e5088082a607af2300005797e79c, /* 1816 */
128'he308e518e11ce7886798c2a787930000, /* 1817 */
128'he8a2c124849300005497e4a6711d8082, /* 1818 */
128'he466e862ec5ef05af456f852fc4e6080, /* 1819 */
128'h338a0a1300004a1789aae0caec86e06a, /* 1820 */
128'h338b0b1300004b17338a8a9300004a97, /* 1821 */
128'h00004c9700050c1b338b8b9300004b97, /* 1822 */
128'h64a660e66446029415634d298bcc8c93, /* 1823 */
128'h6ca26c426be27b027aa27a4279e26906, /* 1824 */
128'hdb8fe06f612541e50513000045176d02, /* 1825 */
128'h89560007c36389524c1cc7914901541c, /* 1826 */
128'h0663d9afe0ef638c855a0fc42603681c, /* 1827 */
128'h00978e63601cd8efe0ef855e85ca0009, /* 1828 */
128'h0000451701a98863d80fe0ef856685e2, /* 1829 */
128'he8221101b77160002ea010ef84450513, /* 1830 */
128'hcfad44014d1cc1414401e04ae426ec06, /* 1831 */
128'hc7ad639cc7bd651ccbad511ccbbd4d5c, /* 1832 */
128'h842a1c0010ef45051c00059384aa892e, /* 1833 */
128'h02a347850ef52c234799c57c57fdcd21, /* 1834 */
128'he65ff0ef0405282303253023e90410f5, /* 1835 */
128'h0000179716f43c238fa78793fffff797, /* 1836 */
128'h26e787930000179718f4302327e78793, /* 1837 */
128'h0247c78385220ea42e23681c18f43423, /* 1838 */
128'h64a2644260e28522e99ff0ef10f40023, /* 1839 */
128'h86930000469717c0106f808261056902, /* 1840 */
128'h0017671302d786b365186294611c78e6, /* 1841 */
128'h553b93ed836d8f3d0127d713e1189736, /* 1842 */
128'h808225018d5d00f717bb40f007bb00f7, /* 1843 */
128'he4061141fc3ff06fa885051300005517, /* 1844 */
128'h0105151bfe9ff0ef842afefff0efe022, /* 1845 */
128'he4061141808201412501640260a28d41, /* 1846 */
128'hfd1ff0ef14020005041bfdbff0efe022, /* 1847 */
128'h87aa80820141640260a28d4115029001, /* 1848 */
128'h8082fb75fee78fa30785fff5c7030585, /* 1849 */
128'h06b30007470300f5873300c78c634781, /* 1850 */
128'hc70387aa8082f76d00e68023078500f5, /* 1851 */
128'h0785fff5c7030585eb09001786930007, /* 1852 */
128'he21987aab7d587b68082fb75fee78fa3, /* 1853 */
128'h963efb7d001786930007c70387b68082, /* 1854 */
128'h99e3d375fee78fa30785fff5c7030585, /* 1855 */
128'hc783000547030585808200078023fec7, /* 1856 */
128'he3994187d79b0187979b40f707bbfff5, /* 1857 */
128'h478100e6146347018082853ef37d0505, /* 1858 */
128'hc78300e587b30007c68300e507b3a015, /* 1859 */
128'he3994187d79b0187979b40f687bb0007, /* 1860 */
128'h000547830ff5f5938082853efee10705, /* 1861 */
128'h80824501bfcd0505c399808200b79363, /* 1862 */
128'hdffd808200b79363000547830ff5f593, /* 1863 */
128'h40a78533e7010007c70387aabfcd0505, /* 1864 */
128'hec06842ae42ee8221101bfcd07858082, /* 1865 */
128'h000547830ff5f593952265a2fe5ff0ef, /* 1866 */
128'h644260e24501fe857be3157d00b78663, /* 1867 */
128'h0007c70300b7856387aa95aa80826105, /* 1868 */
128'h07334781b7fd0785808240a78533e701, /* 1869 */
128'hfed60ee38082853eea990007468300f5, /* 1870 */
128'hbfd5872eb7d50785fa7d000746030705, /* 1871 */
128'ha021872eca890007468300f507334781, /* 1872 */
128'h8082853efa7d00074603070500d60863, /* 1873 */
128'h8fe380824501eb1900054703b7c50785, /* 1874 */
128'h87aeb7e50505fafd0007c6830785fee6, /* 1875 */
128'he519842a84aeec06e426e8221101bfd5, /* 1876 */
128'h85a68522cc1163808887879300005797, /* 1877 */
128'h00005797ef8100044783942afa1ff0ef, /* 1878 */
128'h610564a2644260e2852244018607b623, /* 1879 */
128'h00054783c519f9fff0ef852285a68082, /* 1880 */
128'h84a7b02300005797050500050023c781, /* 1881 */
128'h842ac891e822ec066104e4261101bfd9, /* 1882 */
128'he008050500050023c501f73ff0ef8526, /* 1883 */
128'h4783c11d8082610564a28526644260e2, /* 1884 */
128'h0017c703ce810007c68387aacf990005, /* 1885 */
128'hb7e5078900d780a300e780238082e311, /* 1886 */
128'hf69347a1eb0587aa0075771380824501, /* 1887 */
128'h00c508b387aaffed8f5537fd07220ff5, /* 1888 */
128'h5761003657930106ee6340f88833469d, /* 1889 */
128'h00c79763963e963a97aa078e02e78733, /* 1890 */
128'hfeb78fa30785bfe9fee7bc2307a18082, /* 1891 */
128'heb9d872a8b9d00b567b304b50463b7f5, /* 1892 */
128'h06b30006b80300f586b3a811471d4781, /* 1893 */
128'hfed765e340f606b30106b02307a100f5, /* 1894 */
128'h963a95be078e02e78733576100365793, /* 1895 */
128'h00f586b3808200f61363478100f50733, /* 1896 */
128'hb7e501068023078500f706b30006c803, /* 1897 */
128'he84af406e432ec26852e842af0227179, /* 1898 */
128'h6582892ace1184aa6622dd3ff0efe02e, /* 1899 */
128'hf0ef944a864a8522fff6091300c56463, /* 1900 */
128'h64e269428526740270a200040023f75f, /* 1901 */
128'h00a5e963842ae406e022114180826145, /* 1902 */
128'h883280820141640260a28522f53ff0ef, /* 1903 */
128'h0733fef605e317fd4781fff6461386ae, /* 1904 */
128'h00b7002397220005c58300e685b300f8, /* 1905 */
128'h00e507b3a821478100e614634701b7e5, /* 1906 */
128'h9f9507050006c6830007c78300e586b3, /* 1907 */
128'h4783808200c51363962a8082853ed3f5, /* 1908 */
128'h842af0227179bfc50505feb78de30005, /* 1909 */
128'hd19ff0ef892ee44ef406e84aec26852e, /* 1910 */
128'h008509bbd0dff0ef8522c8990005049b, /* 1911 */
128'h740270a2852244010097db63408987bb, /* 1912 */
128'h852285ca86268082614569a2694264e2, /* 1913 */
128'h0ff5f593962abfe10405d17df83ff0ef, /* 1914 */
128'h00150793000547038082450100c51463, /* 1915 */
128'hef630ff5f59347c1b7ed853efeb70be3, /* 1916 */
128'hc7038082853e4781e60187aa260100c7, /* 1917 */
128'h00757793b7f5367d0785feb71ce30007, /* 1918 */
128'h0007c68387aa00a7083b9f1d4721c39d, /* 1919 */
128'h1702fed819e30007869b0785fcb69de3, /* 1920 */
128'h179300b7e733008597938e19953a9301, /* 1921 */
128'h27018edd00365713020796938fd90107, /* 1922 */
128'hf8b71fe30007c703d24d8a1deb1187aa, /* 1923 */
128'h0a63008785130007b803bfcd367d0785, /* 1924 */
128'hfef51be30785f8b712e30007c70300d8, /* 1925 */
128'h00054703e7c9419cb7f1377d87aabfa5, /* 1926 */
128'h000027970015470306f71e6303000793, /* 1927 */
128'hc6898a850006c68300e786b318478793, /* 1928 */
128'h04d71763078006930ff777130207071b, /* 1929 */
128'hcf950447f7930007c78397ba00254703, /* 1930 */
128'h02f71f630300079300054703c19c47c1, /* 1931 */
128'h4703973e13c707130000271700154783, /* 1932 */
128'h07130ff7f7930207879bc7098b050007, /* 1933 */
128'h8082c19c47a1a809050900e79c630780, /* 1934 */
128'he82211018082fae78fe34741bfed47a9, /* 1935 */
128'h00c16583f61ff0efc632ec06006c842e, /* 1936 */
128'h079b000547030ee80813000028174681, /* 1937 */
128'h9863044678930006460300f806330007, /* 1938 */
128'h7893808261058536644260e2ec050008, /* 1939 */
128'h86b3feb7f4e3fd07879b00088b630046, /* 1940 */
128'hfe07079bc6098a09b7d196be050502d5, /* 1941 */
128'h7139b7e1e008b7cdfc97879b0ff7f793, /* 1942 */
128'h842ae42e00063023f04afc06f426f822, /* 1943 */
128'h744270e25529e90165a2b03ff0ef84b2, /* 1944 */
128'h8522082c892a862e80826121790274a2, /* 1945 */
128'hcb010007c703fe8782e367e2f5dff0ef, /* 1946 */
128'he088fcf718e347a9fd279be307858f81, /* 1947 */
128'h00e6846302d0071300054683b7e94501, /* 1948 */
128'h60a2f23ff0efe40605051141f2dff06f, /* 1949 */
128'h842ee406e02211418082014140a00533, /* 1950 */
128'h04630007c70304b00693601cf0dff0ef, /* 1951 */
128'h60a202d70e630470069300e6ea6302d7, /* 1952 */
128'h069302d7076304d00693808201416402, /* 1953 */
128'h052a069007130017c683fed716e306b0, /* 1954 */
128'h00e69863042007130027c683fce69fe3, /* 1955 */
128'hbfd50789bff1052a052ab7e9e01c078d, /* 1956 */
128'he0dff0efc632ec06006c842ee8221101, /* 1957 */
128'h4703f9a8081300002817468100c16583, /* 1958 */
128'h78930006460300f806330007079b0005, /* 1959 */
128'h61058536644260e2ec05000898630446, /* 1960 */
128'hf4e3fd07879b00088b63004678938082, /* 1961 */
128'hc6098a09b7d196be050502d586b3feb7, /* 1962 */
128'he008b7cdfc97879b0ff7f793fe07079b, /* 1963 */
128'h601cf87ff0ef842ee406e0221141b7e1, /* 1964 */
128'h00e6ea6302d704630007c70304b00693, /* 1965 */
128'h80820141640260a202d70e6304700693, /* 1966 */
128'hfed716e306b0069302d7076304d00693, /* 1967 */
128'hc683fce69fe3052a069007130017c683, /* 1968 */
128'hb7e9e01c078d00e69863042007130027, /* 1969 */
128'he406e0221141bfd50789bff1052a052a, /* 1970 */
128'hfff5c70300a405b3951ff0efe589842a, /* 1971 */
128'h4703973efff58513ec07879300002797, /* 1972 */
128'h80820141557d640260a2e7198b110007, /* 1973 */
128'h00074703973e00054703fea47ae3157d, /* 1974 */
128'h014105054581462960a26402f77d8b11, /* 1975 */
128'h05220085579bfa5ff06f4581d7dff06f, /* 1976 */
128'h46a54781808201419141154211418d5d, /* 1977 */
128'h059b27018082853ee319000547034629, /* 1978 */
128'hfd07879b9fb902f607bb00b6e763fd07, /* 1979 */
128'h00a04563842ee406e0221141b7c50505, /* 1980 */
128'hf0ef357d02b455bb45a900b7f86347a5, /* 1981 */
128'h0513014160a2640202a4753b4529fe7f, /* 1982 */
128'h3b230000471707fe47854e80006f0305, /* 1983 */
128'he822110180823ef73b23000047173ef7, /* 1984 */
128'h85aa84ae862ee4263e84041300004417, /* 1985 */
128'he00c95a660e2600ca1fff0efec066008, /* 1986 */
128'h00004797e42611018082610564a26442, /* 1987 */
128'he04ae8223ac48493000044973bc78793, /* 1988 */
128'hec068d250513000045170004b9036380, /* 1989 */
128'hc0ef85a26088b6ffd0ef85a24124043b, /* 1990 */
128'h8c85051300004517862286aa608ce41f, /* 1991 */
128'hf14025730ff0000f0000100fb55fd0ef, /* 1992 */
128'h8593000025976902834a64a260e26442, /* 1993 */
128'h8432e406e02211418302610525013265, /* 1994 */
128'h640260a28522547d00850363830fa0ef, /* 1995 */
128'h01258413f22271698082450180820141, /* 1996 */
128'hf0ef892eea4aee26f606852289aae64e, /* 1997 */
128'h0505f9aff0ef852600a404b30505fa6f, /* 1998 */
128'hee631ff00793fff5071beabff0ef9526, /* 1999 */
128'hf78ff0ef85222ea7a3230000479704e7, /* 2000 */
128'h9526f6aff0ef656505130000351784aa, /* 2001 */
128'h842af5aff0ef852204a7f2630ff00793, /* 2002 */
128'h00a405b3f4cff0ef6385051300003517, /* 2003 */
128'h741270b2a8dfd0ef8185051300004517, /* 2004 */
128'h4717200007938082615569b2695264f2, /* 2005 */
128'h850a458110000613b75528f725230000, /* 2006 */
128'hf0ef850a5f45859300003597885ff0ef, /* 2007 */
128'h359700f7096302f0079301294703e10f, /* 2008 */
128'h850a85a2e24ff0ef850a7ea585930000, /* 2009 */
128'h858a43902447879300004797e1cff0ef, /* 2010 */
128'h17934405a1dfd0ef7d05051300003517, /* 2011 */
128'h0000471722f7362300004717451101f4, /* 2012 */
128'h00a7942300004797db7ff0ef22f73623, /* 2013 */
128'h4611fea79e2300004797da9ff0ef4501, /* 2014 */
128'h4797eafff0ef854eff05859300004597, /* 2015 */
128'he426ec06e8221101b7991e8797230000, /* 2016 */
128'h84ae450d892a08c7df638432478de04a, /* 2017 */
128'h451708a7956325010004d783d6bff0ef, /* 2018 */
128'h25010024d783d55ff0ef1be555030000, /* 2019 */
128'hdc1ff0ef00448513ffc4059b06a79a63, /* 2020 */
128'h4517f8a7952300004797d39ff0ef4511, /* 2021 */
128'h000047974611d25ff0ef18e555030000, /* 2022 */
128'hf0ef854af6c5859300004597f6a79b23, /* 2023 */
128'h1645d58300004597256000ef4535e2bf, /* 2024 */
128'h4797240000ef02000513d33ff0ef4515, /* 2025 */
128'h0000471727850007d78314e787930000, /* 2026 */
128'h278d439c134787930000479714f71023, /* 2027 */
128'h909fd0ef6dc50513000035170087cf63, /* 2028 */
128'h60e2d5fff06f6105690264a260e26442, /* 2029 */
128'hf022f406717980826105690264a26442, /* 2030 */
128'h0f230115c70300e10fa346890105c703, /* 2031 */
128'h02f70a63478d00d70e6301e1570300e1, /* 2032 */
128'hd06f61456bc505130000351770a27402, /* 2033 */
128'hd0efe42e6945051300003517842a8b7f, /* 2034 */
128'hd8dff06f614570a265a2740285228a7f, /* 2035 */
128'h0113ebfff06f614505c170a241907402, /* 2036 */
128'h842a232130232291342322813823dc01, /* 2037 */
128'h22113c230028218006134581893284ae, /* 2038 */
128'he802c44a08282040061385a6e84ff0ef, /* 2039 */
128'h23813083f63ff0ef8522002cec2ff0ef, /* 2040 */
128'h24010113220139032281348323013403, /* 2041 */
128'h45974611cb8104a7d783000047978082, /* 2042 */
128'he40611418082cf3ff06fe32585930000, /* 2043 */
128'ha70300e57763878e1041e7034ec000ef, /* 2044 */
128'h1007e78310a7a22310e1a02327051001, /* 2045 */
128'h4501808201418d5d91011782150260a2, /* 2046 */
128'hfc1ff0ef84aae426e822ec0611018082, /* 2047 */
128'h150202f407b33e800793428000ef842a, /* 2048 */
128'h610564a28d0502a7d533644260e29101, /* 2049 */
128'h00ef842af95ff0efe022e40611418082, /* 2050 */
128'h60a202f407b324078793000f47b73fc0, /* 2051 */
128'h1101808202a7d5330141910115026402, /* 2052 */
128'h892af63ff0ef84aae04ae426e822ec06, /* 2053 */
128'h24040413000f443702a485333ca000ef, /* 2054 */
128'hfe856ee3f45ff0ef0405944a02855433, /* 2055 */
128'he426110180826105690264a2644260e2, /* 2056 */
128'h68048493842ae04aec06e822009894b7, /* 2057 */
128'hf0ef41240433854a89260084f3638922, /* 2058 */
128'h80826105690264a2644260e2f47dfa1f, /* 2059 */
128'h100007b7808200054503808200b50023, /* 2060 */
128'h4783100007378082020575130147c503, /* 2061 */
128'h07b7808200a70023dfe50207f7930147, /* 2062 */
128'h476d00e78623f8000713000782231000, /* 2063 */
128'h071300e78623470d0007822300e78023, /* 2064 */
128'h808200e788230200071300e78423fc70, /* 2065 */
128'h60a2e50900044503842ae406e0221141, /* 2066 */
128'h2797b7f50405fa5ff0ef808201416402, /* 2067 */
128'h97aa973e811100f57713e2a787930000, /* 2068 */
128'h00f5802300e580a30007c78300074703, /* 2069 */
128'hf0efec068121842a002ce82211018082, /* 2070 */
128'hf0ef00914503f65ff0ef00814503fd1f, /* 2071 */
128'h00814503fb7ff0ef0ff47513002cf5df, /* 2072 */
128'h644260e2f43ff0ef00914503f4bff0ef, /* 2073 */
128'h892af406e84aec26f022717980826105, /* 2074 */
128'hf0ef0ff57513002c0089553b54e14461, /* 2075 */
128'h00914503f13ff0ef346100814503f81f, /* 2076 */
128'h694264e2740270a2fe9410e3f0bff0ef, /* 2077 */
128'h892af406e84aec26f022717980826145, /* 2078 */
128'h0ff57513002c0089553354e103800413, /* 2079 */
128'h4503ed1ff0ef346100814503f3fff0ef, /* 2080 */
128'h64e2740270a2fe9410e3ec9ff0ef0091, /* 2081 */
128'hf13ff0efec06002c1101808261456942, /* 2082 */
128'he9fff0ef00914503ea7ff0ef00814503, /* 2083 */
128'h439cff278793000047978082610560e2, /* 2084 */
128'h842e892aec4efc06f04af426f8227139, /* 2085 */
128'hb0efd9a505130000451702b7856384b2, /* 2086 */
128'h70e2fca7a32300004797c10d2501f3af, /* 2087 */
128'h471757fd8082612169e2790274a27442, /* 2088 */
128'h0000451785ca86260074faf725230000, /* 2089 */
128'h00004797c50d2501814fb0efd6450513, /* 2090 */
128'h0000351785a6049675634632f8a7a823, /* 2091 */
128'h2923000047174785d10fd0ef33450513, /* 2092 */
128'h099b00c4591be05ff0ef4521b775f6f7, /* 2093 */
128'h993e0039791332e78793000037970009, /* 2094 */
128'hbf5d2dc010ef854ede7ff0ef00094503, /* 2095 */
128'h0000100fbf95f287ab23000047979c25, /* 2096 */
128'h8593000025974305f14025730ff0000f, /* 2097 */
128'h859300003597460511418302037eca65, /* 2098 */
128'hd95fa0efe406f0e505130000451703e5, /* 2099 */
128'h014160a22d45051300003517c9092501, /* 2100 */
128'hc78fd0ef2e45051300003517c84fd06f, /* 2101 */
128'h0513000045172f658593000035974605, /* 2102 */
128'h051300003517c5112501db9fa0efc965, /* 2103 */
128'hc48fd0ef2fc5051300003517b7e92ee5, /* 2104 */
128'hea07a22300004797eb65051300000517, /* 2105 */
128'h000047978eaf90efe807ac2300004797, /* 2106 */
128'h059b60a2cb9927818fc9439ce9078793, /* 2107 */
128'hc08fd06f01412d650513000035170005, /* 2108 */
128'hc5112501bc6fb0efc305051300004517, /* 2109 */
128'h000035974605b7952d85051300003517, /* 2110 */
128'h3517c5112501cdbfa0ef4501f7c58593, /* 2111 */
128'hac05051300003517b7992d2505130000, /* 2112 */
128'h1141900200000023ef9ff0efbc4fd0ef, /* 2113 */
128'h0513000f4537a001d81ff0efe4062501, /* 2114 */
128'hdf870713000047178082450180822405, /* 2115 */
128'he30895360017869300756513157d631c, /* 2116 */
128'h110102b506338082953e055e10d00513, /* 2117 */
128'hc509842afd1ff0efe4328532ec06e822, /* 2118 */
128'h6105644260e28522980ff0ef45816622, /* 2119 */
128'he4062625051300003517114180828082, /* 2120 */
128'h450160a2ef7fc0ef20000537b44fd0ef, /* 2121 */
128'hb0002573808245018082450180820141, /* 2122 */
128'h862e86b287361141808202f5553347a9, /* 2123 */
128'hb08fd0efe40624e505130000351785aa, /* 2124 */
128'h952e842ae0221141a001cd3ff0ef4505, /* 2125 */
128'h640260a29522408007b3f57ff0efe406, /* 2126 */
128'h45058082450580824505808201418d7d, /* 2127 */
128'h00c684bb842ef406ec26f02271798082, /* 2128 */
128'h80826145450164e2740270a200961863, /* 2129 */
128'h200404136622e49fc0efe432852285b2, /* 2130 */
128'h808245098082450980824509bff92605, /* 2131 */
128'hf06f8082450180824501808280828082, /* 2132 */
128'h003796934781e426e822ec061101bd3f, /* 2133 */
128'h644260e200c7986300d5043300d584b3, /* 2134 */
128'h036360980004380380826105450164a2, /* 2135 */
128'hd0ef1c250513000035176090600c02e8, /* 2136 */
128'hd0ef1da505130000351785a28626a46f, /* 2137 */
128'h351784aafc26715dbf5d0785a001a36f, /* 2138 */
128'hec56f052f44ef84ae0a21da505130000, /* 2139 */
128'h3997a0afd0ef4401892ee45ee486e85a, /* 2140 */
128'h3b171d2a8a9300003a971ca989930000, /* 2141 */
128'h0b9b9eafd0ef854e4a411dab0b130000, /* 2142 */
128'h1863470187a69defd0ef855685de0004, /* 2143 */
128'h9c8fd0ef855a85de9d0fd0ef854e0327, /* 2144 */
128'h3517fd4417e3040503259963458187a6, /* 2145 */
128'h06b3a0a945019aefd0ef202505130000, /* 2146 */
128'h6394e390fff7c613c299863e8a850087, /* 2147 */
128'h86be8b05639000858733bf6d07a10705, /* 2148 */
128'h00003517058e02d60b63fff7c693c319, /* 2149 */
128'h1985051300003517970fd0ef16c50513, /* 2150 */
128'h79a2794274e2640660a6557d964fd0ef, /* 2151 */
128'h07a10585808261616ba26b426ae27a02, /* 2152 */
128'h020005138aaa6a05fc56e0d27159b751, /* 2153 */
128'he8caf0a2f486f062f45ef85ae4ceeca6, /* 2154 */
128'hb6bff0ef44818bb28b2ee46ee86aec66, /* 2155 */
128'h9793542c0c1300003c179c4a0a134981, /* 2156 */
128'h351703749b6300fb0cb300fa8db30034, /* 2157 */
128'h694670a674068eefd0ef16a505130000, /* 2158 */
128'h86266da26d426ce27c027ba26a0669a6, /* 2159 */
128'he47ff06f61657ae285567b4264e685da, /* 2160 */
128'hc25fe0ef8d2ac2bfe0ef842ac31fe0ef, /* 2161 */
128'h1d1b0105151b0344f7b3c1ffe0ef892a, /* 2162 */
128'h91011402150201a4643300a96533010d, /* 2163 */
128'hf0ef4521ef8100adb02300acb0238d41, /* 2164 */
128'hf0ef0007c50397e20039f7930985ad9f, /* 2165 */
128'hf822fc06e032e42e7139b7ad0485ac9f, /* 2166 */
128'he0ef842abc9fe0ef89aaec4ef04af426, /* 2167 */
128'h151bbb7fe0ef84aabbdfe0ef892abc3f, /* 2168 */
128'h65a2660215028fc18d450109179b0105, /* 2169 */
128'h00e588330037971347818d5d91011782, /* 2170 */
128'h854e790274a270e2744200c79c63974e, /* 2171 */
128'h8ea907856314d8dff06f6121863e69e2, /* 2172 */
128'h7139b7f100e830238f2900083703e314, /* 2173 */
128'h89aaec4ef04af426f822fc06e032e42e, /* 2174 */
128'hb45fe0ef892ab4bfe0ef842ab51fe0ef, /* 2175 */
128'h8d450109179b0105151bb3ffe0ef84aa, /* 2176 */
128'h47818d5d9101178265a2660215028fc1, /* 2177 */
128'h744200c79c63974e00e5883300379713, /* 2178 */
128'hf06f6121863e69e2854e790274a270e2, /* 2179 */
128'h8f0900083703e3148e8907856314d15f, /* 2180 */
128'hf822fc06e032e42e7139b7f100e83023, /* 2181 */
128'he0ef842aad9fe0ef89aaec4ef04af426, /* 2182 */
128'h151bac7fe0ef84aaacdfe0ef892aad3f, /* 2183 */
128'h65a2660215028fc18d450109179b0105, /* 2184 */
128'h00e588330037971347818d5d91011782, /* 2185 */
128'h854e790274a270e2744200c79c63974e, /* 2186 */
128'h86b307856314c9dff06f6121863e69e2, /* 2187 */
128'h00e8302302a7073300083703e31402a6, /* 2188 */
128'hf04af426f822fc06e032e42e7139b7e1, /* 2189 */
128'h892aa57fe0ef842aa5dfe0ef89aaec4e, /* 2190 */
128'h179b0105151ba4bfe0ef84aaa51fe0ef, /* 2191 */
128'h9101178265a2660215028fc18d450109, /* 2192 */
128'h9c63974e00e588330037971347818d5d, /* 2193 */
128'h863e69e2854e790274a270e2744200c7, /* 2194 */
128'hd6b3078563144505e111c21ff06f6121, /* 2195 */
128'h00e8302302a7573300083703e31402a6, /* 2196 */
128'hf04af426f822fc06e032e42e7139b7d1, /* 2197 */
128'h892a9d7fe0ef842a9ddfe0ef89aaec4e, /* 2198 */
128'h179b0105151b9cbfe0ef84aa9d1fe0ef, /* 2199 */
128'h9101178265a2660215028fc18d450109, /* 2200 */
128'h9c63974e00e588330037971347818d5d, /* 2201 */
128'h863e69e2854e790274a270e2744200c7, /* 2202 */
128'h3703e3148ec907856314ba1ff06f6121, /* 2203 */
128'he032e42e7139b7f100e830238f490008, /* 2204 */
128'h965fe0ef89aaec4ef04af426f822fc06, /* 2205 */
128'he0ef84aa959fe0ef892a95ffe0ef842a, /* 2206 */
128'h15028fc18d450109179b0105151b953f, /* 2207 */
128'h0037971347818d5d9101178265a26602, /* 2208 */
128'h74a270e2744200c79c63974e00e58833, /* 2209 */
128'h6314b29ff06f6121863e69e2854e7902, /* 2210 */
128'h00e830238f6900083703e3148ee90785, /* 2211 */
128'hf04af426f822fc06e032e42e7139b7f1, /* 2212 */
128'h892a8e7fe0ef842a8edfe0ef89aaec4e, /* 2213 */
128'h179b0105151b8dbfe0ef84aa8e1fe0ef, /* 2214 */
128'h9081178265a2660214828fc18cc90109, /* 2215 */
128'h1c6396ae00d988330037169347018fc5, /* 2216 */
128'h863a69e2854e790274a270e2744200c7, /* 2217 */
128'h00a83023e28800f70533ab1ff06f6121, /* 2218 */
128'h051300003517892ae8ca7159bfc90705, /* 2219 */
128'hf062f45ef85afc56e0d2e4cef0a2cce5, /* 2220 */
128'hcf9fc0ef44018b3289aeec66eca6f486, /* 2221 */
128'hcc0b8b9300003b97cb8a0a1300003a17, /* 2222 */
128'hc0ef855204000a93cc8c0c1300003c17, /* 2223 */
128'hcc9fc0ef8885855e85a2fff44493cd7f, /* 2224 */
128'h00f905b30036179314fd460140900cb3, /* 2225 */
128'h85a2cabfc0efe43285520566186397ce, /* 2226 */
128'ha17ff0ef854a85ce6622ca3fc0ef8562, /* 2227 */
128'h051300003517fb541be32405e12984aa, /* 2228 */
128'h64e669468526740670a6c83fc0efcd65, /* 2229 */
128'h61656ce27c027ba27b427ae26a0669a6, /* 2230 */
128'he198e3988726c2918766001676938082, /* 2231 */
128'h351784aaeca67159bfc154fdbf590605, /* 2232 */
128'hfc56e0d2e4cee8caf0a2bfa505130000, /* 2233 */
128'h8ab2892ee86af486ec66f062f45ef85a, /* 2234 */
128'h3b17be29899300003997c23fc0ef4401, /* 2235 */
128'h3c17ee2b8b9300003b97ee2b0b130000, /* 2236 */
128'h0a13be2c8c9300003c97bdac0c130000, /* 2237 */
128'hbd03cba500147793bf1fc0ef854e0400, /* 2238 */
128'hfffd45134601bdffc0ef856285a2000b, /* 2239 */
128'h854e05561c6397ca00f485b300361793, /* 2240 */
128'h6622bbbfc0ef856685a2bc3fc0efe432, /* 2241 */
128'h1ae32405e5298d2a92fff0ef852685ca, /* 2242 */
128'h70a6b9bfc0efbee5051300003517fb44, /* 2243 */
128'h7b427ae26a0669a6694664e6856a7406, /* 2244 */
128'h000b3d03808261656d426ce27c027ba2, /* 2245 */
128'he198e398872ac291876a00167693bf49, /* 2246 */
128'h3517842ae8a2711db7e15d7db7790605, /* 2247 */
128'hf05af456f852e0cae4a6b0a505130000, /* 2248 */
128'hc0ef4c018ab284aefc4eec86e862ec5e, /* 2249 */
128'h0b1300003b17af69091300003917b37f, /* 2250 */
128'h854a10000a13b06b8b9300003b97afeb, /* 2251 */
128'hb09fc0ef855a85ce000c099bb15fc0ef, /* 2252 */
128'h17130187e7b38fd9008c1793010c1713, /* 2253 */
128'h8fd9028c17138fd9020c17138fd9018c, /* 2254 */
128'h171346018fd9038c17138fd9030c1713, /* 2255 */
128'he432854a05561763972600e406b30036, /* 2256 */
128'h85a66622abdfc0ef855e85ceac5fc0ef, /* 2257 */
128'hf94c19e30c05e91d89aa831ff0ef8522, /* 2258 */
128'h644660e6a9dfc0efaf05051300003517, /* 2259 */
128'h6be27b027aa27a4279e2690664a6854e, /* 2260 */
128'h59fdb74d0605e29ce31c808261256c42, /* 2261 */
128'ha20505130000351784aaf4a67119bff1, /* 2262 */
128'hf862fc5ee0dae4d6e8d2eccef0caf8a2, /* 2263 */
128'hc0ef44018b32892eec6efc86f06af466, /* 2264 */
128'h8c9300003c97a06a0a1300003a17a47f, /* 2265 */
128'h00003d1703f00c13498507f00b93a0ec, /* 2266 */
128'h85a2a1bfc0ef855208000a93a0cd0d13, /* 2267 */
128'h95b300e99733408b873ba13fc0ef8566, /* 2268 */
128'h1a6397ca00f486b30036179346010089, /* 2269 */
128'hc0ef856a85a29effc0efe43285520566, /* 2270 */
128'he1398daaf5aff0ef852685ca66229e7f, /* 2271 */
128'hc0efa1a5051300003517fb541be32405, /* 2272 */
128'h6a4669e6790674a6856e744670e69c7f, /* 2273 */
128'h61096de27d027ca27c427be26b066aa6, /* 2274 */
128'he398bf610605e28ce38c008c66638082, /* 2275 */
128'h351784aaf4a67119b7f15dfdbfe5e298, /* 2276 */
128'he4d6e8d2eccef0caf8a293a505130000, /* 2277 */
128'h892eec6efc86f06af466f862fc5ee0da, /* 2278 */
128'h920a0a1300003a17961fc0ef44018b32, /* 2279 */
128'h0c13498507f00b93928c8c9300003c97, /* 2280 */
128'h855208000a93926d0d1300003d1703f0, /* 2281 */
128'h408b87bb92dfc0ef856685a2935fc0ef, /* 2282 */
128'hfff6c693fff7c793008996b300f997b3, /* 2283 */
128'h05661a63974a00e485b3003617134601, /* 2284 */
128'h8f9fc0ef856a85a2901fc0efe4328552, /* 2285 */
128'h2405e1398daae6cff0ef852685ca6622, /* 2286 */
128'h8d9fc0ef92c5051300003517fb5417e3, /* 2287 */
128'h6aa66a4669e6790674a6856e744670e6, /* 2288 */
128'h808261096de27d027ca27c427be26b06, /* 2289 */
128'he19ce31cbf610605e194e314008c6663, /* 2290 */
128'h0000351784aaf4a67119b7f15dfdbfe5, /* 2291 */
128'he0dae4d6e8d2eccef0caf8a284c50513, /* 2292 */
128'h8a32892eec6efc86f06af466f862fc5e, /* 2293 */
128'h3c178329899300003997873fc0ef4401, /* 2294 */
128'h08100b134d0507f00a9383ac0c130000, /* 2295 */
128'hc0ef854e834c8c9300003c9703f00b93, /* 2296 */
128'h07bb408a873b83ffc0ef856285a2847f, /* 2297 */
128'h0024079b8f5d00ed173300fd17b3408b, /* 2298 */
128'hc893fff743138fd5008d16b300fd17b3, /* 2299 */
128'h1c6396ca00d48533003616934601fff7, /* 2300 */
128'hc0ef856685a2ffefc0efe432854e0546, /* 2301 */
128'hed298daad6aff0ef852685ca6622ff6f, /* 2302 */
128'h051300003517f8f41be3080007932405, /* 2303 */
128'h790674a6856e744670e6fd2fc0ef8265, /* 2304 */
128'h7d027ca27c427be26b066aa66a4669e6, /* 2305 */
128'h85be008bea6300167813808261096de2, /* 2306 */
128'h85bab7610605e10ce28c85c600080363, /* 2307 */
128'hf0ca7119bf755dfdbfc5859afe080be3, /* 2308 */
128'hfc5ee8d2ecce7365051300002517892a, /* 2309 */
128'he0dae4d6f4a6f8a2fc86ec6ef06af466, /* 2310 */
128'h00002a17f5cfc0ef4b81e03289aef862, /* 2311 */
128'h00002d17724c8c9300002c9771ca0a13, /* 2312 */
128'h003b949b01779c3347854da172cd0d13, /* 2313 */
128'h856685da00848b3bf30fc0ef85524401, /* 2314 */
128'h0036171367824601fffc4a93f24fc0ef, /* 2315 */
128'hc0efe432855206f61063974e00e90833, /* 2316 */
128'h854a85ce6622efefc0ef856a85daf06f, /* 2317 */
128'hfbb41be38c562405e9318b2ac72ff0ef, /* 2318 */
128'h051300002517fafb90e3040007932b85, /* 2319 */
128'h790674a6855a744670e6ed2fc0ef7265, /* 2320 */
128'h7d027ca27c427be26b066aa66a4669e6, /* 2321 */
128'h85d6e11185e200167513808261096de2, /* 2322 */
128'h7175b7e95b7db749060500b83023e30c, /* 2323 */
128'h69850200051384ae892af4cef8cafca6, /* 2324 */
128'he506f86afc66e0e2e4dee8daecd6f0d2, /* 2325 */
128'h4a098ba68beff0ef8acae032f46ee122, /* 2326 */
128'h9c4989934ca131ec0c1300003c174b01, /* 2327 */
128'h003d969367824d81a88d0d1300003d17, /* 2328 */
128'hbb6ff0ef854a85a6866e04fd966396d6, /* 2329 */
128'h251702fa18638aa68bca4785ed4d842a, /* 2330 */
128'h640a60aa8522e1efc0ef69a505130000, /* 2331 */
128'h6c066ba66b466ae67a0679a6794674e6, /* 2332 */
128'hec36b7754a05808261497da27d427ce2, /* 2333 */
128'h954fe0efe82a95afe0ef842a960fe0ef, /* 2334 */
128'h8d5d0105151b664267a294efe0efe42a, /* 2335 */
128'h8d4166e29101140215028c510106161b, /* 2336 */
128'h018786b34781e28828a7b02300003797, /* 2337 */
128'h00230ff6f693078500fb86330006c683, /* 2338 */
128'h4521ef910ba1033df7b3ff9795e300d6, /* 2339 */
128'h97ea8b8d00078b1b001b079bfe7fe0ef, /* 2340 */
128'hbfb1547dbf050d85fd3fe0ef0007c503, /* 2341 */
128'h0200051384ae892af4cef8cafca67175, /* 2342 */
128'hf86afc66e0e2e4dee8daecd6f0d26985, /* 2343 */
128'h8ba6f9dfe0ef8acae032f46ee122e506, /* 2344 */
128'h89934ca1204c0c1300003c174b014a09, /* 2345 */
128'h969367824d81966d0d1300003d179c49, /* 2346 */
128'hf0ef854a85a6866e04fd966396d6003d, /* 2347 */
128'h02fa18638aa68bca4785ed4d842aa94f, /* 2348 */
128'h60aa8522cfcfc0ef5785051300002517, /* 2349 */
128'h6ba66b466ae67a0679a6794674e6640a, /* 2350 */
128'hb7754a05808261497da27d427ce26c06, /* 2351 */
128'he0efe82a838fe0ef842a83efe0efec36, /* 2352 */
128'h0105151b664267a282cfe0efe42a832f, /* 2353 */
128'h66e29101140215028c510106161b8d5d, /* 2354 */
128'h86b34781e28816a7b323000037978d41, /* 2355 */
128'h92c116c2078900fb86330006d6830187, /* 2356 */
128'hef910ba1033df7b3ff9795e300d61023, /* 2357 */
128'h8b8d00078b1b001b079bec5fe0ef4521, /* 2358 */
128'h547dbf050d85eb1fe0ef0007c50397ea, /* 2359 */
128'hfff5861389b2ecce711980826505bfb1, /* 2360 */
128'h0000251785aa842a892e962af0caf8a2, /* 2361 */
128'hf862fc5ee0dae4d6e8d2f4a64b450513, /* 2362 */
128'h5793c1afc0efe436fc86ec6ef06af466, /* 2363 */
128'h4a8b0b1300002b1744854a81e03e0039, /* 2364 */
128'h4a8c0c1300002c174a8b8b9300002b97, /* 2365 */
128'h4b0d0d1300002d174a8c8c9300002c97, /* 2366 */
128'h080a0a1300003a174b0d8d9300002d97, /* 2367 */
128'hbc8fc0ef4a450513000025170299f863, /* 2368 */
128'h6aa66a4669e6790674a68556744670e6, /* 2369 */
128'h808261096de27d027ca27c427be26b06, /* 2370 */
128'h855e85ce00098663ba0fc0ef855a85a6, /* 2371 */
128'hc0ef856a85e6b8efc0ef8562b94fc0ef, /* 2372 */
128'hc0ef856ee129952ff0ef85226582b86f, /* 2373 */
128'h000a358302f74c636722010a2783b76f, /* 2374 */
128'h3783b5afc0ef4265051300002517c985, /* 2375 */
128'h9782852295a20049561300195593008a, /* 2376 */
128'hb7d14a89b3cfc0ef4105051300002517, /* 2377 */
128'hbf890485b2cfc0ef1905051300002517, /* 2378 */
128'hec26f022f4063fe50513000025177179, /* 2379 */
128'h0000251704000593c5dfe0efe44ee84a, /* 2380 */
128'h4185051300002517b00fc0ef3fc50513, /* 2381 */
128'hae8fc0ef43c5051300002517af4fc0ef, /* 2382 */
128'h4441adafc0ef44851405051300002517, /* 2383 */
128'h853346054685008495b3497901f49993, /* 2384 */
128'h740270a2ff2417e3e73ff0ef24050135, /* 2385 */
128'h131b460580828082614569a2694264e2, /* 2386 */
128'h87f245a901f61e1346814881470100c5, /* 2387 */
128'h97aa0007802397aa0007802340000813, /* 2388 */
128'h13e397aa387d0007802397aa00078023, /* 2389 */
128'h26f38e15c020267302b71d632705fe08, /* 2390 */
128'h059302a68733411686b33e800513c000, /* 2391 */
128'h473302a767b302b345bb02c747334000, /* 2392 */
128'h10e3a3afc06f3d6505130000251702a7, /* 2393 */
128'he4061141bf51c00028f3c02026f3fac7, /* 2394 */
128'hf0ef4509f75ff0ef4505f7bff0ef4501, /* 2395 */
128'h4541f63ff0ef4521f69ff0ef4511f6ff, /* 2396 */
128'he388400007b791011502bff1f5dff0ef, /* 2397 */
128'h400007b7808225016388400007b78082, /* 2398 */
128'h7b88400007b7808225016b880007b823, /* 2399 */
128'h8d510106161b8d5d0085979b80822501, /* 2400 */
128'h871b4000063747812581f788400007b7, /* 2401 */
128'h7a98400006b73e80079300b76f630007, /* 2402 */
128'h80827388400007b7ffe537fdc3198b09, /* 2403 */
128'hbfc1f618078500076703973600279713, /* 2404 */
128'h35fd00b7d763842a4785e406e0221141, /* 2405 */
128'h879300002797883dfedff0ef0045551b, /* 2406 */
128'he06f014160a2640200044503943e3467, /* 2407 */
128'h151b67050185579b9d3d00b007b7a5df, /* 2408 */
128'he8228fd9058565133007071311010085, /* 2409 */
128'hec06c43e454d458946010034842ec62a, /* 2410 */
128'hf49ff0ef454d460100344589f55ff0ef, /* 2411 */
128'h00d5802300f556b357610380079385a2, /* 2412 */
128'h80826105644260e2fee79ae3058537e1, /* 2413 */
128'hec86ec5ef05af456f852e0cae4a6711d, /* 2414 */
128'hff860a1b490184b28aae8b2afc4ee8a2, /* 2415 */
128'h008a853b012b09b30009041b40000bb7, /* 2416 */
128'h16024084863bf6dff0ef002c03446863, /* 2417 */
128'h64a6644660e6f1dfd0ef9201854e002c, /* 2418 */
128'h808261256be27b027aa27a4279e26906, /* 2419 */
128'hb0230921f3bff0ef00c4541b85ce2421, /* 2420 */
128'he486f2a5051300002517715dbf4d008b, /* 2421 */
128'he45ee85aec56f052f44ef84afc26e0a2, /* 2422 */
128'hd17f70eff6c5051300000517864fc0ef, /* 2423 */
128'h89930000199744014905e9b50005059b, /* 2424 */
128'h0ab7e9ab0b1300002b174bc1097e3169, /* 2425 */
128'hea5ff0ef0004051b45a101000a370010, /* 2426 */
128'hc50397ca009407b34481822fc0ef854e, /* 2427 */
128'h808fc0ef854ee8bff0ef048545890007, /* 2428 */
128'hfd4415e3ffdfb0ef9456855aff7494e3, /* 2429 */
128'h6b426ae27a0279a2794274e260a66406, /* 2430 */
128'h794274e260a66406b19fe06f61616ba2, /* 2431 */
128'h0513000025176ba26b426ae27a0279a2, /* 2432 */
128'h2505051300002517fc1fb06f6161e8e5, /* 2433 */
128'hec4ef04af426f822fc067139901fe06f, /* 2434 */
128'h0513000025178b9fe0efe05ae456e852, /* 2435 */
128'h00002917400009b744018dffe0ef18e5, /* 2436 */
128'h059b639097ce00341793449518c90913, /* 2437 */
128'h80effe9416e3f6ffb0ef0405854a0004, /* 2438 */
128'h400004b728cb0b1300002b174901d02f, /* 2439 */
128'h178a0a1300002a17168a8a9300002a97, /* 2440 */
128'he09c090585560007c783016907b34991, /* 2441 */
128'hb823f2bfb0ef8622240125816080608c, /* 2442 */
128'hfd391be3f1dfb0ef25818552688c0004, /* 2443 */
128'h071702f7646347190054579b0ff47413, /* 2444 */
128'h878297ba439c97ba078a6d2707130000, /* 2445 */
128'he0ef8522eedfb0ef1385051300002517, /* 2446 */
128'hed9fb0ef1345051300002517a001a39f, /* 2447 */
128'h1305051300002517b7f5e53ff0ef8522, /* 2448 */
128'h051300002517bfe9b9dff0efec5fb0ef, /* 2449 */
128'h00002517b7e1d30f80efeb3fb0ef12e5, /* 2450 */
128'h0000bf5dc75ff0efea1fb0ef12c50513, /* 2451 */
128'h00000000000000000000000000000000, /* 2452 */
128'h00000000000000000000000000000000, /* 2453 */
128'h00000000000000000000000000000000, /* 2454 */
128'h00000000000000000000000000000000, /* 2455 */
128'h00000000000000000000000000000000, /* 2456 */
128'h00000000000000000000000000000000, /* 2457 */
128'h00000000000000000000000000000000, /* 2458 */
128'h00000000000000000000000000000000, /* 2459 */
128'h00000000000000000000000000000000, /* 2460 */
128'h00000000000000000000000000000000, /* 2461 */
128'h00000000000000000000000000000000, /* 2462 */
128'h00000000000000000000000000000000, /* 2463 */
128'h08082828282828080808080808080808, /* 2464 */
128'h08080808080808080808080808080808, /* 2465 */
128'h101010101010101010101010101010a0, /* 2466 */
128'h10101010101004040404040404040404, /* 2467 */
128'h01010101010101010141414141414110, /* 2468 */
128'h10101010100101010101010101010101, /* 2469 */
128'h02020202020202020242424242424210, /* 2470 */
128'h08101010100202020202020202020202, /* 2471 */
128'h00000000000000000000000000000000, /* 2472 */
128'h00000000000000000000000000000000, /* 2473 */
128'h101010101010101010101010101010a0, /* 2474 */
128'h10101010101010101010101010101010, /* 2475 */
128'h01010101010101010101010101010101, /* 2476 */
128'h02010101010101011001010101010101, /* 2477 */
128'h02020202020202020202020202020202, /* 2478 */
128'h02020202020202021002020202020202, /* 2479 */
128'hc1bdceee242070dbe8c7b756d76aa478, /* 2480 */
128'hfd469501a83046134787c62af57c0faf, /* 2481 */
128'h895cd7beffff5bb18b44f7af698098d8, /* 2482 */
128'h49b40821a679438efd9871936b901122, /* 2483 */
128'he9b6c7aa265e5a51c040b340f61e2562, /* 2484 */
128'he7d3fbc8d8a1e68102441453d62f105d, /* 2485 */
128'h455a14edf4d50d87c33707d621e1cde6, /* 2486 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /* 2487 */
128'hfde5380c6d9d61228771f681fffa3942, /* 2488 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /* 2489 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /* 2490 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /* 2491 */
128'hfc93a039ab9423a7432aff97f4292244, /* 2492 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /* 2493 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /* 2494 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /* 2495 */
128'h0c07020d08030e09040f0a05000b0601, /* 2496 */
128'h020f0c090603000d0a0704010e0b0805, /* 2497 */
128'h09020b040d060f08010a030c050e0700, /* 2498 */
128'h6c5f7465735f64735f63736972776f6c, /* 2499 */
128'h6e67696c615f64730000000000006465, /* 2500 */
128'h645f6b6c635f64730000000000000000, /* 2501 */
128'h69747465735f64730000000000007669, /* 2502 */
128'h735f646d635f6473000000000000676e, /* 2503 */
128'h74657365725f64730000000074726174, /* 2504 */
128'h6e636b6c625f64730000000000000000, /* 2505 */
128'h69736b6c625f64730000000000000074, /* 2506 */
128'h6f656d69745f6473000000000000657a, /* 2507 */
128'h655f7172695f64730000000000007475, /* 2508 */
128'h5f63736972776f6c000000000000006e, /* 2509 */
128'h00000000646d635f74726174735f6473, /* 2510 */
128'h746e695f746961775f63736972776f6c, /* 2511 */
128'h000000000067616c665f747075727265, /* 2512 */
128'h00007172695f64735f63736972776f6c, /* 2513 */
128'h695f646d635f64735f63736972776f6c, /* 2514 */
128'h5f63736972776f6c0000000000007172, /* 2515 */
128'h007172695f646e655f617461645f6473, /* 2516 */
128'h00000000bffe9d8800000000bffeb0c0, /* 2517 */
128'h004c4b40004c4b400030000020000000, /* 2518 */
128'h6d6d5f6472616f62000000020000ffff, /* 2519 */
128'h00000000bffe4ecc0064637465675f63, /* 2520 */
128'h00000000bffe4d3a00000000bffe4adc, /* 2521 */
128'h00000000000000000000000000000000, /* 2522 */
128'hffffbab6ffffbab2ffffbab2ffffba8e, /* 2523 */
128'hffffbabaffffbabaffffbabaffffbaba, /* 2524 */
128'hffffcadcffffcad6ffffcad0ffffc92c, /* 2525 */
128'h00000000bffeb3e800000000bffeb3d8, /* 2526 */
128'h00000000bffeb41000000000bffeb3f8, /* 2527 */
128'h00000000bffeb44000000000bffeb428, /* 2528 */
128'h00000000bffeb47000000000bffeb458, /* 2529 */
128'h00000000bffeb4a000000000bffeb488, /* 2530 */
128'h00000000bffeb4d000000000bffeb4b8, /* 2531 */
128'h40040300400402004004010040040000, /* 2532 */
128'h40050000400405004004040140040400, /* 2533 */
128'h30000000000000030000000040050100, /* 2534 */
128'h60000000000000053000000000000001, /* 2535 */
128'h70000000000000027000000000000004, /* 2536 */
128'h00000001400000007000000000000000, /* 2537 */
128'h00000005000000012000000000000006, /* 2538 */
128'h20000000000000020000000040000000, /* 2539 */
128'h00000000100000000000000100000000, /* 2540 */
128'h1e19140f0d0c0a000000000000000000, /* 2541 */
128'h000186a00000271050463c37322d2823, /* 2542 */
128'h017d7840017d784000989680000f4240, /* 2543 */
128'h031975000319750002faf080018cba80, /* 2544 */
128'h02faf08005f5e10002faf080017d7840, /* 2545 */
128'h00000020000000000bebc2000c65d400, /* 2546 */
128'h00000200000001000000008000000040, /* 2547 */
128'h00002000000010000000080000000400, /* 2548 */
128'h0000c000000080000000600000004000, /* 2549 */
128'h37363534333231300002000000010000, /* 2550 */
128'h2043534952776f4c4645444342413938, /* 2551 */
128'h746f6f622d7520646573696d696e696d, /* 2552 */
128'h00000000647261432d445320726f6620, /* 2553 */
128'hfffff952fffff968fffff954fffff940, /* 2554 */
128'h00000000fffff98cfffff952fffff97a, /* 2555 */
128'he00600003800000039080000edfe0dd0, /* 2556 */
128'h00000000100000001100000028000000, /* 2557 */
128'h0000000000000000a806000059010000, /* 2558 */
128'h00000000010000000000000000000000, /* 2559 */
128'h02000000000000000400000003000000, /* 2560 */
128'h020000000f0000000400000003000000, /* 2561 */
128'h2c6874651b0000001400000003000000, /* 2562 */
128'h007665642d657261622d656e61697261, /* 2563 */
128'h2c687465260000001000000003000000, /* 2564 */
128'h0100000000657261622d656e61697261, /* 2565 */
128'h1a0000000300000000006e65736f6863, /* 2566 */
128'h303140747261752f636f732f2c000000, /* 2567 */
128'h0000003030323531313a303030303030, /* 2568 */
128'h00000000737570630100000002000000, /* 2569 */
128'h01000000000000000400000003000000, /* 2570 */
128'h000000000f0000000400000003000000, /* 2571 */
128'h40787d01380000000400000003000000, /* 2572 */
128'h03000000000000304075706301000000, /* 2573 */
128'h0300000080f0fa024b00000004000000, /* 2574 */
128'h03000000007570635b00000004000000, /* 2575 */
128'h03000000000000006700000004000000, /* 2576 */
128'h0000000079616b6f6b00000005000000, /* 2577 */
128'h7a6874651b0000001300000003000000, /* 2578 */
128'h0000766373697200656e61697261202c, /* 2579 */
128'h34367672720000000b00000003000000, /* 2580 */
128'h0b000000030000000000636466616d69, /* 2581 */
128'h0000393376732c76637369727c000000, /* 2582 */
128'h01000000850000000000000003000000, /* 2583 */
128'h6f72746e6f632d747075727265746e69, /* 2584 */
128'h04000000030000000000000072656c6c, /* 2585 */
128'h0000000003000000010000008f000000, /* 2586 */
128'h1b0000000f00000003000000a0000000, /* 2587 */
128'h000063746e692d7570632c7663736972, /* 2588 */
128'h01000000b50000000400000003000000, /* 2589 */
128'h01000000bb0000000400000003000000, /* 2590 */
128'h01000000020000000200000002000000, /* 2591 */
128'h0030303030303030384079726f6d656d, /* 2592 */
128'h6f6d656d5b0000000700000003000000, /* 2593 */
128'h67000000100000000300000000007972, /* 2594 */
128'h00000040000000000000008000000000, /* 2595 */
128'h0300000000636f730100000002000000, /* 2596 */
128'h03000000020000000000000004000000, /* 2597 */
128'h03000000020000000f00000004000000, /* 2598 */
128'h616972612c6874651b0000001f000000, /* 2599 */
128'h706d697300636f732d657261622d656e, /* 2600 */
128'h000000000300000000007375622d656c, /* 2601 */
128'h303240746e696c6301000000c3000000, /* 2602 */
128'h0d000000030000000000003030303030, /* 2603 */
128'h30746e696c632c76637369721b000000, /* 2604 */
128'hca000000100000000300000000000000, /* 2605 */
128'h07000000010000000300000001000000, /* 2606 */
128'h00000000670000001000000003000000, /* 2607 */
128'h0300000000000c000000000000000002, /* 2608 */
128'h006c6f72746e6f63de00000008000000, /* 2609 */
128'h7075727265746e690100000002000000, /* 2610 */
128'h3030634072656c6c6f72746e6f632d74, /* 2611 */
128'h04000000030000000000000030303030, /* 2612 */
128'h04000000030000000000000000000000, /* 2613 */
128'h0c00000003000000010000008f000000, /* 2614 */
128'h003063696c702c76637369721b000000, /* 2615 */
128'h03000000a00000000000000003000000, /* 2616 */
128'h0b00000001000000ca00000010000000, /* 2617 */
128'h10000000030000000900000001000000, /* 2618 */
128'h000000000000000c0000000067000000, /* 2619 */
128'he8000000040000000300000000000004, /* 2620 */
128'hfb000000040000000300000007000000, /* 2621 */
128'hb5000000040000000300000003000000, /* 2622 */
128'hbb000000040000000300000002000000, /* 2623 */
128'h75626564010000000200000002000000, /* 2624 */
128'h0000304072656c6c6f72746e6f632d67, /* 2625 */
128'h637369721b0000001000000003000000, /* 2626 */
128'h03000000003331302d67756265642c76, /* 2627 */
128'hffff000001000000ca00000008000000, /* 2628 */
128'h00000000670000001000000003000000, /* 2629 */
128'h03000000001000000000000000000000, /* 2630 */
128'h006c6f72746e6f63de00000008000000, /* 2631 */
128'h30303140747261750100000002000000, /* 2632 */
128'h08000000030000000000003030303030, /* 2633 */
128'h03000000003035373631736e1b000000, /* 2634 */
128'h00000010000000006700000010000000, /* 2635 */
128'h04000000030000000010000000000000, /* 2636 */
128'h040000000300000080f0fa024b000000, /* 2637 */
128'h040000000300000000c2010006010000, /* 2638 */
128'h04000000030000000200000014010000, /* 2639 */
128'h04000000030000000100000025010000, /* 2640 */
128'h04000000030000000200000030010000, /* 2641 */
128'h0100000002000000040000003a010000, /* 2642 */
128'h3030303240636d6d2d63736972776f6c, /* 2643 */
128'h10000000030000000000000030303030, /* 2644 */
128'h00000000000000200000000067000000, /* 2645 */
128'h14010000040000000300000000000100, /* 2646 */
128'h25010000040000000300000002000000, /* 2647 */
128'h1b0000000c0000000300000002000000, /* 2648 */
128'h0200000000636d6d2d63736972776f6c, /* 2649 */
128'h406874652d63736972776f6c01000000, /* 2650 */
128'h03000000000000003030303030303033, /* 2651 */
128'h2d63736972776f6c1b0000000c000000, /* 2652 */
128'h5b000000080000000300000000687465, /* 2653 */
128'h0400000003000000006b726f7774656e, /* 2654 */
128'h04000000030000000200000014010000, /* 2655 */
128'h06000000030000000300000025010000, /* 2656 */
128'h0300000000007fe3023e180047010000, /* 2657 */
128'h00000030000000006700000010000000, /* 2658 */
128'h01000000020000000080000000000000, /* 2659 */
128'h303440646e7277682d63736972776f6c, /* 2660 */
128'h0e000000030000000000303030303030, /* 2661 */
128'h6e7277682d63736972776f6c1b000000, /* 2662 */
128'h67000000100000000300000000000064, /* 2663 */
128'h00100000000000000000004000000000, /* 2664 */
128'h09000000020000000200000002000000, /* 2665 */
128'h2300736c6c65632d7373657264646123, /* 2666 */
128'h61706d6f6300736c6c65632d657a6973, /* 2667 */
128'h6f647473006c65646f6d00656c626974, /* 2668 */
128'h65736162656d697400687461702d7475, /* 2669 */
128'h6b636f6c630079636e6575716572662d, /* 2670 */
128'h63697665640079636e6575716572662d, /* 2671 */
128'h75746174730067657200657079745f65, /* 2672 */
128'h2d756d6d006173692c76637369720073, /* 2673 */
128'h230074696c70732d626c740065707974, /* 2674 */
128'h00736c6c65632d747075727265746e69, /* 2675 */
128'h6f72746e6f632d747075727265746e69, /* 2676 */
128'h646e6168702c78756e696c0072656c6c, /* 2677 */
128'h727265746e69007365676e617200656c, /* 2678 */
128'h6572006465646e657478652d73747075, /* 2679 */
128'h616d2c76637369720073656d616e2d67, /* 2680 */
128'h766373697200797469726f6972702d78, /* 2681 */
128'h70732d746e6572727563007665646e2c, /* 2682 */
128'h61702d747075727265746e6900646565, /* 2683 */
128'h0073747075727265746e6900746e6572, /* 2684 */
128'h6f692d6765720074666968732d676572, /* 2685 */
128'h63616d2d6c61636f6c0068746469772d, /* 2686 */
128'h0000000000000000737365726464612d, /* 2687 */
128'h0000000000203a642520656369766544, /* 2688 */
128'h00203a6425206563697665642073250a, /* 2689 */
128'h00000000203a6425206563697665440a, /* 2690 */
128'h000a656369766564206e776f6e6b6e75, /* 2691 */
128'h00000a2973252c73252870756b6f6f6c, /* 2692 */
128'h7265206c616e7265746e692070636864, /* 2693 */
128'h00000000000000000a7025202c726f72, /* 2694 */
128'h5145525f5043484420676e69646e6553, /* 2695 */
128'h4b434120504348440000000a54534555, /* 2696 */
128'h696c432050434844000000000000000a, /* 2697 */
128'h203a7373657264644120504920746e65, /* 2698 */
128'h0000000a64252e64252e64252e642520, /* 2699 */
128'h73657264644120504920726576726553, /* 2700 */
128'h0a64252e64252e64252e642520203a73, /* 2701 */
128'h6120726574756f520000000000000000, /* 2702 */
128'h252e64252e642520203a737365726464, /* 2703 */
128'h6b73616d2074654e0000000a64252e64, /* 2704 */
128'h64252e642520203a7373657264646120, /* 2705 */
128'h697420657361654c000a64252e64252e, /* 2706 */
128'h7364253a6d64253a686425203d20656d, /* 2707 */
128'h3d206e69616d6f44000000000000000a, /* 2708 */
128'h4820746e65696c4300000a2273252220, /* 2709 */
128'h000a22732522203d20656d616e74736f, /* 2710 */
128'h000000000a44455050494b53204b4341, /* 2711 */
128'h000000000000000a4b414e2050434844, /* 2712 */
128'h73657264646120646574736575716552, /* 2713 */
128'h0000000000000a646573756665722073, /* 2714 */
128'h000000000000000a732520726f727245, /* 2715 */
128'h6e6f6974706f2064656c646e61686e75, /* 2716 */
128'h656c646e61686e55000000000a642520, /* 2717 */
128'h64252065646f63706f20504348442064, /* 2718 */
128'h20676e69646e6553000000000000000a, /* 2719 */
128'h000a595245564f435349445f50434844, /* 2720 */
128'h00000000000a29732528726f72726570, /* 2721 */
128'h3a2043414d2073250000000030687465, /* 2722 */
128'h3a583230253a583230253a5832302520, /* 2723 */
128'h000a583230253a583230253a58323025, /* 2724 */
128'h484420646e65732074276e646c756f43, /* 2725 */
128'h206e6f20595245564f43534944205043, /* 2726 */
128'h00000a7325203a732520656369766564, /* 2727 */
128'h5043484420726f6620676e6974696157, /* 2728 */
128'h2020202020202020000a524546464f5f, /* 2729 */
128'h00000000000063250000000000000020, /* 2730 */
128'h0000005832302520000000000000002e, /* 2731 */
128'h00000000732573250000000000000a0a, /* 2732 */
128'h00000000007325203a646c697542202c, /* 2733 */
128'h73257a4820756c250000000000007325, /* 2734 */
128'h0000000000756c250000000000000000, /* 2735 */
128'h0073257a4863252000000000646c252e, /* 2736 */
128'h00000000007325736574794220756c25, /* 2737 */
128'h00003a786c3830250073254269632520, /* 2738 */
128'h000a73252020202000786c6c2a302520, /* 2739 */
128'h000000203a5d64255b6e6f6974636553, /* 2740 */
128'h727265207974696e6173207264646170, /* 2741 */
128'h2c7825286e666c6500000a702520726f, /* 2742 */
128'h000000000a3b29782578302c78257830, /* 2743 */
128'h782578302c302c7825287465736d656d, /* 2744 */
128'h464f5f4f4c43414d00000000000a3b29, /* 2745 */
128'h464f5f494843414d0000000054455346, /* 2746 */
128'h46464f5f524c50540000000054455346, /* 2747 */
128'h46464f5f534346540000000000544553, /* 2748 */
128'h4c5254434f49444d0000000000544553, /* 2749 */
128'h46464f5f534346520054455346464f5f, /* 2750 */
128'h5346464f5f5253520000000000544553, /* 2751 */
128'h46464f5f444142520000000000005445, /* 2752 */
128'h46464f5f524c50520000000000544553, /* 2753 */
128'h000000003f3f3f3f0000000000544553, /* 2754 */
128'h000064252b54455346464f5f524c5052, /* 2755 */
128'h6f746f72502050490000000000000047, /* 2756 */
128'h00000000000000000a50495049203d20, /* 2757 */
128'h6f746f72502050490000000000000054, /* 2758 */
128'h6f746f7250205049000a504745203d20, /* 2759 */
128'h6165682074736574000a505550203d20, /* 2760 */
128'h6e6f6320747365740000000a3a726564, /* 2761 */
128'h6f746f7250205049000a3a73746e6574, /* 2762 */
128'h6f746f7250205049000a504449203d20, /* 2763 */
128'h6f746f725020504900000a5054203d20, /* 2764 */
128'h00000000000000000a50434344203d20, /* 2765 */
128'h6f746f72502050490000000000000036, /* 2766 */
128'h00000000000000000a50565352203d20, /* 2767 */
128'h000a455247203d206f746f7250205049, /* 2768 */
128'h000a505345203d206f746f7250205049, /* 2769 */
128'h00000a4841203d206f746f7250205049, /* 2770 */
128'h000a50544d203d206f746f7250205049, /* 2771 */
128'h5054454542203d206f746f7250205049, /* 2772 */
128'h6f746f72502050490000000000000a48, /* 2773 */
128'h000000000000000a5041434e45203d20, /* 2774 */
128'h6f746f7250205049000000000000004d, /* 2775 */
128'h00000000000000000a504d4f43203d20, /* 2776 */
128'h0a50544353203d206f746f7250205049, /* 2777 */
128'h6f746f72502050490000000000000000, /* 2778 */
128'h00000000000a4554494c504455203d20, /* 2779 */
128'h0a534c504d203d206f746f7250205049, /* 2780 */
128'h6f746f72502050490000000000000000, /* 2781 */
128'h6f746f7270205049000a574152203d20, /* 2782 */
128'h2820646574726f707075736e75203d20, /* 2783 */
128'h79745f6f746f7270000000000a297825, /* 2784 */
128'h0000000000000a78257830203d206570, /* 2785 */
128'h727265746e692064656c646e61686e75, /* 2786 */
128'h414d2070757465530000000a21747075, /* 2787 */
128'h4d454f2049505351000a726464612043, /* 2788 */
128'h0000000000000a7825203d205d64255b, /* 2789 */
128'h00000a786c253a786c25203d2043414d, /* 2790 */
128'h3025203d20737365726464612043414d, /* 2791 */
128'h3230253a783230253a783230253a7832, /* 2792 */
128'h0000000a2e783230253a783230253a78, /* 2793 */
128'h75727265746e692074656e7265687445, /* 2794 */
128'h0a646c25203d20737574617473207470, /* 2795 */
128'h65687420746f6f420000000000000000, /* 2796 */
128'h2e6d6172676f727020646564616f6c20, /* 2797 */
128'h2c657962646f6f4700000000000a2e2e, /* 2798 */
128'h000000000a2e2e2e207265746f6f6220, /* 2799 */
128'h00007f7c5d5b3f3e3d3c3b3a2c2b2a22, /* 2800 */
128'h007f7c5d5b3f3e3d3c3b3a2e2c2b2a22, /* 2801 */
128'h66656463626139383736353433323130, /* 2802 */
128'h72776f6c2f6372730000000000000000, /* 2803 */
128'h00000000000000632e636d6d5f637369, /* 2804 */
128'h61625f6473203d3d20657361625f6473, /* 2805 */
128'h5f63736972776f6c00726464615f6573, /* 2806 */
128'h000a74756f656d6974207325203a6473, /* 2807 */
128'h616d202c6465766f6d65722064726143, /* 2808 */
128'h6425206f74206465676e616863206b73, /* 2809 */
128'h736e692064726143000000000000000a, /* 2810 */
128'h6e616863206b73616d202c6465747265, /* 2811 */
128'h0000000000000a6425206f7420646567, /* 2812 */
128'h25207461206465746165726320636d6d, /* 2813 */
128'h0000000a7825203d2074736f68202c78, /* 2814 */
128'h0000000000006f4e0000000000736559, /* 2815 */
128'h002020203a434d4d0000000052444420, /* 2816 */
128'h00000000000a7325203a656369766544, /* 2817 */
128'h3a4449207265727574636166756e614d, /* 2818 */
128'h0a7825203a4d454f000000000a782520, /* 2819 */
128'h6325203a656d614e0000000000000000, /* 2820 */
128'h0000000000000a206325632563256325, /* 2821 */
128'h00000a6425203a646565705320737542, /* 2822 */
128'h25203a79746963617061432068676948, /* 2823 */
128'h79746963617061430000000000000a73, /* 2824 */
128'h7464695720737542000000000000203a, /* 2825 */
128'h000000000a73257469622d6425203a68, /* 2826 */
128'h0000007825782520000000203a78250a, /* 2827 */
128'h00000000000064735f63736972776f6c, /* 2828 */
128'h0000000065646f6d206e776f6e6b6e55, /* 2829 */
128'h7830203a726f72724520737574617453, /* 2830 */
128'h2074756f656d69540000000a58383025, /* 2831 */
128'h616572206472616320676e6974696177, /* 2832 */
128'h6c69616620636d6d00000000000a7964, /* 2833 */
128'h6d6320706f747320646e6573206f7420, /* 2834 */
128'h6f6c62203a434d4d0000000000000a64, /* 2835 */
128'h20786c257830207265626d756e206b63, /* 2836 */
128'h6c2578302878616d2073646565637865, /* 2837 */
128'h203d3e20434d4d6500000000000a2978, /* 2838 */
128'h726f6620646572697571657220342e34, /* 2839 */
128'h642072657375206465636e61686e6520, /* 2840 */
128'h000000000000000a6165726120617461, /* 2841 */
128'h757320746f6e2073656f642064726143, /* 2842 */
128'h696e6f697469747261702074726f7070, /* 2843 */
128'h656f64206472614300000000000a676e, /* 2844 */
128'h20434820656e6966656420746f6e2073, /* 2845 */
128'h00000a657a69732070756f7267205057, /* 2846 */
128'h636e61686e6520617461642072657355, /* 2847 */
128'h5720434820746f6e2061657261206465, /* 2848 */
128'h696c6120657a69732070756f72672050, /* 2849 */
128'h72617020692550470000000a64656e67, /* 2850 */
128'h505720434820746f6e206e6f69746974, /* 2851 */
128'h67696c6120657a69732070756f726720, /* 2852 */
128'h656f642064726143000000000a64656e, /* 2853 */
128'h6e652074726f7070757320746f6e2073, /* 2854 */
128'h657475626972747461206465636e6168, /* 2855 */
128'h6e65206c61746f54000000000000000a, /* 2856 */
128'h6563786520657a6973206465636e6168, /* 2857 */
128'h20752528206d756d6978616d20736465, /* 2858 */
128'h656f64206472614300000a297525203e, /* 2859 */
128'h6f682074726f7070757320746f6e2073, /* 2860 */
128'h61702064656c6c6f72746e6f63207473, /* 2861 */
128'h6572206574697277206e6f6974697472, /* 2862 */
128'h6e6974746573207974696c696261696c, /* 2863 */
128'h726c61206472614300000000000a7367, /* 2864 */
128'h64656e6f697469747261702079646165, /* 2865 */
128'h206f6e203a434d4d000000000000000a, /* 2866 */
128'h0000000a746e65736572702064726163, /* 2867 */
128'h73657220746f6e206469642064726143, /* 2868 */
128'h20656761746c6f76206f7420646e6f70, /* 2869 */
128'h00000000000000000a217463656c6573, /* 2870 */
128'h7463656c6573206f7420656c62616e75, /* 2871 */
128'h00000000000000000a65646f6d206120, /* 2872 */
128'h646e756f66206473635f747865206f4e, /* 2873 */
128'h78363025206e614d0000000000000a21, /* 2874 */
128'h000000783430257834302520726e5320, /* 2875 */
128'h00000000632563256325632563256325, /* 2876 */
128'h6167656c20434d4d00000064252e6425, /* 2877 */
128'h636167654c2044530000000000007963, /* 2878 */
128'h6867694820434d4d0000000000000079, /* 2879 */
128'h0000297a484d36322820646565705320, /* 2880 */
128'h35282064656570532068676948204453, /* 2881 */
128'h6867694820434d4d000000297a484d30, /* 2882 */
128'h0000297a484d32352820646565705320, /* 2883 */
128'h7a484d32352820323552444420434d4d, /* 2884 */
128'h31524453205348550000000000000029, /* 2885 */
128'h00000000000000297a484d3532282032, /* 2886 */
128'h7a484d30352820353252445320534855, /* 2887 */
128'h35524453205348550000000000000029, /* 2888 */
128'h000000000000297a484d303031282030, /* 2889 */
128'h7a484d30352820303552444420534855, /* 2890 */
128'h31524453205348550000000000000029, /* 2891 */
128'h0000000000297a484d38303228203430, /* 2892 */
128'h0000297a484d30303228203030325348, /* 2893 */
128'h6f6e2064252065636976654420434d4d, /* 2894 */
128'h00000000000000000a646e756f662074, /* 2895 */
128'h00000000434d4d650000000000004453, /* 2896 */
128'h000000297325282000006425203a7325, /* 2897 */
128'h6e656c20656c69460000000000636d6d, /* 2898 */
128'h000000000000000a6425203d20687467, /* 2899 */
128'h0a7325203d202964252c70252835646d, /* 2900 */
128'h20747365757165520000000000000000, /* 2901 */
128'h25202e676e6f6c206f6f742068746170, /* 2902 */
128'h000000000000002f00000000000a646c, /* 2903 */
128'h6b636f6c62202c22732522203a717277, /* 2904 */
128'h00000000000000000a64253d657a6973, /* 2905 */
128'h646e6520656c69662065766965636552, /* 2906 */
128'h775f656c646e61680000000000000a2e, /* 2907 */
128'h00000000000a2e64656c6c6163207172, /* 2908 */
128'h65706f2050544654206c6167656c6c49, /* 2909 */
128'h00000000000000000a2e6e6f69746172, /* 2910 */
128'h25203d206465726975716572206e656c, /* 2911 */
128'h000a7825203d206c6175746361202c58, /* 2912 */
128'h206f74206c696146000000005c2d2f7c, /* 2913 */
128'h2172657669726420445320746e756f6d, /* 2914 */
128'h6f6f622064616f4c000000000000000a, /* 2915 */
128'h726f6d656d206f746e69206e69622e74, /* 2916 */
128'h6e69622e746f6f620000000000000a79, /* 2917 */
128'h742064656c6961460000000000000000, /* 2918 */
128'h0000000a21746f6f62206e65706f206f, /* 2919 */
128'h20524444206f7420666c652064616f6c, /* 2920 */
128'h6461657220666c65000a79726f6d656d, /* 2921 */
128'h646f6320687469772064656c69616620, /* 2922 */
128'h206f74206c6961660000000064252065, /* 2923 */
128'h000000000021656c69662065736f6c63, /* 2924 */
128'h6420746e756f6d75206f74206c696166, /* 2925 */
128'h20746f6f622d750a00000000216b7369, /* 2926 */
128'h67617473207473726966206465736162, /* 2927 */
128'h00000a726564616f6c20746f6f622065, /* 2928 */
128'h696166207325206e6f69747265737361, /* 2929 */
128'h696c202c732520656c6966202c64656c, /* 2930 */
128'h206e6f6974636e7566202c642520656e, /* 2931 */
128'h3a4552554c49414600000000000a7325, /* 2932 */
128'h74612078257830203d21207825783020, /* 2933 */
128'h00000a2e782578302074657366666f20, /* 2934 */
128'h7025203d203270202c7025203d203170, /* 2935 */
128'h2020202020202020000000000000000a, /* 2936 */
128'h08080808080808080000000000202020, /* 2937 */
128'h20676e69747465730000000000080808, /* 2938 */
128'h20676e69747365740000000000007525, /* 2939 */
128'h3a4552554c4941460000000000007525, /* 2940 */
128'h64612064616220656c626973736f7020, /* 2941 */
128'h666f20746120656e696c207373657264, /* 2942 */
128'h00000000000a2e782578302074657366, /* 2943 */
128'h7478656e206f7420676e697070696b53, /* 2944 */
128'h000000000000000a2e2e2e7473657420, /* 2945 */
128'h20202020200808080808080808080808, /* 2946 */
128'h08080808080808080808202020202020, /* 2947 */
128'h00000000000820080000000000000008, /* 2948 */
128'h78302073692065676e61722074736574, /* 2949 */
128'h00000000000a70257830206f74207025, /* 2950 */
128'h000000000075252f00752520706f6f4c, /* 2951 */
128'h6441206b637574530000000000000a3a, /* 2952 */
128'h0000203a732520200000007373657264, /* 2953 */
128'h00000a2e656e6f4400000000000a6b6f, /* 2954 */
128'h4d415244206c6174656d20657261420a, /* 2955 */
128'h65747365746d656d00000a7473657420, /* 2956 */
128'h20302e332e34206e6f69737265762072, /* 2957 */
128'h000000000000000a297469622d642528, /* 2958 */
128'h30322029432820746867697279706f43, /* 2959 */
128'h2073656c7261684320323130322d3130, /* 2960 */
128'h000000000000000a2e6e6f62617a6143, /* 2961 */
128'h74207265646e75206465736e6563694c, /* 2962 */
128'h50206c6172656e654720554e47206568, /* 2963 */
128'h65762065736e6563694c2063696c6275, /* 2964 */
128'h0a2e29796c6e6f282032206e6f697372, /* 2965 */
128'h5f676e696b726f770000000000000000, /* 2966 */
128'h20646c25202c424b6425203d20746573, /* 2967 */
128'h6c25202c736e6f697463757274736e69, /* 2968 */
128'h203d20495043202c73656c6379632064, /* 2969 */
128'h00000000000000000a646c252e646c25, /* 2970 */
128'h46454443424139383736353433323130, /* 2971 */
128'h6f57206f6c6c65480000000000000000, /* 2972 */
128'h205d64255b70777300000a0d21646c72, /* 2973 */
128'h73206863746977530000000a5825203d, /* 2974 */
128'h000a58252c5825203d20676e69747465, /* 2975 */
128'h5825203d2064656573206d6f646e6152, /* 2976 */
128'h0a746f6f62204453000000000000000a, /* 2977 */
128'h6f6f6220495053510000000000000000, /* 2978 */
128'h736574204d4152440000000000000a74, /* 2979 */
128'h6f6f6220505446540000000000000a74, /* 2980 */
128'h65742065686361430000000000000a74, /* 2981 */
128'h00000a0d7061727400000000000a7473, /* 2982 */
128'h00000002464c457fcccccccccccccccd, /* 2983 */
128'h1032547698badcfeefcdab8967452301, /* 2984 */
128'h5851f42d4c957f2d1000000020000000, /* 2985 */
128'haaaaaaaaaaaaaaaa5555555555555555, /* 2986 */
128'h00004b4d47545045000000030f060301, /* 2987 */
128'h000000003000000000000000004b4d47, /* 2988 */
128'h00000000ffffffff0000000000000000, /* 2989 */
128'h0000646d635f6473000000000c000000, /* 2990 */
128'h00000000bffeb36800006772615f6473, /* 2991 */
128'h000000000000000000000000cc33aa55, /* 2992 */
128'h00000000000000000000000000000000, /* 2993 */
128'h00000000000000000000000000000000, /* 2994 */
128'h00000000000000000000000000000000, /* 2995 */
128'h00000000000000000000000000000000, /* 2996 */
128'h00000000000000000000000000000000, /* 2997 */
128'h00000000000000000000000000000000, /* 2998 */
128'h00000000000000000000000000000000, /* 2999 */
128'h00000000000000000000000000000000, /* 3000 */
128'h00000000000000000000000000000000, /* 3001 */
128'h00000000000000000000000000000000, /* 3002 */
128'h00000000000000000000000000000000, /* 3003 */
128'h00000000000000000000000000000000, /* 3004 */
128'h00000000000000000000000000000000, /* 3005 */
128'h00000000000000000000000000000000, /* 3006 */
128'h00000000000000000000000000000000, /* 3007 */
128'h000000002f7c5c2d00000000ffffffff, /* 3008 */
128'hffffffff0000000600000000bffeb520, /* 3009 */
128'h00000000bffe70f40000000000000000, /* 3010 */
128'h000000000000000000000000000000b6, /* 3011 */
128'h00000000000000000000000000000000, /* 3012 */
128'h00000000000000000000000000000000, /* 3013 */
128'h00000000000000000000000000000000, /* 3014 */
128'h00000000000000000000000000000000, /* 3015 */
128'h00000000000000000000000000000000, /* 3016 */
128'h00000000000000000000000000000000, /* 3017 */
128'h00000000000000000000000000000000, /* 3018 */
128'h00000000000000000000000000000000, /* 3019 */
128'h00000000000000000000000000000000, /* 3020 */
128'h00000000000000000000000000000000, /* 3021 */
128'h00000000000000000000000000000000, /* 3022 */
128'h00000000000000000000000000000000, /* 3023 */
128'h00000000000000000000000000000000, /* 3024 */
128'h00000000000000000000000000000000, /* 3025 */
128'h00000000000000000000000000000000, /* 3026 */
128'h00000000000000000000000000000000, /* 3027 */
128'h00000000000000000000000000000000, /* 3028 */
128'h00000000000000000000000000000000, /* 3029 */
128'h00000000000000000000000000000000, /* 3030 */
128'h00000000000000000000000000000000, /* 3031 */
128'h00000000000000000000000000000000, /* 3032 */
128'h00000000000000000000000000000000, /* 3033 */
128'h00000000000000000000000000000000, /* 3034 */
128'h00000000000000000000000000000000, /* 3035 */
128'h00000000000000000000000000000000, /* 3036 */
128'h00000000000000000000000000000000, /* 3037 */
128'h00000000000000000000000000000000, /* 3038 */
128'h00000000000000000000000000000000, /* 3039 */
128'h00000000000000000000000000000000, /* 3040 */
128'h00000000000000000000000000000000, /* 3041 */
128'h00000000000000000000000000000000, /* 3042 */
128'h00000000000000000000000000000000, /* 3043 */
128'h00000000000000000000000000000000, /* 3044 */
128'h00000000000000000000000000000000, /* 3045 */
128'h00000000000000000000000000000000, /* 3046 */
128'h00000000000000000000000000000000, /* 3047 */
128'h00000000000000000000000000000000, /* 3048 */
128'h00000000000000000000000000000000, /* 3049 */
128'h00000000000000000000000000000000, /* 3050 */
128'h00000000000000000000000000000000, /* 3051 */
128'h00000000000000000000000000000000, /* 3052 */
128'h00000000000000000000000000000000, /* 3053 */
128'h00000000000000000000000000000000, /* 3054 */
128'h00000000000000000000000000000000, /* 3055 */
128'h00000000000000000000000000000000, /* 3056 */
128'h00000000000000000000000000000000, /* 3057 */
128'h00000000000000000000000000000000, /* 3058 */
128'h00000000000000000000000000000000, /* 3059 */
128'h00000000000000000000000000000000, /* 3060 */
128'h00000000000000000000000000000000, /* 3061 */
128'h00000000000000000000000000000000, /* 3062 */
128'h00000000000000000000000000000000, /* 3063 */
128'h00000000000000000000000000000000, /* 3064 */
128'h00000000000000000000000000000000, /* 3065 */
128'h00000000000000000000000000000000, /* 3066 */
128'h00000000000000000000000000000000, /* 3067 */
128'h00000000000000000000000000000000, /* 3068 */
128'h00000000000000000000000000000000, /* 3069 */
128'h00000000000000000000000000000000, /* 3070 */
128'h00000000000000000000000000000000, /* 3071 */
128'h00000000000000000000000000000000, /* 3072 */
128'h00000000000000000000000000000000, /* 3073 */
128'h00000000000000000000000000000000, /* 3074 */
128'h00000000000000000000000000000000, /* 3075 */
128'h00000000000000000000000000000000, /* 3076 */
128'h00000000000000000000000000000000, /* 3077 */
128'h00000000000000000000000000000000, /* 3078 */
128'h00000000000000000000000000000000, /* 3079 */
128'h00000000000000000000000000000000, /* 3080 */
128'h00000000000000000000000000000000, /* 3081 */
128'h00000000000000000000000000000000, /* 3082 */
128'h00000000000000000000000000000000, /* 3083 */
128'h00000000000000000000000000000000, /* 3084 */
128'h00000000000000000000000000000000, /* 3085 */
128'h00000000000000000000000000000000, /* 3086 */
128'h00000000000000000000000000000000, /* 3087 */
128'h00000000000000000000000000000000, /* 3088 */
128'h00000000000000000000000000000000, /* 3089 */
128'h00000000000000000000000000000000, /* 3090 */
128'h00000000000000000000000000000000, /* 3091 */
128'h00000000000000000000000000000000, /* 3092 */
128'h00000000000000000000000000000000, /* 3093 */
128'h00000000000000000000000000000000, /* 3094 */
128'h00000000000000000000000000000000, /* 3095 */
128'h00000000000000000000000000000000, /* 3096 */
128'h00000000000000000000000000000000, /* 3097 */
128'h00000000000000000000000000000000, /* 3098 */
128'h00000000000000000000000000000000, /* 3099 */
128'h00000000000000000000000000000000, /* 3100 */
128'h00000000000000000000000000000000, /* 3101 */
128'h00000000000000000000000000000000, /* 3102 */
128'h00000000000000000000000000000000, /* 3103 */
128'h00000000000000000000000000000000, /* 3104 */
128'h00000000000000000000000000000000, /* 3105 */
128'h00000000000000000000000000000000, /* 3106 */
128'h00000000000000000000000000000000, /* 3107 */
128'h00000000000000000000000000000000, /* 3108 */
128'h00000000000000000000000000000000, /* 3109 */
128'h00000000000000000000000000000000, /* 3110 */
128'h00000000000000000000000000000000, /* 3111 */
128'h00000000000000000000000000000000, /* 3112 */
128'h00000000000000000000000000000000, /* 3113 */
128'h00000000000000000000000000000000, /* 3114 */
128'h00000000000000000000000000000000, /* 3115 */
128'h00000000000000000000000000000000, /* 3116 */
128'h00000000000000000000000000000000, /* 3117 */
128'h00000000000000000000000000000000, /* 3118 */
128'h00000000000000000000000000000000, /* 3119 */
128'h00000000000000000000000000000000, /* 3120 */
128'h00000000000000000000000000000000, /* 3121 */
128'h00000000000000000000000000000000, /* 3122 */
128'h00000000000000000000000000000000, /* 3123 */
128'h00000000000000000000000000000000, /* 3124 */
128'h00000000000000000000000000000000, /* 3125 */
128'h00000000000000000000000000000000, /* 3126 */
128'h00000000000000000000000000000000, /* 3127 */
128'h00000000000000000000000000000000, /* 3128 */
128'h00000000000000000000000000000000, /* 3129 */
128'h00000000000000000000000000000000, /* 3130 */
128'h00000000000000000000000000000000, /* 3131 */
128'h00000000000000000000000000000000, /* 3132 */
128'h00000000000000000000000000000000, /* 3133 */
128'h00000000000000000000000000000000, /* 3134 */
128'h00000000000000000000000000000000, /* 3135 */
128'h00000000000000000000000000000000, /* 3136 */
128'h00000000000000000000000000000000, /* 3137 */
128'h00000000000000000000000000000000, /* 3138 */
128'h00000000000000000000000000000000, /* 3139 */
128'h00000000000000000000000000000000, /* 3140 */
128'h00000000000000000000000000000000, /* 3141 */
128'h00000000000000000000000000000000, /* 3142 */
128'h00000000000000000000000000000000, /* 3143 */
128'h00000000000000000000000000000000, /* 3144 */
128'h00000000000000000000000000000000, /* 3145 */
128'h00000000000000000000000000000000, /* 3146 */
128'h00000000000000000000000000000000, /* 3147 */
128'h00000000000000000000000000000000, /* 3148 */
128'h00000000000000000000000000000000, /* 3149 */
128'h00000000000000000000000000000000, /* 3150 */
128'h00000000000000000000000000000000, /* 3151 */
128'h00000000000000000000000000000000, /* 3152 */
128'h00000000000000000000000000000000, /* 3153 */
128'h00000000000000000000000000000000, /* 3154 */
128'h00000000000000000000000000000000, /* 3155 */
128'h00000000000000000000000000000000, /* 3156 */
128'h00000000000000000000000000000000, /* 3157 */
128'h00000000000000000000000000000000, /* 3158 */
128'h00000000000000000000000000000000, /* 3159 */
128'h00000000000000000000000000000000, /* 3160 */
128'h00000000000000000000000000000000, /* 3161 */
128'h00000000000000000000000000000000, /* 3162 */
128'h00000000000000000000000000000000, /* 3163 */
128'h00000000000000000000000000000000, /* 3164 */
128'h00000000000000000000000000000000, /* 3165 */
128'h00000000000000000000000000000000, /* 3166 */
128'h00000000000000000000000000000000, /* 3167 */
128'h00000000000000000000000000000000, /* 3168 */
128'h00000000000000000000000000000000, /* 3169 */
128'h00000000000000000000000000000000, /* 3170 */
128'h00000000000000000000000000000000, /* 3171 */
128'h00000000000000000000000000000000, /* 3172 */
128'h00000000000000000000000000000000, /* 3173 */
128'h00000000000000000000000000000000, /* 3174 */
128'h00000000000000000000000000000000, /* 3175 */
128'h00000000000000000000000000000000, /* 3176 */
128'h00000000000000000000000000000000, /* 3177 */
128'h00000000000000000000000000000000, /* 3178 */
128'h00000000000000000000000000000000, /* 3179 */
128'h00000000000000000000000000000000, /* 3180 */
128'h00000000000000000000000000000000, /* 3181 */
128'h00000000000000000000000000000000, /* 3182 */
128'h00000000000000000000000000000000, /* 3183 */
128'h00000000000000000000000000000000, /* 3184 */
128'h00000000000000000000000000000000, /* 3185 */
128'h00000000000000000000000000000000, /* 3186 */
128'h00000000000000000000000000000000, /* 3187 */
128'h00000000000000000000000000000000, /* 3188 */
128'h00000000000000000000000000000000, /* 3189 */
128'h00000000000000000000000000000000, /* 3190 */
128'h00000000000000000000000000000000, /* 3191 */
128'h00000000000000000000000000000000, /* 3192 */
128'h00000000000000000000000000000000, /* 3193 */
128'h00000000000000000000000000000000, /* 3194 */
128'h00000000000000000000000000000000, /* 3195 */
128'h00000000000000000000000000000000, /* 3196 */
128'h00000000000000000000000000000000, /* 3197 */
128'h00000000000000000000000000000000, /* 3198 */
128'h00000000000000000000000000000000, /* 3199 */
128'h00000000000000000000000000000000, /* 3200 */
128'h00000000000000000000000000000000, /* 3201 */
128'h00000000000000000000000000000000, /* 3202 */
128'h00000000000000000000000000000000, /* 3203 */
128'h00000000000000000000000000000000, /* 3204 */
128'h00000000000000000000000000000000, /* 3205 */
128'h00000000000000000000000000000000, /* 3206 */
128'h00000000000000000000000000000000, /* 3207 */
128'h00000000000000000000000000000000, /* 3208 */
128'h00000000000000000000000000000000, /* 3209 */
128'h00000000000000000000000000000000, /* 3210 */
128'h00000000000000000000000000000000, /* 3211 */
128'h00000000000000000000000000000000, /* 3212 */
128'h00000000000000000000000000000000, /* 3213 */
128'h00000000000000000000000000000000, /* 3214 */
128'h00000000000000000000000000000000, /* 3215 */
128'h00000000000000000000000000000000, /* 3216 */
128'h00000000000000000000000000000000, /* 3217 */
128'h00000000000000000000000000000000, /* 3218 */
128'h00000000000000000000000000000000, /* 3219 */
128'h00000000000000000000000000000000, /* 3220 */
128'h00000000000000000000000000000000, /* 3221 */
128'h00000000000000000000000000000000, /* 3222 */
128'h00000000000000000000000000000000, /* 3223 */
128'h00000000000000000000000000000000, /* 3224 */
128'h00000000000000000000000000000000, /* 3225 */
128'h00000000000000000000000000000000, /* 3226 */
128'h00000000000000000000000000000000, /* 3227 */
128'h00000000000000000000000000000000, /* 3228 */
128'h00000000000000000000000000000000, /* 3229 */
128'h00000000000000000000000000000000, /* 3230 */
128'h00000000000000000000000000000000, /* 3231 */
128'h00000000000000000000000000000000, /* 3232 */
128'h00000000000000000000000000000000, /* 3233 */
128'h00000000000000000000000000000000, /* 3234 */
128'h00000000000000000000000000000000, /* 3235 */
128'h00000000000000000000000000000000, /* 3236 */
128'h00000000000000000000000000000000, /* 3237 */
128'h00000000000000000000000000000000, /* 3238 */
128'h00000000000000000000000000000000, /* 3239 */
128'h00000000000000000000000000000000, /* 3240 */
128'h00000000000000000000000000000000, /* 3241 */
128'h00000000000000000000000000000000, /* 3242 */
128'h00000000000000000000000000000000, /* 3243 */
128'h00000000000000000000000000000000, /* 3244 */
128'h00000000000000000000000000000000, /* 3245 */
128'h00000000000000000000000000000000, /* 3246 */
128'h00000000000000000000000000000000, /* 3247 */
128'h00000000000000000000000000000000, /* 3248 */
128'h00000000000000000000000000000000, /* 3249 */
128'h00000000000000000000000000000000, /* 3250 */
128'h00000000000000000000000000000000, /* 3251 */
128'h00000000000000000000000000000000, /* 3252 */
128'h00000000000000000000000000000000, /* 3253 */
128'h00000000000000000000000000000000, /* 3254 */
128'h00000000000000000000000000000000, /* 3255 */
128'h00000000000000000000000000000000, /* 3256 */
128'h00000000000000000000000000000000, /* 3257 */
128'h00000000000000000000000000000000, /* 3258 */
128'h00000000000000000000000000000000, /* 3259 */
128'h00000000000000000000000000000000, /* 3260 */
128'h00000000000000000000000000000000, /* 3261 */
128'h00000000000000000000000000000000, /* 3262 */
128'h00000000000000000000000000000000, /* 3263 */
128'h00000000000000000000000000000000, /* 3264 */
128'h00000000000000000000000000000000, /* 3265 */
128'h00000000000000000000000000000000, /* 3266 */
128'h00000000000000000000000000000000, /* 3267 */
128'h00000000000000000000000000000000, /* 3268 */
128'h00000000000000000000000000000000, /* 3269 */
128'h00000000000000000000000000000000, /* 3270 */
128'h00000000000000000000000000000000, /* 3271 */
128'h00000000000000000000000000000000, /* 3272 */
128'h00000000000000000000000000000000, /* 3273 */
128'h00000000000000000000000000000000, /* 3274 */
128'h00000000000000000000000000000000, /* 3275 */
128'h00000000000000000000000000000000, /* 3276 */
128'h00000000000000000000000000000000, /* 3277 */
128'h00000000000000000000000000000000, /* 3278 */
128'h00000000000000000000000000000000, /* 3279 */
128'h00000000000000000000000000000000, /* 3280 */
128'h00000000000000000000000000000000, /* 3281 */
128'h00000000000000000000000000000000, /* 3282 */
128'h00000000000000000000000000000000, /* 3283 */
128'h00000000000000000000000000000000, /* 3284 */
128'h00000000000000000000000000000000, /* 3285 */
128'h00000000000000000000000000000000, /* 3286 */
128'h00000000000000000000000000000000, /* 3287 */
128'h00000000000000000000000000000000, /* 3288 */
128'h00000000000000000000000000000000, /* 3289 */
128'h00000000000000000000000000000000, /* 3290 */
128'h00000000000000000000000000000000, /* 3291 */
128'h00000000000000000000000000000000, /* 3292 */
128'h00000000000000000000000000000000, /* 3293 */
128'h00000000000000000000000000000000, /* 3294 */
128'h00000000000000000000000000000000, /* 3295 */
128'h00000000000000000000000000000000, /* 3296 */
128'h00000000000000000000000000000000, /* 3297 */
128'h00000000000000000000000000000000, /* 3298 */
128'h00000000000000000000000000000000, /* 3299 */
128'h00000000000000000000000000000000, /* 3300 */
128'h00000000000000000000000000000000, /* 3301 */
128'h00000000000000000000000000000000, /* 3302 */
128'h00000000000000000000000000000000, /* 3303 */
128'h00000000000000000000000000000000, /* 3304 */
128'h00000000000000000000000000000000, /* 3305 */
128'h00000000000000000000000000000000, /* 3306 */
128'h00000000000000000000000000000000, /* 3307 */
128'h00000000000000000000000000000000, /* 3308 */
128'h00000000000000000000000000000000, /* 3309 */
128'h00000000000000000000000000000000, /* 3310 */
128'h00000000000000000000000000000000, /* 3311 */
128'h00000000000000000000000000000000, /* 3312 */
128'h00000000000000000000000000000000, /* 3313 */
128'h00000000000000000000000000000000, /* 3314 */
128'h00000000000000000000000000000000, /* 3315 */
128'h00000000000000000000000000000000, /* 3316 */
128'h00000000000000000000000000000000, /* 3317 */
128'h00000000000000000000000000000000, /* 3318 */
128'h00000000000000000000000000000000, /* 3319 */
128'h00000000000000000000000000000000, /* 3320 */
128'h00000000000000000000000000000000, /* 3321 */
128'h00000000000000000000000000000000, /* 3322 */
128'h00000000000000000000000000000000, /* 3323 */
128'h00000000000000000000000000000000, /* 3324 */
128'h00000000000000000000000000000000, /* 3325 */
128'h00000000000000000000000000000000, /* 3326 */
128'h00000000000000000000000000000000, /* 3327 */
128'h00000000000000000000000000000000, /* 3328 */
128'h00000000000000000000000000000000, /* 3329 */
128'h00000000000000000000000000000000, /* 3330 */
128'h00000000000000000000000000000000, /* 3331 */
128'h00000000000000000000000000000000, /* 3332 */
128'h00000000000000000000000000000000, /* 3333 */
128'h00000000000000000000000000000000, /* 3334 */
128'h00000000000000000000000000000000, /* 3335 */
128'h00000000000000000000000000000000, /* 3336 */
128'h00000000000000000000000000000000, /* 3337 */
128'h00000000000000000000000000000000, /* 3338 */
128'h00000000000000000000000000000000, /* 3339 */
128'h00000000000000000000000000000000, /* 3340 */
128'h00000000000000000000000000000000, /* 3341 */
128'h00000000000000000000000000000000, /* 3342 */
128'h00000000000000000000000000000000, /* 3343 */
128'h00000000000000000000000000000000, /* 3344 */
128'h00000000000000000000000000000000, /* 3345 */
128'h00000000000000000000000000000000, /* 3346 */
128'h00000000000000000000000000000000, /* 3347 */
128'h00000000000000000000000000000000, /* 3348 */
128'h00000000000000000000000000000000, /* 3349 */
128'h00000000000000000000000000000000, /* 3350 */
128'h00000000000000000000000000000000, /* 3351 */
128'h00000000000000000000000000000000, /* 3352 */
128'h00000000000000000000000000000000, /* 3353 */
128'h00000000000000000000000000000000, /* 3354 */
128'h00000000000000000000000000000000, /* 3355 */
128'h00000000000000000000000000000000, /* 3356 */
128'h00000000000000000000000000000000, /* 3357 */
128'h00000000000000000000000000000000, /* 3358 */
128'h00000000000000000000000000000000, /* 3359 */
128'h00000000000000000000000000000000, /* 3360 */
128'h00000000000000000000000000000000, /* 3361 */
128'h00000000000000000000000000000000, /* 3362 */
128'h00000000000000000000000000000000, /* 3363 */
128'h00000000000000000000000000000000, /* 3364 */
128'h00000000000000000000000000000000, /* 3365 */
128'h00000000000000000000000000000000, /* 3366 */
128'h00000000000000000000000000000000, /* 3367 */
128'h00000000000000000000000000000000, /* 3368 */
128'h00000000000000000000000000000000, /* 3369 */
128'h00000000000000000000000000000000, /* 3370 */
128'h00000000000000000000000000000000, /* 3371 */
128'h00000000000000000000000000000000, /* 3372 */
128'h00000000000000000000000000000000, /* 3373 */
128'h00000000000000000000000000000000, /* 3374 */
128'h00000000000000000000000000000000, /* 3375 */
128'h00000000000000000000000000000000, /* 3376 */
128'h00000000000000000000000000000000, /* 3377 */
128'h00000000000000000000000000000000, /* 3378 */
128'h00000000000000000000000000000000, /* 3379 */
128'h00000000000000000000000000000000, /* 3380 */
128'h00000000000000000000000000000000, /* 3381 */
128'h00000000000000000000000000000000, /* 3382 */
128'h00000000000000000000000000000000, /* 3383 */
128'h00000000000000000000000000000000, /* 3384 */
128'h00000000000000000000000000000000, /* 3385 */
128'h00000000000000000000000000000000, /* 3386 */
128'h00000000000000000000000000000000, /* 3387 */
128'h00000000000000000000000000000000, /* 3388 */
128'h00000000000000000000000000000000, /* 3389 */
128'h00000000000000000000000000000000, /* 3390 */
128'h00000000000000000000000000000000, /* 3391 */
128'h00000000000000000000000000000000, /* 3392 */
128'h00000000000000000000000000000000, /* 3393 */
128'h00000000000000000000000000000000, /* 3394 */
128'h00000000000000000000000000000000, /* 3395 */
128'h00000000000000000000000000000000, /* 3396 */
128'h00000000000000000000000000000000, /* 3397 */
128'h00000000000000000000000000000000, /* 3398 */
128'h00000000000000000000000000000000, /* 3399 */
128'h00000000000000000000000000000000, /* 3400 */
128'h00000000000000000000000000000000, /* 3401 */
128'h00000000000000000000000000000000, /* 3402 */
128'h00000000000000000000000000000000, /* 3403 */
128'h00000000000000000000000000000000, /* 3404 */
128'h00000000000000000000000000000000, /* 3405 */
128'h00000000000000000000000000000000, /* 3406 */
128'h00000000000000000000000000000000, /* 3407 */
128'h00000000000000000000000000000000, /* 3408 */
128'h00000000000000000000000000000000, /* 3409 */
128'h00000000000000000000000000000000, /* 3410 */
128'h00000000000000000000000000000000, /* 3411 */
128'h00000000000000000000000000000000, /* 3412 */
128'h00000000000000000000000000000000, /* 3413 */
128'h00000000000000000000000000000000, /* 3414 */
128'h00000000000000000000000000000000, /* 3415 */
128'h00000000000000000000000000000000, /* 3416 */
128'h00000000000000000000000000000000, /* 3417 */
128'h00000000000000000000000000000000, /* 3418 */
128'h00000000000000000000000000000000, /* 3419 */
128'h00000000000000000000000000000000, /* 3420 */
128'h00000000000000000000000000000000, /* 3421 */
128'h00000000000000000000000000000000, /* 3422 */
128'h00000000000000000000000000000000, /* 3423 */
128'h00000000000000000000000000000000, /* 3424 */
128'h00000000000000000000000000000000, /* 3425 */
128'h00000000000000000000000000000000, /* 3426 */
128'h00000000000000000000000000000000, /* 3427 */
128'h00000000000000000000000000000000, /* 3428 */
128'h00000000000000000000000000000000, /* 3429 */
128'h00000000000000000000000000000000, /* 3430 */
128'h00000000000000000000000000000000, /* 3431 */
128'h00000000000000000000000000000000, /* 3432 */
128'h00000000000000000000000000000000, /* 3433 */
128'h00000000000000000000000000000000, /* 3434 */
128'h00000000000000000000000000000000, /* 3435 */
128'h00000000000000000000000000000000, /* 3436 */
128'h00000000000000000000000000000000, /* 3437 */
128'h00000000000000000000000000000000, /* 3438 */
128'h00000000000000000000000000000000, /* 3439 */
128'h00000000000000000000000000000000, /* 3440 */
128'h00000000000000000000000000000000, /* 3441 */
128'h00000000000000000000000000000000, /* 3442 */
128'h00000000000000000000000000000000, /* 3443 */
128'h00000000000000000000000000000000, /* 3444 */
128'h00000000000000000000000000000000, /* 3445 */
128'h00000000000000000000000000000000, /* 3446 */
128'h00000000000000000000000000000000, /* 3447 */
128'h00000000000000000000000000000000, /* 3448 */
128'h00000000000000000000000000000000, /* 3449 */
128'h00000000000000000000000000000000, /* 3450 */
128'h00000000000000000000000000000000, /* 3451 */
128'h00000000000000000000000000000000, /* 3452 */
128'h00000000000000000000000000000000, /* 3453 */
128'h00000000000000000000000000000000, /* 3454 */
128'h00000000000000000000000000000000, /* 3455 */
128'h00000000000000000000000000000000, /* 3456 */
128'h00000000000000000000000000000000, /* 3457 */
128'h00000000000000000000000000000000, /* 3458 */
128'h00000000000000000000000000000000, /* 3459 */
128'h00000000000000000000000000000000, /* 3460 */
128'h00000000000000000000000000000000, /* 3461 */
128'h00000000000000000000000000000000, /* 3462 */
128'h00000000000000000000000000000000, /* 3463 */
128'h00000000000000000000000000000000, /* 3464 */
128'h00000000000000000000000000000000, /* 3465 */
128'h00000000000000000000000000000000, /* 3466 */
128'h00000000000000000000000000000000, /* 3467 */
128'h00000000000000000000000000000000, /* 3468 */
128'h00000000000000000000000000000000, /* 3469 */
128'h00000000000000000000000000000000, /* 3470 */
128'h00000000000000000000000000000000, /* 3471 */
128'h00000000000000000000000000000000, /* 3472 */
128'h00000000000000000000000000000000, /* 3473 */
128'h00000000000000000000000000000000, /* 3474 */
128'h00000000000000000000000000000000, /* 3475 */
128'h00000000000000000000000000000000, /* 3476 */
128'h00000000000000000000000000000000, /* 3477 */
128'h00000000000000000000000000000000, /* 3478 */
128'h00000000000000000000000000000000, /* 3479 */
128'h00000000000000000000000000000000, /* 3480 */
128'h00000000000000000000000000000000, /* 3481 */
128'h00000000000000000000000000000000, /* 3482 */
128'h00000000000000000000000000000000, /* 3483 */
128'h00000000000000000000000000000000, /* 3484 */
128'h00000000000000000000000000000000, /* 3485 */
128'h00000000000000000000000000000000, /* 3486 */
128'h00000000000000000000000000000000, /* 3487 */
128'h00000000000000000000000000000000, /* 3488 */
128'h00000000000000000000000000000000, /* 3489 */
128'h00000000000000000000000000000000, /* 3490 */
128'h00000000000000000000000000000000, /* 3491 */
128'h00000000000000000000000000000000, /* 3492 */
128'h00000000000000000000000000000000, /* 3493 */
128'h00000000000000000000000000000000, /* 3494 */
128'h00000000000000000000000000000000, /* 3495 */
128'h00000000000000000000000000000000, /* 3496 */
128'h00000000000000000000000000000000, /* 3497 */
128'h00000000000000000000000000000000, /* 3498 */
128'h00000000000000000000000000000000, /* 3499 */
128'h00000000000000000000000000000000, /* 3500 */
128'h00000000000000000000000000000000, /* 3501 */
128'h00000000000000000000000000000000, /* 3502 */
128'h00000000000000000000000000000000, /* 3503 */
128'h00000000000000000000000000000000, /* 3504 */
128'h00000000000000000000000000000000, /* 3505 */
128'h00000000000000000000000000000000, /* 3506 */
128'h00000000000000000000000000000000, /* 3507 */
128'h00000000000000000000000000000000, /* 3508 */
128'h00000000000000000000000000000000, /* 3509 */
128'h00000000000000000000000000000000, /* 3510 */
128'h00000000000000000000000000000000, /* 3511 */
128'h00000000000000000000000000000000, /* 3512 */
128'h00000000000000000000000000000000, /* 3513 */
128'h00000000000000000000000000000000, /* 3514 */
128'h00000000000000000000000000000000, /* 3515 */
128'h00000000000000000000000000000000, /* 3516 */
128'h00000000000000000000000000000000, /* 3517 */
128'h00000000000000000000000000000000, /* 3518 */
128'h00000000000000000000000000000000, /* 3519 */
128'h00000000000000000000000000000000, /* 3520 */
128'h00000000000000000000000000000000, /* 3521 */
128'h00000000000000000000000000000000, /* 3522 */
128'h00000000000000000000000000000000, /* 3523 */
128'h00000000000000000000000000000000, /* 3524 */
128'h00000000000000000000000000000000, /* 3525 */
128'h00000000000000000000000000000000, /* 3526 */
128'h00000000000000000000000000000000, /* 3527 */
128'h00000000000000000000000000000000, /* 3528 */
128'h00000000000000000000000000000000, /* 3529 */
128'h00000000000000000000000000000000, /* 3530 */
128'h00000000000000000000000000000000, /* 3531 */
128'h00000000000000000000000000000000, /* 3532 */
128'h00000000000000000000000000000000, /* 3533 */
128'h00000000000000000000000000000000, /* 3534 */
128'h00000000000000000000000000000000, /* 3535 */
128'h00000000000000000000000000000000, /* 3536 */
128'h00000000000000000000000000000000, /* 3537 */
128'h00000000000000000000000000000000, /* 3538 */
128'h00000000000000000000000000000000, /* 3539 */
128'h00000000000000000000000000000000, /* 3540 */
128'h00000000000000000000000000000000, /* 3541 */
128'h00000000000000000000000000000000, /* 3542 */
128'h00000000000000000000000000000000, /* 3543 */
128'h00000000000000000000000000000000, /* 3544 */
128'h00000000000000000000000000000000, /* 3545 */
128'h00000000000000000000000000000000, /* 3546 */
128'h00000000000000000000000000000000, /* 3547 */
128'h00000000000000000000000000000000, /* 3548 */
128'h00000000000000000000000000000000, /* 3549 */
128'h00000000000000000000000000000000, /* 3550 */
128'h00000000000000000000000000000000, /* 3551 */
128'h00000000000000000000000000000000, /* 3552 */
128'h00000000000000000000000000000000, /* 3553 */
128'h00000000000000000000000000000000, /* 3554 */
128'h00000000000000000000000000000000, /* 3555 */
128'h00000000000000000000000000000000, /* 3556 */
128'h00000000000000000000000000000000, /* 3557 */
128'h00000000000000000000000000000000, /* 3558 */
128'h00000000000000000000000000000000, /* 3559 */
128'h00000000000000000000000000000000, /* 3560 */
128'h00000000000000000000000000000000, /* 3561 */
128'h00000000000000000000000000000000, /* 3562 */
128'h00000000000000000000000000000000, /* 3563 */
128'h00000000000000000000000000000000, /* 3564 */
128'h00000000000000000000000000000000, /* 3565 */
128'h00000000000000000000000000000000, /* 3566 */
128'h00000000000000000000000000000000, /* 3567 */
128'h00000000000000000000000000000000, /* 3568 */
128'h00000000000000000000000000000000, /* 3569 */
128'h00000000000000000000000000000000, /* 3570 */
128'h00000000000000000000000000000000, /* 3571 */
128'h00000000000000000000000000000000, /* 3572 */
128'h00000000000000000000000000000000, /* 3573 */
128'h00000000000000000000000000000000, /* 3574 */
128'h00000000000000000000000000000000, /* 3575 */
128'h00000000000000000000000000000000, /* 3576 */
128'h00000000000000000000000000000000, /* 3577 */
128'h00000000000000000000000000000000, /* 3578 */
128'h00000000000000000000000000000000, /* 3579 */
128'h00000000000000000000000000000000, /* 3580 */
128'h00000000000000000000000000000000, /* 3581 */
128'h00000000000000000000000000000000, /* 3582 */
128'h00000000000000000000000000000000, /* 3583 */
128'h00000000000000000000000000000000, /* 3584 */
128'h00000000000000000000000000000000, /* 3585 */
128'h00000000000000000000000000000000, /* 3586 */
128'h00000000000000000000000000000000, /* 3587 */
128'h00000000000000000000000000000000, /* 3588 */
128'h00000000000000000000000000000000, /* 3589 */
128'h00000000000000000000000000000000, /* 3590 */
128'h00000000000000000000000000000000, /* 3591 */
128'h00000000000000000000000000000000, /* 3592 */
128'h00000000000000000000000000000000, /* 3593 */
128'h00000000000000000000000000000000, /* 3594 */
128'h00000000000000000000000000000000, /* 3595 */
128'h00000000000000000000000000000000, /* 3596 */
128'h00000000000000000000000000000000, /* 3597 */
128'h00000000000000000000000000000000, /* 3598 */
128'h00000000000000000000000000000000, /* 3599 */
128'h00000000000000000000000000000000, /* 3600 */
128'h00000000000000000000000000000000, /* 3601 */
128'h00000000000000000000000000000000, /* 3602 */
128'h00000000000000000000000000000000, /* 3603 */
128'h00000000000000000000000000000000, /* 3604 */
128'h00000000000000000000000000000000, /* 3605 */
128'h00000000000000000000000000000000, /* 3606 */
128'h00000000000000000000000000000000, /* 3607 */
128'h00000000000000000000000000000000, /* 3608 */
128'h00000000000000000000000000000000, /* 3609 */
128'h00000000000000000000000000000000, /* 3610 */
128'h00000000000000000000000000000000, /* 3611 */
128'h00000000000000000000000000000000, /* 3612 */
128'h00000000000000000000000000000000, /* 3613 */
128'h00000000000000000000000000000000, /* 3614 */
128'h00000000000000000000000000000000, /* 3615 */
128'h00000000000000000000000000000000, /* 3616 */
128'h00000000000000000000000000000000, /* 3617 */
128'h00000000000000000000000000000000, /* 3618 */
128'h00000000000000000000000000000000, /* 3619 */
128'h00000000000000000000000000000000, /* 3620 */
128'h00000000000000000000000000000000, /* 3621 */
128'h00000000000000000000000000000000, /* 3622 */
128'h00000000000000000000000000000000, /* 3623 */
128'h00000000000000000000000000000000, /* 3624 */
128'h00000000000000000000000000000000, /* 3625 */
128'h00000000000000000000000000000000, /* 3626 */
128'h00000000000000000000000000000000, /* 3627 */
128'h00000000000000000000000000000000, /* 3628 */
128'h00000000000000000000000000000000, /* 3629 */
128'h00000000000000000000000000000000, /* 3630 */
128'h00000000000000000000000000000000, /* 3631 */
128'h00000000000000000000000000000000, /* 3632 */
128'h00000000000000000000000000000000, /* 3633 */
128'h00000000000000000000000000000000, /* 3634 */
128'h00000000000000000000000000000000, /* 3635 */
128'h00000000000000000000000000000000, /* 3636 */
128'h00000000000000000000000000000000, /* 3637 */
128'h00000000000000000000000000000000, /* 3638 */
128'h00000000000000000000000000000000, /* 3639 */
128'h00000000000000000000000000000000, /* 3640 */
128'h00000000000000000000000000000000, /* 3641 */
128'h00000000000000000000000000000000, /* 3642 */
128'h00000000000000000000000000000000, /* 3643 */
128'h00000000000000000000000000000000, /* 3644 */
128'h00000000000000000000000000000000, /* 3645 */
128'h00000000000000000000000000000000, /* 3646 */
128'h00000000000000000000000000000000, /* 3647 */
128'h00000000000000000000000000000000, /* 3648 */
128'h00000000000000000000000000000000, /* 3649 */
128'h00000000000000000000000000000000, /* 3650 */
128'h00000000000000000000000000000000, /* 3651 */
128'h00000000000000000000000000000000, /* 3652 */
128'h00000000000000000000000000000000, /* 3653 */
128'h00000000000000000000000000000000, /* 3654 */
128'h00000000000000000000000000000000, /* 3655 */
128'h00000000000000000000000000000000, /* 3656 */
128'h00000000000000000000000000000000, /* 3657 */
128'h00000000000000000000000000000000, /* 3658 */
128'h00000000000000000000000000000000, /* 3659 */
128'h00000000000000000000000000000000, /* 3660 */
128'h00000000000000000000000000000000, /* 3661 */
128'h00000000000000000000000000000000, /* 3662 */
128'h00000000000000000000000000000000, /* 3663 */
128'h00000000000000000000000000000000, /* 3664 */
128'h00000000000000000000000000000000, /* 3665 */
128'h00000000000000000000000000000000, /* 3666 */
128'h00000000000000000000000000000000, /* 3667 */
128'h00000000000000000000000000000000, /* 3668 */
128'h00000000000000000000000000000000, /* 3669 */
128'h00000000000000000000000000000000, /* 3670 */
128'h00000000000000000000000000000000, /* 3671 */
128'h00000000000000000000000000000000, /* 3672 */
128'h00000000000000000000000000000000, /* 3673 */
128'h00000000000000000000000000000000, /* 3674 */
128'h00000000000000000000000000000000, /* 3675 */
128'h00000000000000000000000000000000, /* 3676 */
128'h00000000000000000000000000000000, /* 3677 */
128'h00000000000000000000000000000000, /* 3678 */
128'h00000000000000000000000000000000, /* 3679 */
128'h00000000000000000000000000000000, /* 3680 */
128'h00000000000000000000000000000000, /* 3681 */
128'h00000000000000000000000000000000, /* 3682 */
128'h00000000000000000000000000000000, /* 3683 */
128'h00000000000000000000000000000000, /* 3684 */
128'h00000000000000000000000000000000, /* 3685 */
128'h00000000000000000000000000000000, /* 3686 */
128'h00000000000000000000000000000000, /* 3687 */
128'h00000000000000000000000000000000, /* 3688 */
128'h00000000000000000000000000000000, /* 3689 */
128'h00000000000000000000000000000000, /* 3690 */
128'h00000000000000000000000000000000, /* 3691 */
128'h00000000000000000000000000000000, /* 3692 */
128'h00000000000000000000000000000000, /* 3693 */
128'h00000000000000000000000000000000, /* 3694 */
128'h00000000000000000000000000000000, /* 3695 */
128'h00000000000000000000000000000000, /* 3696 */
128'h00000000000000000000000000000000, /* 3697 */
128'h00000000000000000000000000000000, /* 3698 */
128'h00000000000000000000000000000000, /* 3699 */
128'h00000000000000000000000000000000, /* 3700 */
128'h00000000000000000000000000000000, /* 3701 */
128'h00000000000000000000000000000000, /* 3702 */
128'h00000000000000000000000000000000, /* 3703 */
128'h00000000000000000000000000000000, /* 3704 */
128'h00000000000000000000000000000000, /* 3705 */
128'h00000000000000000000000000000000, /* 3706 */
128'h00000000000000000000000000000000, /* 3707 */
128'h00000000000000000000000000000000, /* 3708 */
128'h00000000000000000000000000000000, /* 3709 */
128'h00000000000000000000000000000000, /* 3710 */
128'h00000000000000000000000000000000, /* 3711 */
128'h00000000000000000000000000000000, /* 3712 */
128'h00000000000000000000000000000000, /* 3713 */
128'h00000000000000000000000000000000, /* 3714 */
128'h00000000000000000000000000000000, /* 3715 */
128'h00000000000000000000000000000000, /* 3716 */
128'h00000000000000000000000000000000, /* 3717 */
128'h00000000000000000000000000000000, /* 3718 */
128'h00000000000000000000000000000000, /* 3719 */
128'h00000000000000000000000000000000, /* 3720 */
128'h00000000000000000000000000000000, /* 3721 */
128'h00000000000000000000000000000000, /* 3722 */
128'h00000000000000000000000000000000, /* 3723 */
128'h00000000000000000000000000000000, /* 3724 */
128'h00000000000000000000000000000000, /* 3725 */
128'h00000000000000000000000000000000, /* 3726 */
128'h00000000000000000000000000000000, /* 3727 */
128'h00000000000000000000000000000000, /* 3728 */
128'h00000000000000000000000000000000, /* 3729 */
128'h00000000000000000000000000000000, /* 3730 */
128'h00000000000000000000000000000000, /* 3731 */
128'h00000000000000000000000000000000, /* 3732 */
128'h00000000000000000000000000000000, /* 3733 */
128'h00000000000000000000000000000000, /* 3734 */
128'h00000000000000000000000000000000, /* 3735 */
128'h00000000000000000000000000000000, /* 3736 */
128'h00000000000000000000000000000000, /* 3737 */
128'h00000000000000000000000000000000, /* 3738 */
128'h00000000000000000000000000000000, /* 3739 */
128'h00000000000000000000000000000000, /* 3740 */
128'h00000000000000000000000000000000, /* 3741 */
128'h00000000000000000000000000000000, /* 3742 */
128'h00000000000000000000000000000000, /* 3743 */
128'h00000000000000000000000000000000, /* 3744 */
128'h00000000000000000000000000000000, /* 3745 */
128'h00000000000000000000000000000000, /* 3746 */
128'h00000000000000000000000000000000, /* 3747 */
128'h00000000000000000000000000000000, /* 3748 */
128'h00000000000000000000000000000000, /* 3749 */
128'h00000000000000000000000000000000, /* 3750 */
128'h00000000000000000000000000000000, /* 3751 */
128'h00000000000000000000000000000000, /* 3752 */
128'h00000000000000000000000000000000, /* 3753 */
128'h00000000000000000000000000000000, /* 3754 */
128'h00000000000000000000000000000000, /* 3755 */
128'h00000000000000000000000000000000, /* 3756 */
128'h00000000000000000000000000000000, /* 3757 */
128'h00000000000000000000000000000000, /* 3758 */
128'h00000000000000000000000000000000, /* 3759 */
128'h00000000000000000000000000000000, /* 3760 */
128'h00000000000000000000000000000000, /* 3761 */
128'h00000000000000000000000000000000, /* 3762 */
128'h00000000000000000000000000000000, /* 3763 */
128'h00000000000000000000000000000000, /* 3764 */
128'h00000000000000000000000000000000, /* 3765 */
128'h00000000000000000000000000000000, /* 3766 */
128'h00000000000000000000000000000000, /* 3767 */
128'h00000000000000000000000000000000, /* 3768 */
128'h00000000000000000000000000000000, /* 3769 */
128'h00000000000000000000000000000000, /* 3770 */
128'h00000000000000000000000000000000, /* 3771 */
128'h00000000000000000000000000000000, /* 3772 */
128'h00000000000000000000000000000000, /* 3773 */
128'h00000000000000000000000000000000, /* 3774 */
128'h00000000000000000000000000000000, /* 3775 */
128'h00000000000000000000000000000000, /* 3776 */
128'h00000000000000000000000000000000, /* 3777 */
128'h00000000000000000000000000000000, /* 3778 */
128'h00000000000000000000000000000000, /* 3779 */
128'h00000000000000000000000000000000, /* 3780 */
128'h00000000000000000000000000000000, /* 3781 */
128'h00000000000000000000000000000000, /* 3782 */
128'h00000000000000000000000000000000, /* 3783 */
128'h00000000000000000000000000000000, /* 3784 */
128'h00000000000000000000000000000000, /* 3785 */
128'h00000000000000000000000000000000, /* 3786 */
128'h00000000000000000000000000000000, /* 3787 */
128'h00000000000000000000000000000000, /* 3788 */
128'h00000000000000000000000000000000, /* 3789 */
128'h00000000000000000000000000000000, /* 3790 */
128'h00000000000000000000000000000000, /* 3791 */
128'h00000000000000000000000000000000, /* 3792 */
128'h00000000000000000000000000000000, /* 3793 */
128'h00000000000000000000000000000000, /* 3794 */
128'h00000000000000000000000000000000, /* 3795 */
128'h00000000000000000000000000000000, /* 3796 */
128'h00000000000000000000000000000000, /* 3797 */
128'h00000000000000000000000000000000, /* 3798 */
128'h00000000000000000000000000000000, /* 3799 */
128'h00000000000000000000000000000000, /* 3800 */
128'h00000000000000000000000000000000, /* 3801 */
128'h00000000000000000000000000000000, /* 3802 */
128'h00000000000000000000000000000000, /* 3803 */
128'h00000000000000000000000000000000, /* 3804 */
128'h00000000000000000000000000000000, /* 3805 */
128'h00000000000000000000000000000000, /* 3806 */
128'h00000000000000000000000000000000, /* 3807 */
128'h00000000000000000000000000000000, /* 3808 */
128'h00000000000000000000000000000000, /* 3809 */
128'h00000000000000000000000000000000, /* 3810 */
128'h00000000000000000000000000000000, /* 3811 */
128'h00000000000000000000000000000000, /* 3812 */
128'h00000000000000000000000000000000, /* 3813 */
128'h00000000000000000000000000000000, /* 3814 */
128'h00000000000000000000000000000000, /* 3815 */
128'h00000000000000000000000000000000, /* 3816 */
128'h00000000000000000000000000000000, /* 3817 */
128'h00000000000000000000000000000000, /* 3818 */
128'h00000000000000000000000000000000, /* 3819 */
128'h00000000000000000000000000000000, /* 3820 */
128'h00000000000000000000000000000000, /* 3821 */
128'h00000000000000000000000000000000, /* 3822 */
128'h00000000000000000000000000000000, /* 3823 */
128'h00000000000000000000000000000000, /* 3824 */
128'h00000000000000000000000000000000, /* 3825 */
128'h00000000000000000000000000000000, /* 3826 */
128'h00000000000000000000000000000000, /* 3827 */
128'h00000000000000000000000000000000, /* 3828 */
128'h00000000000000000000000000000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00000000000000000000000000000000, /* 3840 */
128'h00000000000000000000000000000000, /* 3841 */
128'h00000000000000000000000000000000, /* 3842 */
128'h00000000000000000000000000000000, /* 3843 */
128'h00000000000000000000000000000000, /* 3844 */
128'h00000000000000000000000000000000, /* 3845 */
128'h00000000000000000000000000000000, /* 3846 */
128'h00000000000000000000000000000000, /* 3847 */
128'h00000000000000000000000000000000, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule

