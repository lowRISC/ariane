/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'hfffe8e93100e8e9b05f5eeb711249c63, /*    1 */
128'h011111133ff1011b00004137fe0e9ee3, /*    2 */
128'h00008297000280e70ce2829300008297, /*    3 */
128'h000280e713050513000005170f428293, /*    4 */
128'hbb5606130000c617fb05859300000597, /*    5 */
128'h000f4eb7011696933ff6869b000046b7, /*    6 */
128'h0085b703fffe8e930005b703240e8e9b, /*    7 */
128'hff81011301b111130110011bfe0e9ae3, /*    8 */
128'h0085b70300e6b0230005b7030006b703, /*    9 */
128'h0185b70300e6b8230105b70300e6b423, /*   10 */
128'hfcc5cce3020686930205859300e6bc23, /*   11 */
128'h40b787b300d787b30147879300000797, /*   12 */
128'h30579073090787930000079700078067, /*   13 */
128'h3b8606130000c617c20585930000c597, /*   14 */
128'h0005bc230005b8230005b4230005b023, /*   15 */
128'h020004b703f090effec5c6e302058593, /*   16 */
128'h02000937004484930124a02300100913, /*   17 */
128'h3440297310500073ff24c6e34009091b, /*   18 */
128'hf1402973020004b7fe090ae300897913, /*   19 */
128'h0004a903000920230099093300291913, /*   20 */
128'h4009091b0200093700448493fe091ee3, /*   21 */
128'h1050007334102373342022f3ff24c6e3, /*   22 */
128'h41206d6f7266206f6c6c6548ffdff06f, /*   23 */
128'h617720657361656c502021656e616972, /*   24 */
128'h000a2e2e2e746e656d6f6d2061207469, /*   25 */
128'h00000000000000000000000000000000, /*   26 */
128'h00000000000000000000000000000000, /*   27 */
128'h00000000000000000000000000000000, /*   28 */
128'h00000000000000000000000000000000, /*   29 */
128'h00000000000000000000000000000000, /*   30 */
128'h00000000000000000000000000000000, /*   31 */
128'hd963454c0005cc635735c28587ae6914, /*   32 */
128'he21c97b6470102a787b30a00051300b7, /*   33 */
128'h853e85b200030563018533038082853a, /*   34 */
128'h908686930000c697b7edfda007138302, /*   35 */
128'h87930000c79762949d0707130000c717, /*   36 */
128'h87b30280069302d787bb878d8f999c67, /*   37 */
128'h47148082853a470100e7956397ba02d7, /*   38 */
128'hf0efe4061141b7f502870713fea68de3, /*   39 */
128'hbfe545018082014160a26108c509fbbf, /*   40 */
128'hf0efe852ec4ef04af426f822fc067139, /*   41 */
128'h0000ba17440144814985892acd31f9bf, /*   42 */
128'he091450100f44d6300c9278348ca0a13, /*   43 */
128'h61216a4269e2790274a2744270e25535, /*   44 */
128'h67a2ed19f29ff0ef854a85a200308082, /*   45 */
128'h50ef8552000995632485cb990087c783, /*   46 */
128'h0513bf652405274080ef498165224c40, /*   47 */
128'hf2dff0efe42ef406f0227179b7c1fda0, /*   48 */
128'h842aee7ff0ef083065a2c105fda00413, /*   49 */
128'h00f7096300c547030ff007936562e911, /*   50 */
128'h547980826145740270a2852223a080ef, /*   51 */
128'hf0efec4ef04af426f822fc067139bfd5, /*   52 */
128'h0000a9970ff00913440184aacd01eebf, /*   53 */
128'h74a2744270e200f4496344dc5a498993, /*   54 */
128'hf0ef852685a200308082612169e27902, /*   55 */
128'h85a20127896300c7c78367a2ed09e83f, /*   56 */
128'hb7d924051d4080ef6522420050ef854e, /*   57 */
128'he8dff0ef892eec26f406e84af0227179, /*   58 */
128'he45ff0ef84aa85ca0030c11dfda00413, /*   59 */
128'h548505130000a517864a608ced01842a, /*   60 */
128'h740270a28522196080ef65223e2050ef, /*   61 */
128'hf406ec26f022717980826145694264e2, /*   62 */
128'h85a6842ac11dfda00413e47ff0ef84ae, /*   63 */
128'hcf63445c3aa050ef520505130000a517, /*   64 */
128'h543515c080ef51e505130000a51700f4, /*   65 */
128'h003085228082614564e2740270a28522, /*   66 */
128'h130080ef6522f565842adcfff0ef85a6, /*   67 */
128'h5479fcf71be30ff0079300c7c70367a2, /*   68 */
128'he50965a2de1ff0eff406e42e7179bfc1, /*   69 */
128'hf96dd97ff0ef08308082614570a24501, /*   70 */
128'he42eec064108842ae8221101bfc56562, /*   71 */
128'h852200030e6302053303c919db9ff0ef, /*   72 */
128'h60e2fda005138302610560e265a26442, /*   73 */
128'h0000b7977139bfdd4501808261056442, /*   74 */
128'h04130000b417f426f822639c69478793, /*   75 */
128'h043b840d8c0574e484930000b4977564, /*   76 */
128'h892afc06e852ec4ef04a0280079302f4, /*   77 */
128'h942602f4043345ea0a130000aa1789ae, /*   78 */
128'h69e2790274a2744270e2450100849b63, /*   79 */
128'h2a6050ef855285ca6090808261216a42, /*   80 */
128'hbfc902848493c5016d3060ef854a608c, /*   81 */
128'hb7e16522f569cdbff0ef852685ce0030, /*   82 */
128'h84b68432e42efc06f04af426f8227139, /*   83 */
128'hcb5ff0ef083065a2c115cf7ff0ef893a, /*   84 */
128'h70e2978285a2615c862686ca6562e519, /*   85 */
128'hbfc5fda0051380826121790274a27442, /*   86 */
128'h84b68432e42efc06f04af426f8227139, /*   87 */
128'hc75ff0ef083065a2c115cb7ff0ef893a, /*   88 */
128'h70e2978285a2655c862686ca6562e519, /*   89 */
128'hbfc5fda0051380826121790274a27442, /*   90 */
128'hc7dff0ef84b2e42ef822fc06f4267139, /*   91 */
128'h701ce509c39ff0ef842a083065a2c105, /*   92 */
128'h8082612174a2744270e2978285a66562, /*   93 */
128'h2785c3190017f713419cbfcdfda00513, /*   94 */
128'hd71b8e5927a106220086571b419cc19c, /*   95 */
128'h0ff77713c19c0087d7138ed906a20086, /*   96 */
128'h122300d5112300c510238fd90087979b, /*   97 */
128'hf022f4067179419c80820005132300f5, /*   98 */
128'h419c00f510230457879b6785c19c27d1, /*   99 */
128'h0087979b0ff777130087d713c632842a, /*  100 */
128'hc4360509084c57fd460900f11a238fd9, /*  101 */
128'h05130161059346097bd060ef00f11b23, /*  102 */
128'h00041323082c462147c17af060ef0044, /*  103 */
128'h00f404a347c579b060efec3e00840513, /*  104 */
128'h785060ef00c4051300041523006c4611, /*  105 */
128'h01440693779060ef01040513002c4611, /*  106 */
128'hfed79ce39f31ffe7d6030789470187a2, /*  107 */
128'h9fb94107d71b9fb9934117424107579b, /*  108 */
128'h80826145740270a200f41523fff7c793, /*  109 */
128'h97b64721678563944b8787930000b797, /*  110 */
128'hc7bb27850077e793fff6079b8007bc23, /*  111 */
128'h678500f747630005071b6805450102e7, /*  112 */
128'h00e588b300351713808280c6b82396be, /*  113 */
128'hbfe1050501173023973697420008b883, /*  114 */
128'he406450185aa86220005841be0221141, /*  115 */
128'h717980820141640260a28522fa1ff0ef, /*  116 */
128'he436f4064619051984b2842aec26f022, /*  117 */
128'h6b5060ef85b64619852266a26c1060ef, /*  118 */
128'h00e4859b70a27402852200f4162347a1, /*  119 */
128'h6785737dc5010113fadff06f614564e2, /*  120 */
128'h38913c233a113423392138233a813023, /*  121 */
128'h3761382337513c233941302339313423, /*  122 */
128'h35a1382335913c233781302337713423, /*  123 */
128'hd00007b7943e747d978a911a35078793, /*  124 */
128'hf0040023e0040023ca040b23ce042023, /*  125 */
128'h00e7ea63892a5800073797aad0040023, /*  126 */
128'ha0017b9040ef15e505130000a51785aa, /*  127 */
128'h871374fd678524f71d63478900054703, /*  128 */
128'h970a350787139abacd848a93970a3507, /*  129 */
128'h49818a368cb28baed0048c13cb848b13, /*  130 */
128'hcd03013907b395ca0f0985939c3a9b3a, /*  131 */
128'h89bb058902a0071329890f07c7830015, /*  132 */
128'h22e78f63471904f76b6326e78b6301a9, /*  133 */
128'hcc848513470d2ae78963470502f76263, /*  134 */
128'h40ef262505130000a51785be22e78763, /*  135 */
128'hfee794e3473d22e783634731bf4d7350, /*  136 */
128'h953e866ae0048513978a350787936785, /*  137 */
128'h03600713b769e00d002357f060ef9d22, /*  138 */
128'h20e78e630330071300f76e6322e78163, /*  139 */
128'haac94605cb648513fae798e303500713, /*  140 */
128'hf8e79ce30ff0071324e7856303800713, /*  141 */
128'h8363479924f58363747d479500614583, /*  142 */
128'h16079263000ca7833af59f63478938f5, /*  143 */
128'h0593ce4405134985978a350a87936a85, /*  144 */
128'h8793507060ef013ca023953e46110109, /*  145 */
128'h953e461101490593ce840513978a350a, /*  146 */
128'h54e25a5203c505130000a5174f1060ef, /*  147 */
128'hcf840913978a350a8793671040efde02, /*  148 */
128'h03a3478d47b060ef854a55fd4619993e, /*  149 */
128'h978a350a879346f115231350079300f1, /*  150 */
128'h46c1051385a6460594becb740493c2a6, /*  151 */
128'h879346f106a30320079349f060efc0d2, /*  152 */
128'h051346114a1195becf040593978a350a, /*  153 */
128'h09a30360079347b060ef4741072346f1, /*  154 */
128'h461195becf440593978a350a879346f1, /*  155 */
128'h460557fd459060ef47410a2347510513, /*  156 */
128'h0d23000103a346f10ca347b1051385a6, /*  157 */
128'h45810f0006131020079343f060ef4731, /*  158 */
128'h1d23101007933dd060efde3e37a10513, /*  159 */
128'h36f10e233961051385de4799464136f1, /*  160 */
128'h679946f113232637879377e1411060ef, /*  161 */
128'h0413978a350a879346f1142335378793, /*  162 */
128'h051385a20440061304300693943ecec4, /*  163 */
128'h35e1051385a2460156fdba5ff0ef3721, /*  164 */
128'hcf3ff0ef0e8885de86ca5672bd9ff0ef, /*  165 */
128'h398134833a0134033a813083911a6305, /*  166 */
128'h37813a8338013a033881398339013903, /*  167 */
128'h35813c8336013c0336813b8337013b03, /*  168 */
128'h4611cd04851380823b01011335013d03, /*  169 */
128'h87936785a00d953e978a350787936785, /*  170 */
128'h60ef9d22953e866af0048513978a3507, /*  171 */
128'h355060ef85564611b3bdf00d00233630, /*  172 */
128'h978a350787936785bfdd855a4611b395, /*  173 */
128'hce045783339060ef4611953ece048513, /*  174 */
128'h578300f411238fd90087979b0087d71b, /*  175 */
128'h00f410238fd90087979b0087d71bce24, /*  176 */
128'h866ab749cc048513bb39cef42023401c, /*  177 */
128'h2783b321d00d00232fd060ef9d228562, /*  178 */
128'h0000a51700fa2023478512079a63000a, /*  179 */
128'h0e8801090593461146f040efe4c50513, /*  180 */
128'hcb840513978a3504879364852d1060ef, /*  181 */
128'h353147032b9060ef014905934611953e, /*  182 */
128'h0000a517350145833511460335214683, /*  183 */
128'h00a146833501578342f040efe1c50513, /*  184 */
128'h352157831cf71e230000b71700914603, /*  185 */
128'h0000b717e1c505130000a51700814583, /*  186 */
128'h01b147033fb040ef00b147031cf71323, /*  187 */
128'h0000a517018145830191460301a14683, /*  188 */
128'h01214683013147033df040efe1c50513, /*  189 */
128'he20505130000a5170101458301114603, /*  190 */
128'h05130000a51755c2010157833c3040ef, /*  191 */
128'hb7170121578316f713230000b717e2e5, /*  192 */
128'hf6bb02f5d63b03c0079314f71e230000, /*  193 */
128'h02f5d5bbe107879b678502f6763b02f5, /*  194 */
128'h95bee0040593978a35048793383040ef, /*  195 */
128'h3504879336b040efe08505130000a517, /*  196 */
128'he00505130000a51795be978af0040593, /*  197 */
128'h40efe0a505130000a517bbf5353040ef, /*  198 */
128'h20234785de0794e3000a2783b3fd3450, /*  199 */
128'ha517329040efdfe505130000a51700fa, /*  200 */
128'h35078793678531d040efe02505130000, /*  201 */
128'he08505130000a51795be978ad0040593, /*  202 */
128'hb34d2f9040efe0e505130000a517bf45, /*  203 */
128'hf852fc4ee0cae4a6e8a2ec86711d737d, /*  204 */
128'h6a85e22505130000a517911a89aaf456, /*  205 */
128'h0493978a020a8793747d2d1040efca02, /*  206 */
128'hb7970d9060ef852655fd461994beff84, /*  207 */
128'hc83e4a05fef40913439ce82787930000, /*  208 */
128'h993e978a020a879312f11d2313500793, /*  209 */
128'h07930f7060ef014107a31a68460585ca, /*  210 */
128'h020a879312f10f23479112f10ea30370, /*  211 */
128'h60ef13f10513461195beff040593978a, /*  212 */
128'h14f101a314510513460585ca57fd0d30, /*  213 */
128'h0fc007930b9060ef000107a315410223, /*  214 */
128'h057060efca3e04a1051345810f000613, /*  215 */
128'h05134641479985ce04f1152310100793, /*  216 */
128'h2637879377e108b060ef04f106230661, /*  217 */
128'h879312f11c2335378793679912f11b23, /*  218 */
128'h06930421051385a2943e1451978a020a, /*  219 */
128'h02e1051385a2821ff0ef044006130430, /*  220 */
128'h85ce86a610084652855ff0ef460156fd, /*  221 */
128'h64a66446450160e6911a630596fff0ef, /*  222 */
128'ha51785aa808261257aa27a4279e26906, /*  223 */
128'hf0a2f48671591ad0406fd12505130000, /*  224 */
128'h05a1051384aa81010113e4cee8caeca6, /*  225 */
128'h60efd602e83eec3ae442893689b2e046, /*  226 */
128'h6762747d97ba81078793101867857f20, /*  227 */
128'h0521051385a2864a86ba943e7fc40413, /*  228 */
128'h863e86c285a267c26822f94ff0efd64e, /*  229 */
128'h85a6180856326882fc4ff0ef03e10513, /*  230 */
128'h7406450170a67f0101138ddff0ef86c6, /*  231 */
128'he222e606716d8082616569a6694664e6, /*  232 */
128'h00254703003547830045480300554883, /*  233 */
128'h85930000a597842a0005460300154683, /*  234 */
128'h85220f9040efc76505130000a517c765, /*  235 */
128'h85930000a597860ac10d842ae01ff0ef, /*  236 */
128'h85220d9040efc7e505130000a517c565, /*  237 */
128'hc98505130000a51780826151641260b2, /*  238 */
128'h7159b7cd0bb040efe007a8230000b797, /*  239 */
128'hec66f062f45ef85afc56e0d2e4ceeca6, /*  240 */
128'h44818aae89aae46ee8caf0a2f486e86a, /*  241 */
128'hc70b0b130000ab17940a0a130000ba17, /*  242 */
128'h0000ac97c7cc0c130000ac1706000b93, /*  243 */
128'h035441630004841bfff58d1bc6cc8c93, /*  244 */
128'h7b427ae26a0669a6694664e6740670a6, /*  245 */
128'hc01d808261656da26d426ce27c027ba2, /*  246 */
128'hff04891303b040ef855ae39d00f47793, /*  247 */
128'h7b0505130000a51702879d630009079b, /*  248 */
128'hc583009987b301d040ef8552023040ef, /*  249 */
128'h1263009040efc16505130000a5170007, /*  250 */
128'h87b3a80500f979134d81fffd4913068d, /*  251 */
128'he7630ff7f793fe05879b0007c5830129, /*  252 */
128'h40ef8562b75d09057de040ef856600fb, /*  253 */
128'hff2dcce32d857cc040ef8552bfdd7d40, /*  254 */
128'h079b4124093b7bc040ef00f4f913855a, /*  255 */
128'h40ef732505130000a51700f45a630009, /*  256 */
128'h879b0007c583012987b3bf1504857a40, /*  257 */
128'h786040ef856600fbe7630ff7f793fe05, /*  258 */
128'hec267179bfdd77c040ef8562b7f10905, /*  259 */
128'ha697893289ae84b6f022f406e44ee84a, /*  260 */
128'hb68686930000a697c5093ba686930000, /*  261 */
128'hb60606130000a6170187071300009717, /*  262 */
128'h5d6300098f63842a6fe040ef854a85a6, /*  263 */
128'hb48606130000a61786ce40a485bb0095, /*  264 */
128'h00f44463ffe4879b9c296e0040ef954a, /*  265 */
128'hb18585930000a59700890533ffd4841b, /*  266 */
128'h69a2694264e2854a740270a22bc060ef, /*  267 */
128'h7115f73ff06f4581862e86b280826145, /*  268 */
128'h002cfebff0efed8645050c800613002c, /*  269 */
128'h450160ee6ca040efb00505130000a517, /*  270 */
128'h6963862e9ff787133b9ad7b78082612d, /*  271 */
128'h079304a7676323f78713000f47b704a7, /*  272 */
128'h0000b7173e80079346890ca7fc633e70, /*  273 */
128'hec0600074903e04a97361101a7470713, /*  274 */
128'h690264a260e2644202091663e426e822, /*  275 */
128'h6660406f6105aa6505130000a51785aa, /*  276 */
128'hbf7d240787934685b7d9a00787934681, /*  277 */
128'h47293e800793c81502f555b302f57433, /*  278 */
128'h0713cf3902f4773346a547a90687e263, /*  279 */
128'h743302f457b30640071300877d630630, /*  280 */
128'h0000a517943e001444130324341302e4, /*  281 */
128'ha51785a2c80160c040ef84b2a5c50513, /*  282 */
128'h862660e264425fc040efa52505130000, /*  283 */
128'h6105a42505130000a517690264a285ca, /*  284 */
128'hf46302f45733bf6102e454335e20406f, /*  285 */
128'h0000a51785aabf554401bf51843a0086, /*  286 */
128'h86bb459958d94701862ebfa19fc50513, /*  287 */
128'h1702cf8500f557b3883e03c6879b02e8, /*  288 */
128'he426972e1101976585930000b5979301, /*  289 */
128'h60e26442e495e04ae822ec0600074483, /*  290 */
128'h61059da505130000a51785aa690264a2, /*  291 */
128'h0000a51785aafab71ce327055720406f, /*  292 */
128'hfff7471301071733577db7f59c450513, /*  293 */
128'h03b6869b02e505334729c10d44018d79, /*  294 */
128'h746301045433942a472500d414334405, /*  295 */
128'h970505130000a51785be078514590087, /*  296 */
128'h05130000a51785a2c801520040ef8932, /*  297 */
128'h690285a6864a60e26442510040ef9665, /*  298 */
128'h4f60406f610596e505130000a51764a2, /*  299 */
128'hf54ef94ae1a202c7073b8cbafce67155, /*  300 */
128'he162e55ee95aed56f152fd26e586f8ea, /*  301 */
128'hf66384368d3289ae892a04000793f4ee, /*  302 */
128'h4cc1000c956302ccdcbb04000c9300e7, /*  303 */
128'h001a849b020d1a13001d1a9b03acdcbb, /*  304 */
128'h0000ab9791cb0b130000ab17020a5a13, /*  305 */
128'h4501e00d7dcc0c1300008c17884b8b93, /*  306 */
128'h6b4a6aea7a0a79aa794a74ea640e60ae, /*  307 */
128'h85ca808261697da67d467ce66c0a6baa, /*  308 */
128'h00040d9b45a040ef8d8505130000a517, /*  309 */
128'h482146914781874e000c8d9b008cf463, /*  310 */
128'h9381020d979305b66b630007861b4889, /*  311 */
128'h083803bd06bb0d9de56399be034787b3, /*  312 */
128'h0b079c630006881b02e0089385ba4781, /*  313 */
128'h8c23e036894505130000a51797ba1098, /*  314 */
128'h9281168241b4043b6682400040effa07, /*  315 */
128'h02dd1963b79d557dd13d10a070ef9936, /*  316 */
128'h1602c19095aa26010828002795934310, /*  317 */
128'h67023c8040efe03ae43e855a85d69201, /*  318 */
128'h1963bf9d4691482107859752488967a2, /*  319 */
128'hbfd1e19095aa0828003795936310010d, /*  320 */
128'h164208280017959300075603011d1d63, /*  321 */
128'h082c00074603bf6d00c5902395aa9241, /*  322 */
128'he03e855eb76500c580230ff6761395be, /*  323 */
128'hbf253cfdfe97eae327856782136070ef, /*  324 */
128'h0005450300cc053300074603bfdd4781, /*  325 */
128'h54634186561b0186161bc51909757513, /*  326 */
128'h87aa1582b70d07052785011700230006, /*  327 */
128'h8f8d25058082e21c00b7f46345019181, /*  328 */
128'h0088458189aa04000613fd4e7115bfd5, /*  329 */
128'hed5ef15af556f952e1cae5a6e9a2ed86, /*  330 */
128'h07130000a71767869982e16ae566e962, /*  331 */
128'h440106e79d63557983e107e2631868e7, /*  332 */
128'h9b9776ab0b1300009b174a8503800a13, /*  333 */
128'h9d1708000cb780000c377a2b8b930000, /*  334 */
128'h656600f464630781578377ad0d130000, /*  335 */
128'h9dbd0028038006137786028a05bba091, /*  336 */
128'h855a85a2cfbd77c20957926347a29982, /*  337 */
128'h018487b37482040908637922292040ef, /*  338 */
128'h40ef71a505130000951785a60397e863, /*  339 */
128'h7a4a79ea690e64ae644e60ee55752740, /*  340 */
128'h8082612d6d0a6caa6c4a6bea7b0a7aaa, /*  341 */
128'h061b45c224a040ef856a86ca85a66642, /*  342 */
128'h79020097ff6377a274c2998285260009, /*  343 */
128'h8626228040ef855e85ca993e86268c9d, /*  344 */
128'h057e4505bfb1240503e060ef854a4581, /*  345 */
128'h780707130000a7178082400005378082, /*  346 */
128'he30895360017869300756513157d631c, /*  347 */
128'h67858082953e057e450597aa20000537, /*  348 */
128'h871308a74463862a0ce5076382078713, /*  349 */
128'h496306e60b636c650513000095178087, /*  350 */
128'hc3ad6a250513000095178006079b04c7, /*  351 */
128'hc963722505130000951787f787936785, /*  352 */
128'h000095979e3d11417c07879b77fd04c7, /*  353 */
128'h40efe4066e4505130000a51771458593, /*  354 */
128'h808201416d4505130000a51760a21600, /*  355 */
128'h00e60a63674505130000951781078713, /*  356 */
128'hfaf612e3674505130000951781878793, /*  357 */
128'h09e36925051300009517830787138082, /*  358 */
128'h0513000095178287879300c74963fee6, /*  359 */
128'h680505130000951783878713bfe966e5, /*  360 */
128'h680505130000951784078793fce608e3, /*  361 */
128'hf022717980826365051300009517bf75, /*  362 */
128'h07bb00a5893b440184aaf406e84aec26, /*  363 */
128'h942a904114420104551302f044634099, /*  364 */
128'h1542fff54513740270a2952201045513, /*  365 */
128'h0068460985a6808261459141694264e2, /*  366 */
128'h979b0087d71b048900c15783731050ef, /*  367 */
128'hbf45943e93c117c200f117238fd90087, /*  368 */
128'h8793f44ef84afc26e486e0a26785715d, /*  369 */
128'h0e636dd7879367a13cf50463842e8067, /*  370 */
128'h082884b205e9440799638005079b0af5, /*  371 */
128'ha517461985ca006409136df050ef4611, /*  372 */
128'h0793017445836cb050ef5d2505130000, /*  373 */
128'h1cf5816347b108b7e76332f5886302e0, /*  374 */
128'h478502b7e3631af58263479104b7e563, /*  375 */
128'h83635ba5051300009517478910f58463, /*  376 */
128'ha415018040ef756505130000951702f5, /*  377 */
128'h5c0505130000951747a118f581634799, /*  378 */
128'h2cf5816347f5a4297ff030effef591e3, /*  379 */
128'h0000951747d916f5896347c500b7ed63, /*  380 */
128'h856302100793bf6dfef580e35dc50513, /*  381 */
128'h051300009517faf596e3029007932af5, /*  382 */
128'h04b7e2632cf5816306200793b7c95f65, /*  383 */
128'h02f0079300b7ef632af5816303300793, /*  384 */
128'h5f850513000095170320079328f58663, /*  385 */
128'h079328f5836305c00793b7bdf8f58ae3, /*  386 */
128'hbf91f6f58de360e505130000951705e0, /*  387 */
128'h0670079300b7ef6328f5856308400793, /*  388 */
128'h620505130000951706c0079326f58a63, /*  389 */
128'h079326f5876308900793b73df4f58ae3, /*  390 */
128'h9517f0f59ce30880079326f588630ff0, /*  391 */
128'h0000a79701e45703b73d62a505130000, /*  392 */
128'h12f713634dc989930000a9974e47d783, /*  393 */
128'h10f71b634ce7d7830000a79702045703, /*  394 */
128'h0000a597461956b050ef852285ca4619, /*  395 */
128'h012301a4578355b050ef854a49c58593, /*  396 */
128'h859b01c4578300f41f23020412230204, /*  397 */
128'h1d230009d78302f4102302240513fde4, /*  398 */
128'h579bdb3ff0ef00f41e230029d78300f4, /*  399 */
128'h862602a4122300a11e238d5d05220085, /*  400 */
128'h051300009517a06ddcdfe0ef450185a2, /*  401 */
128'h9517b56143c5051300009517bd4942e5, /*  402 */
128'h0264470302444783bdbd44a505130000, /*  403 */
128'h01c1178300f10e230254478300f10ea3, /*  404 */
128'h470300e10e2327810274470300e10ea3, /*  405 */
128'h0e230234470300e10ea301c119030224, /*  406 */
128'ha79704e79b6301c156830450071300e1, /*  407 */
128'h85930000a597461947e23ad79f230000, /*  408 */
128'h2f230000a71739e505130000a5173965, /*  409 */
128'h0000a79766a2476247d050efe43638f7, /*  410 */
128'h60ef450102a40593ff89061b37478793, /*  411 */
128'h8082616179a2794274e2640660a65a00, /*  412 */
128'h2f230000a71747e204e6946304300713, /*  413 */
128'ha797c799439c362787930000a79734f7, /*  414 */
128'h86930000a697f7e9439c352787930000, /*  415 */
128'h85930000a597342606130000a6173466, /*  416 */
128'h4d200713b765d73fe0ef02a405133465, /*  417 */
128'h587030ef364505130000951702e79863, /*  418 */
128'h3605051300009517ccaff0ef852285a6, /*  419 */
128'hbf95cb4ff0ef02a4051385ca573030ef, /*  420 */
128'h17fd67c101e45703f6e787e35fe00713, /*  421 */
128'ha5974611f4f70de302045703f6f701e3, /*  422 */
128'h9517b7993a9050ef0868302585930000, /*  423 */
128'h3405051300009517b33d33a505130000, /*  424 */
128'h00009517bb293565051300009517b315, /*  425 */
128'hb31937a5051300009517bb0136450513, /*  426 */
128'h051300009517b9f53805051300009517, /*  427 */
128'h9517b1e53ac5051300009517b9cd39e5, /*  428 */
128'h3e85051300009517b9f93c2505130000, /*  429 */
128'h0265d703b1e93f65051300009517b9d1, /*  430 */
128'h278484930000a4972807d7830000a797, /*  431 */
128'h26a7d7830000a7970285d703ecf711e3, /*  432 */
128'h016589930205891320000793eaf719e3, /*  433 */
128'h46192f7050ef854a85ce461900f59a23, /*  434 */
128'h46192e7050ef854e228585930000a597, /*  435 */
128'h2d5050ef00640513218585930000a597, /*  436 */
128'h061301c457832cb050ef852285ca4619, /*  437 */
128'hd78302f4142301e4578302f4132302a0, /*  438 */
128'h079300f41f230024d78300f41e230004, /*  439 */
128'h05130000951785aab36900f416236080, /*  440 */
128'hb603430017b7bba54601421030ef37e5, /*  441 */
128'h00f674132601608130239f0101138307, /*  442 */
128'h879b0387f5930034179b66858387b703, /*  443 */
128'h5e913c23639c97ae430005b79fad8406, /*  444 */
128'h849b5f200513fee7881b278160113423, /*  445 */
128'h00c5163b101005138a1d09056c63ffc7, /*  446 */
128'h07130000a717c34927018f71fff74713, /*  447 */
128'h871b700776130084171beb3d431814e7, /*  448 */
128'h969b00d100a345d495ba070e9f318006, /*  449 */
128'h550300d100230086d69b0106d69b0106, /*  450 */
128'h1e63806686936685c6918005069b0001, /*  451 */
128'h43000837860a27850077e79337ed02d5, /*  452 */
128'h983a00369813974285b246814037d79b, /*  453 */
128'h0006881bff063c230621068500083803, /*  454 */
128'h430017b70405a9bff0ef8626fef845e3, /*  455 */
128'h3483852660013403608130838287b823, /*  456 */
128'he8220c2007b711018082610101135f81, /*  457 */
128'hb703430014b747812401ec06e42643c0, /*  458 */
128'h00009517e7990206c163033716938304, /*  459 */
128'h60e2c3c00c2007b72ef030ef26450513, /*  460 */
128'hbfc14785ec3ff0ef8082610564a26442, /*  461 */
128'h0000a597461184ae8432ec26f0227179, /*  462 */
128'h0000a797129050eff406006808458593, /*  463 */
128'ha89785a6862247b20007a80303c78793, /*  464 */
128'h0693026757030000a717022888930000, /*  465 */
128'h85228e0ff0ef02e505130000a5170450, /*  466 */
128'h05220085579b8082614564e2740270a2, /*  467 */
128'h0185579b0185171b8082914115428d5d, /*  468 */
128'h8fd98f750085571bf00686938fd966c1, /*  469 */
128'h808225018d5d8d7900ff07370085151b, /*  470 */
128'h4585460100740207879b070007b7715d, /*  471 */
128'hf44ef84ae0a2fc26e486c63e04b00513, /*  472 */
128'h05130000951784aa099070efec56f052, /*  473 */
128'hc31101079713fff4c793211030ef19e5, /*  474 */
128'ha7175785f8f70e230000a71757b9ecc5, /*  475 */
128'hf8f705230000a7175789f8f709a30000, /*  476 */
128'h0000a7175791f8f700a30000a717578d, /*  477 */
128'ha797fe056513893d027070eff6f70c23, /*  478 */
128'hf5a585930000a5974611f6a783a30000, /*  479 */
128'hf48585930000a597460901f050ef0048, /*  480 */
128'h06374722f31ff0ef451200f050ef0028, /*  481 */
128'h77138ff183210087179bf00606130100, /*  482 */
128'hb02317c29101430016b78fd915020ff7, /*  483 */
128'h8086b7838006b78380f6b42393c180a6, /*  484 */
128'h79a2794274e282f6b42347a1640660a6, /*  485 */
128'h0000aa175ae14401808261616ae27a02, /*  486 */
128'h863b49190d49899300009997ee4a0a13, /*  487 */
128'h061b0405854e0004059b014407b3028a, /*  488 */
128'h30ef00c780230ff6761300c4d6330286, /*  489 */
128'h8007b603430017b7bf81fd241ee31150, /*  490 */
128'h8f4d91c115c20080073771398087b583, /*  491 */
128'he05ae456e852ec4ef04af426f822fc06, /*  492 */
128'h0d7030ef08c505130000951780e7b423, /*  493 */
128'he6c7c7830000a797e73747030000a717, /*  494 */
128'he5a6c6830000a697e65848030000a817, /*  495 */
128'he485c5830000a597e51646030000a617, /*  496 */
128'h0000a41709b030ef0605051300009517, /*  497 */
128'h89930000a997448100044783e3440413, /*  498 */
128'haa1700144783e2f703230000a717e0e9, /*  499 */
128'he0f708a30000a7176a89e02a0a130000, /*  500 */
128'h0000a7174300193700262b3700244783, /*  501 */
128'hdef709a30000a71700344783def70f23, /*  502 */
128'h00544783def704230000a71700444783, /*  503 */
128'hda079a230000a797dcf70ea30000a717, /*  504 */
128'hda07a8230000a797da07a4230000a797, /*  505 */
128'hd807ac230000a797da07a2230000a797, /*  506 */
128'h0493ed1fe0ef8522e78d0009a783e4a9, /*  507 */
128'h37830207456303379713830937835a0b, /*  508 */
128'hbfc5bc1ff0effc075de3033797138309, /*  509 */
128'h84937c9050ef4501dff154fd000a2783, /*  510 */
128'h4783b7d914fdb7e9ba7ff0efbfc1710a, /*  511 */
128'h4503002547838f5d07a2000547030015, /*  512 */
128'h4781808225018d5d05628fd907c20035, /*  513 */
128'h468300f58733808200e613630007871b, /*  514 */
128'h9e29b7d500d70023078500f507330007, /*  515 */
128'hfeb50fa30505808200f613630005079b, /*  516 */
128'h8413e04ae426ec06e8221101495cbfc5, /*  517 */
128'h451502000613478101853903cfb50095, /*  518 */
128'h0007470300f9073346ad02e008934821, /*  519 */
128'h0007831b0e50071300a7146302c70063, /*  520 */
128'h040500e4002304050114002301031563, /*  521 */
128'h84ae01c9051300b94783fcd79be30785, /*  522 */
128'h470301994783c088f4bff0ef00f58423, /*  523 */
128'h0179478300f492238fd90087979b0189, /*  524 */
128'h002300f493238fd90087979b01694703, /*  525 */
128'h611c80826105690264a2644260e20004, /*  526 */
128'h0007468303a0061302000593cf99873e, /*  527 */
128'h00d706630017869300c6986302d5fc63, /*  528 */
128'h577d46050007c683b7dd0705a00d577d, /*  529 */
128'h871b078900b666630ff6f593fd06869b, /*  530 */
128'hc50747030000a7178082853ae11c0006, /*  531 */
128'hd683c70d0007c703cb85611cc915bfd5, /*  532 */
128'hc503e406114102e69063008557030067, /*  533 */
128'h4525c391450100157793402060ef0017, /*  534 */
128'hc68301b5c783808245258082014160a2, /*  535 */
128'h1d630006879b8edd0087979b470d01a5, /*  536 */
128'h8fd10087179b0145c6030155c70300e5, /*  537 */
128'hf02271798082853e27818fd50107979b, /*  538 */
128'h03450993e052e84af4065904e44eec26, /*  539 */
128'h390060ef85ce8626468500154503842a, /*  540 */
128'h40f487bb000402234c58505ce1312501, /*  541 */
128'h69a2694264e2740270a2450100e7eb63, /*  542 */
128'hff2a74e34a0500344903808261456a02, /*  543 */
128'h60ef85ce86269cbd4685001445034c5c, /*  544 */
128'hc39900454783b7f94505b7e5397d34e0, /*  545 */
128'hec06e8221101591c80824501f8dff06f, /*  546 */
128'hf0ef892e84aa02b787634401e04ae426, /*  547 */
128'h864a46850014c503ec190005041bfddf, /*  548 */
128'h597d4405c11925012d6060ef03448593, /*  549 */
128'h6105690264a2644260e285220324a823, /*  550 */
128'h022357fde04ae426ec06e82211018082, /*  551 */
128'h4783e52d2501fa3ff0ef842ad91c0005, /*  552 */
128'h979b8fd90087979b4509232447032334, /*  553 */
128'h02e79f63a55707134107d79b776d0107, /*  554 */
128'h010005370005079bd4bff0ef06a40513, /*  555 */
128'h0127f7b31465049300544537fff50913, /*  556 */
128'h2501d25ff0ef0864051300978c634501, /*  557 */
128'h64a2644260e200a035338d0501257533, /*  558 */
128'hf44ef84a715dbfcd450d808261056902, /*  559 */
128'h89aa00053023ec56f052fc26e0a2e486, /*  560 */
128'h171302054e6347adddbff0ef8932852e, /*  561 */
128'h84aa638097baa56787930000a7970035, /*  562 */
128'h4503c79d000447830089b023c01547b1, /*  563 */
128'h00090563e38500157793222060ef0014, /*  564 */
128'h79a2794274e2640660a647a9c1118911, /*  565 */
128'h00230ff4f51380826161853e6ae27a02, /*  566 */
128'h478d00157713136060ef00a400a30004, /*  567 */
128'hf0ef85224581f571891100090463fb79, /*  568 */
128'h0a131fa40913848a04f51a634785ee5f, /*  569 */
128'hf0ef854ac7894501ffc9478389a623a4, /*  570 */
128'hff2a14e30991094100a9a0232501c51f, /*  571 */
128'h85d2000a076345090004aa0301048913, /*  572 */
128'h470dfe9915e30491c10dea1ff0ef8522, /*  573 */
128'hf6e505e34785470dbf8500e519634785, /*  574 */
128'h03f4470304044783b78547b5c1194a01, /*  575 */
128'h07134107d79b0107979b8fd90087979b, /*  576 */
128'h999b04a4478304b44983fee791e32000, /*  577 */
128'h0444448329811a09876300f9e9b30089, /*  578 */
128'hf793009401a3fff4879b470501342e23, /*  579 */
128'h03e30124012304144903faf769e30ff7, /*  580 */
128'h4a83ffc100f977b3fff9079b2901fa09, /*  581 */
128'h142300faeab3008a9a9b045447830464, /*  582 */
128'h0474478304844503ffbd00faf7930154, /*  583 */
128'h47030434478314050e638d5d0085151b, /*  584 */
128'h033486bbdfa98fd90087979b25010424, /*  585 */
128'h63e3873200d7063b9f3d004ad71b2781, /*  586 */
128'hf3266ce384ae032655bb40c5063bf4c5, /*  587 */
128'h39331955694100b67763490516556605, /*  588 */
128'hd458014787bb24890147073b090900b9, /*  589 */
128'h93e310e91163470dd05c03442023cc04, /*  590 */
128'h0024949bd408b09ff0ef06040513f00a, /*  591 */
128'hc81c57fdee99e6e30094d49b1ff4849b, /*  592 */
128'h08f91963478d00f402a3f8000793c45c, /*  593 */
128'h979b8fd90087979b0644470306544783, /*  594 */
128'h001a059b06e79b6347054107d79b0107, /*  595 */
128'h470323344783e13d2501ce7ff0ef8522, /*  596 */
128'h0107979b8fd90087979b000402a32324, /*  597 */
128'h051304e79263a55707134107d79b776d, /*  598 */
128'h252787932501416157b7a8dff0ef0344, /*  599 */
128'h614177b7a77ff0ef2184051302f51763, /*  600 */
128'hf0ef21c4051300f51c63272787932501, /*  601 */
128'h9797c448a57ff0ef22040513c808a61f, /*  602 */
128'h0000971793c117c227857dc7d7830000, /*  603 */
128'h00042a230124002300f413237cf71723, /*  604 */
128'h0005099ba27ff0ef05840513b3514781, /*  605 */
128'he00a84e3b545a19ff0ef05440513b5b1, /*  606 */
128'hb7090014949b00f915634789d41c9fb5, /*  607 */
128'hbdcd9cbd0017d79b8885029787bb478d, /*  608 */
128'h2501c01ff0ef842ae426ec06e8221101, /*  609 */
128'h005447030cf71063478d00044703ed69, /*  610 */
128'h458120000613034404930af71b634785, /*  611 */
128'h079322f40923055007939fdff0ef8526, /*  612 */
128'h0aa302f40a230520079322f409a3faa0, /*  613 */
128'h481c20f40da302f40b230610079302f4, /*  614 */
128'h0107971b20e40d2302e40ba304100713, /*  615 */
128'h20e40ea320f40e230087571b0107571b, /*  616 */
128'h0f23445c20f40fa30187d79b0107d71b, /*  617 */
128'h0087571b0107571b0107971b501020e4, /*  618 */
128'h22e400a322f400230720069300144503, /*  619 */
128'h0ca320d40c230187d79b0107d71b2605, /*  620 */
128'h85a64685d81022f401a322e4012320d4, /*  621 */
128'h4581460100144503000402a367d050ef, /*  622 */
128'h64a2644260e200a035332501671050ef, /*  623 */
128'hf963377985beffe5879b4d1880826105, /*  624 */
128'h80829d3d02b787bb55480025478300e7, /*  625 */
128'he84a71794d180eb7f563478580824501, /*  626 */
128'h470302e5f963892ae44eec26f022f406, /*  627 */
128'h08d70d63468d06d70b63842e46890005, /*  628 */
128'h0094d59b9cad515c0015d49b00f71e63, /*  629 */
128'h740270a257fdc9112501ac7ff0ef9dbd, /*  630 */
128'h0249278380826145853e69a2694264e2, /*  631 */
128'h9dbd94ca1ff4f4930099d59b0014899b, /*  632 */
128'hf993f5792501a93ff0ef0344c483854a, /*  633 */
128'h8fc50087979b880503494783994e1ff9, /*  634 */
128'hd59b515cbf4d93d117d2bf658391c019, /*  635 */
128'h0014141bf1452501a65ff0ef9dbd0085, /*  636 */
128'h979b034945030359478399221fe47413, /*  637 */
128'hf0ef9dbd0075d59b515cb7618fc90087, /*  638 */
128'h05131fc575130024151bf93d2501a3bf, /*  639 */
128'hbfb9024557931512ffaff0ef954a0345, /*  640 */
128'hfc06f04a4544f42671398082853e4785, /*  641 */
128'h892a478500b51523e456e852ec4ef822, /*  642 */
128'h69e2790274a2744270e2450900f49c63, /*  643 */
128'hfee4f4e34f98611c808261216aa26a42, /*  644 */
128'h579800e69463470d0007c683e0a9842e, /*  645 */
128'h009928235788fce477e30087d703eb0d, /*  646 */
128'h0009378300f92a239fa90044579bd171, /*  647 */
128'h450100893c23943e034787930416883d, /*  648 */
128'h350309924a855a7d0027c98384bab75d, /*  649 */
128'hbf7d2501e5dff0ef0134766385a60009, /*  650 */
128'hf69afce301448c630005049be75ff0ef, /*  651 */
128'hbfc14134043bf6f4f7e34f9c00093783, /*  652 */
128'hec06e426e822110100a55583b7954505, /*  653 */
128'h6008484ce4950005049bf35ff0ef842a, /*  654 */
128'h020006136c08ec990005049b939ff0ef, /*  655 */
128'h601c00e7802357156c1cf3cff0ef4581, /*  656 */
128'h610564a28526644260e200e782234705, /*  657 */
128'hf04af426f822fc06e852ec4e71398082, /*  658 */
128'h4a0984aa4d1c0ab9f5634a094985e456, /*  659 */
128'h8f63842e89324709000547830af5f063, /*  660 */
128'h0015d99b093794630ee78863470d0ae7, /*  661 */
128'h8bdff0ef9dbd0099d59b00b989bb515c, /*  662 */
128'h779300198a9b8805060a166300050a1b, /*  663 */
128'h0347c783013487b3cc191ff9f9930ff9, /*  664 */
128'h8fd98ff50049179b00f7f71316c16685, /*  665 */
128'h00f48223478502f98a2399a60ff7f793, /*  666 */
128'h0a1b86fff0ef9dbd8526009ad59b50dc, /*  667 */
128'h0049591bc40d1ffafa93000a1f630005, /*  668 */
128'h00f482234785032a8a239aa60ff97913, /*  669 */
128'h6aa26a4269e2790274a28552744270e2, /*  670 */
128'h0089591b0347c783015487b380826121, /*  671 */
128'hd59b515cb7e90127e9339bc100f97913, /*  672 */
128'hfc0a12e300050a1b815ff0ef9dbd0085, /*  673 */
128'h191b03240a2394261fe474130014141b, /*  674 */
128'h822303240aa30089591b0109591b0109, /*  675 */
128'hfdcff0ef9dbd0075d59b515cbf790134, /*  676 */
128'h1fc474130024141bf80a16e300050a1b, /*  677 */
128'h06372501d96ff0ef85569aa603440a93, /*  678 */
128'h94260109179b2901012569338d71f000, /*  679 */
128'h00fa80a30087d79b03240a230107d79b, /*  680 */
128'h012a81a300fa81230189591b0109579b, /*  681 */
128'he852f04af822fc06ec4ef4267139bf79, /*  682 */
128'h0009056300c52903e99189ae84aae456, /*  683 */
128'h041bc5bff0efa815490502f96d634d1c, /*  684 */
128'h744270e2852244050087ed6347850005, /*  685 */
128'h57fd808261216aa26a4269e2790274a2, /*  686 */
128'h4a05844afef461e3894e4c9c08f40263, /*  687 */
128'h4401012a646300f4676324054c9c5afd, /*  688 */
128'hc9012501c0dff0ef852685a24409b7e9, /*  689 */
128'h0637b7cdfd241de3fb450ae305550a63, /*  690 */
128'he9052501debff0ef852685a2167d1000, /*  691 */
128'h37fdf8e788e3577dc4c0489c02099063, /*  692 */
128'hbfb500f482a30017e7930054c783c89c, /*  693 */
128'h4785dd612501dbdff0ef852685ce8622, /*  694 */
128'h00a55903f04a7139b795547df6f514e3, /*  695 */
128'he852ec4ef426030917932905f822fc06, /*  696 */
128'h790274a2744270e24511eb9993c1e456, /*  697 */
128'h7993d7ed495c808261216aa26a4269e2, /*  698 */
128'h61082785480c00099d63842a8a2e00f9, /*  699 */
128'hfcf775e30009071b00855783e18dc85c, /*  700 */
128'hec1c97ce03478793012415230996601c, /*  701 */
128'hfab337fd00495a9b00254783bf5d4501, /*  702 */
128'h47850005049bb2fff0effc0a9fe30157, /*  703 */
128'h450500f4946357fdbf4945090097e463, /*  704 */
128'h480cf60a0ee306f4e0634d1c6008b761, /*  705 */
128'h8be34785d4bd451d0005049be83ff0ef, /*  706 */
128'h2501de0ff0ef6008fcf48de357fdfcf4, /*  707 */
128'hf0ef034505134581200006136008f579, /*  708 */
128'h2823aabff0ef855285a600043a03bf0f, /*  709 */
128'h591c00faed630025478360084a0502aa, /*  710 */
128'ha89ff0ef85a6c8046008d91c415787bb, /*  711 */
128'hf1412501d24ff0ef01450223b7b9c848, /*  712 */
128'hf8227139b7e9db1c27855b1c2a856018, /*  713 */
128'hc783e05ae456e852ec4ef04afc06f426, /*  714 */
128'h071300e78663842e84aa02f007130005, /*  715 */
128'h000447030004a62304050ce7946305c0, /*  716 */
128'h099305c00a9302f00a130ce7f06347fd, /*  717 */
128'h0d5784630d478663000447834b2102e0, /*  718 */
128'hb42ff0ef854a02000593462d0204b903, /*  719 */
128'h00144783013900230d37966300044783, /*  720 */
128'h0024478300f900a302e007930b379463, /*  721 */
128'h02000793943a09479b63470d1d378963, /*  722 */
128'h19632501adfff0ef8526458100f905a3, /*  723 */
128'h11632501ce0ff0ef608848cc492d1005, /*  724 */
128'h00b7478312078063000747836c981005, /*  725 */
128'h00f58633078500f706b3708cef898ba1, /*  726 */
128'h852645810cd60a63fff646030006c683, /*  727 */
128'hc55c4bdc611ca0e1dd5d2501df9ff0ef, /*  728 */
128'h0004bc232501a81ff0ef85264581bf35, /*  729 */
128'h6b026aa26a4269e2790274a2744270e2, /*  730 */
128'hf75787e3b7b54709b73d040580826121, /*  731 */
128'hb78d02400793943a12f6e76302000693, /*  732 */
128'ha8c948e502000313478145a147014681, /*  733 */
128'h954a9101020695130027e793a2110505, /*  734 */
128'h0200051392011602a865268500e50023, /*  735 */
128'h00094683c6e5460100e5736346119432, /*  736 */
128'h9f6300e90023471500e695630e500713, /*  737 */
128'h946347118bb10ff7f7930027979b0165, /*  738 */
128'h0037f713bded00c905a30086661300e7, /*  739 */
128'hf1279de3b7c501066613fed714e34685, /*  740 */
128'hf713f4e513e34711c51500b7c783709c, /*  741 */
128'h0004bc230004a623cb990207f7930047, /*  742 */
128'h4515f315bfd94511b72d4501e6070ae3, /*  743 */
128'hdbe58bc100b5c7836c8cfbe58b91b705, /*  744 */
128'h9a63b5a1c4c8ae4ff0ef0007c503609c, /*  745 */
128'h873245ad46a10ff7f7930027979b0565, /*  746 */
128'h7de3000747039722930117020017061b, /*  747 */
128'hf263fd370ae3f35709e3f3470be3f2e3, /*  748 */
128'h851700054c634185551b0187151b02b6, /*  749 */
128'h19e300080663000548030c2505130000, /*  750 */
128'hf3e30ff57513fbf7051bb5754519ef07, /*  751 */
128'h3701eca8efe30ff57513f9f7051beea8, /*  752 */
128'hec26f0227179bdc10ff777130017e793, /*  753 */
128'h0e500913451184aef406842ae44ee84a, /*  754 */
128'haecff0ef6008a0b1c90de199484c49bd, /*  755 */
128'h00b7c783c3210007c7036c1ce1292501, /*  756 */
128'h17e18bfd033780630327026303f7f793, /*  757 */
128'h64e2740270a2450100979a630017b793, /*  758 */
128'hbfdff0ef852245818082614569a26942, /*  759 */
128'h1101bfe54511b7cd00042a23d9452501, /*  760 */
128'h250187dff0ef842ae426ec06e8224581, /*  761 */
128'h2501a7eff0ef6008484c0e500493e50d, /*  762 */
128'h4585cb9900978d630007c7836c1ced09, /*  763 */
128'h00f513634791dd792501bb7ff0ef8522, /*  764 */
128'he82211018082610564a2644260e2451d, /*  765 */
128'he49d0005049bfa9ff0ef842aec06e426, /*  766 */
128'h6c08e0850005049ba34ff0ef6008484c, /*  767 */
128'h462d6c08700c838ff0ef458102000613, /*  768 */
128'h644260e200e782234705601c80eff0ef, /*  769 */
128'h4d1c08b7f06347858082610564a28526, /*  770 */
128'h842ae052e44eec26f406e84af0227179, /*  771 */
128'hf0ef852285ca59fd4a0506f5f063892e, /*  772 */
128'h64e2740270a24501e8910005049bed6f, /*  773 */
128'h8c6303448c63808261456a0269a26942, /*  774 */
128'hfd7125018abff0ef852285ca46010334, /*  775 */
128'he79300544783c81c278501378a63481c, /*  776 */
128'hfaf4e7e30004891b4c1c00f402a30017, /*  777 */
128'h713980824509bf4d4505bf5d4509bf65, /*  778 */
128'h832ff0eff42ee432e82efc061028ec2a, /*  779 */
128'h8733050ecb4787930000979704054263, /*  780 */
128'hc319676200070023c3196622631800a7, /*  781 */
128'h18634785cb114501e39897aa00070023, /*  782 */
128'h70e22501a02ff0ef0828080c460100f6, /*  783 */
128'hfca6e122e5067175bfe5452d80826121, /*  784 */
128'h302316050c63e42eecd6f0d2f4cef8ca, /*  785 */
128'h9ceff0ef1028002c8a7984aa89320005, /*  786 */
128'hb61ff0efe4be1028083c65a2e91d2501, /*  787 */
128'h799301c977934519e011e11964062501, /*  788 */
128'h102800f517634791c11510078e6301f9, /*  789 */
128'h794674e6640a60aac9052501e7dff0ef, /*  790 */
128'h451d00b44783808261496ae67a0679a6, /*  791 */
128'h00897913fff9452100497793f3fd8bc5, /*  792 */
128'h07937a220089e9936406a02108090a63, /*  793 */
128'h072300f40ca300f408a3021007130460, /*  794 */
128'h0ba300040b2300e40823000407a30004, /*  795 */
128'h0ea300040e23000405a300e40c230004, /*  796 */
128'h85a2000a450300040fa300040f230004, /*  797 */
128'h0a2300040da300040d234785f9bfe0ef, /*  798 */
128'h036300fa02230005091b00040aa30004, /*  799 */
128'h2501e1fff0ef030a2a83855285ca0209, /*  800 */
128'h80cff0ef0125262385d6397d7522fd21, /*  801 */
128'h79220209e993c3990089f793f1392501, /*  802 */
128'h85a3d09c01348523f4800309278385a2, /*  803 */
128'h01c40513c8c8f35fe0ef000945030004, /*  804 */
128'hae230004a623c88800695783daffe0ef, /*  805 */
128'h1de3bdf5450100f494230124b0230004, /*  806 */
128'hee0716e30107f713451100b44783ee05, /*  807 */
128'hec079ee3451d8b85fa0900e300297913, /*  808 */
128'he4d6e8d2eccef8a27119bdd14525bf51, /*  809 */
128'hf06af466f862fc5ee0daf0caf4a6fc86, /*  810 */
128'he0ef8ab6e4328a2e842a0006a023ec6e, /*  811 */
128'h662200b44783000998630005099be85f, /*  812 */
128'h790674a6854e744670e60007899bc39d, /*  813 */
128'h7d027ca27c427be26b066aa66a4669e6, /*  814 */
128'h16078c638b8500a44783808261096de2, /*  815 */
128'h00f67463893e40f907bb445c01042903, /*  816 */
128'h03040b131ff00c1320000b930006091b, /*  817 */
128'h120791631ff777934458fa090ae35cfd, /*  818 */
128'h01a7fd3337fd0025478300975d1b6008, /*  819 */
128'hec6347854848eb11020d19630ffd7d13, /*  820 */
128'hf0ef4c0cbfb5498900f405a3478900a7, /*  821 */
128'h00f405a3478501951763b7e52501bc6f, /*  822 */
128'hf0efe43e853e4c0c601ccc08b7954985, /*  823 */
128'h8dc200a6083b000d061bd5792501b86f, /*  824 */
128'h873b0099549b0027c683072c7a6367a2, /*  825 */
128'h86a60017c50341a684bb00e6f46300c4, /*  826 */
128'h00a44783f9452501176050ef85d28642, /*  827 */
128'h0097fc6341b507bb4c48c3850407f793, /*  828 */
128'h955285da20000613910115020097951b, /*  829 */
128'h9a3e9381020497930094949bc3ffe0ef, /*  830 */
128'h9fa5000aa783c45c9fa54099093b445c, /*  831 */
128'h00a44703050601634c50bf3900faa023, /*  832 */
128'he44285da46850017c503c30d04077713, /*  833 */
128'hf793682200a44783f131250113c050ef, /*  834 */
128'h0017c50386424685601c00f40523fbf7, /*  835 */
128'h444c01b42e23f10d25010e8050ef85da, /*  836 */
128'h0127746340bb873b1ff5f5930009049b, /*  837 */
128'he0ef855295a28626030585930007049b, /*  838 */
128'heccef0caf8a27119b585499dbf9dbb1f, /*  839 */
128'hf466f862fc5ee0daf4a6fc86e4d6e8d2, /*  840 */
128'h8ab689328a2e842a0006a023ec6ef06a, /*  841 */
128'h00b44783000997630005099bca3fe0ef, /*  842 */
128'h790674a6854e744670e60007899bc39d, /*  843 */
128'h7d027ca27c427be26b066aa66a4669e6, /*  844 */
128'h1a0782638b8900a44783808261096de2, /*  845 */
128'h0c1320000b9304f76e630127873b445c, /*  846 */
128'h77930409046344585cfd03040b131ff0, /*  847 */
128'h0025478300975d1b6008140794631ff7, /*  848 */
128'hef01040d1a630ffd7d1301a7fd3337fd, /*  849 */
128'h05a3478902e798634705cb914581485c, /*  850 */
128'h0005079bd6aff0ef4c0cb749498900f4, /*  851 */
128'he79300a4478312f76b634818445cf3fd, /*  852 */
128'h05a3478501979763b78500f405230207, /*  853 */
128'h4783c85ce311cc1c4858bf89498500f4, /*  854 */
128'hc50346854c50601cc38d0407f79300a4, /*  855 */
128'h00a44783f96925017d9040ef85da0017, /*  856 */
128'he43e853e4c0c601c00f40523fbf7f793, /*  857 */
128'h00a8063b000d081bd1592501964ff0ef, /*  858 */
128'h0099549b0027c683072c7a6367a28db2, /*  859 */
128'h0017c50341a684bb00e6f4630104873b, /*  860 */
128'h87bb4c4cf1492501789040ef85d286a6, /*  861 */
128'h0613918115820097959b0297f26341b5, /*  862 */
128'hf79300a44783a29fe0ef855a95d22000, /*  863 */
128'h9381020497930094949b00f40523fbf7, /*  864 */
128'h000aa783c45c9fa54099093b445c9a3e, /*  865 */
128'h481400c70e634c58bdc900faa0239fa5, /*  866 */
128'h40ef85da46850017c50300d77a634458, /*  867 */
128'h0009049b444801b42e23fd0125016ed0, /*  868 */
128'h0007049b0127746340ab873b1ff57513, /*  869 */
128'h47839b5fe0ef952285d2862603050513, /*  870 */
128'hb5f1c81cbf4100f405230407e79300a4, /*  871 */
128'hab7fe0ef842ae406e0221141bd15499d, /*  872 */
128'hf793cf610207f71300a44783e16d2501, /*  873 */
128'h05930017c50346854c50601cc3950407, /*  874 */
128'hf79300a44783ed4d25016ab040ef0304, /*  875 */
128'h2501b5ffe0ef6008500c00f40523fbf7, /*  876 */
128'h00e785a30207671300b7c703741ce155, /*  877 */
128'h8e230086d69b0106d69b0107169b4818, /*  878 */
128'h8f230187571b0107569b00d78ea300e7, /*  879 */
128'h00078ba300078b23485800e78fa300d7, /*  880 */
128'h00e78a230107571b0107169b00e78d23, /*  881 */
128'h00e78aa30087571b0107571b0107171b, /*  882 */
128'h0086d69b00e78c23021007130106d69b, /*  883 */
128'h0007892300e78ca300d78da304600713, /*  884 */
128'h0523fdf7f793600800a44783000789a3, /*  885 */
128'he06f014160a2640200f50223478500f4, /*  886 */
128'he022114180820141640260a24505ea3f, /*  887 */
128'he0ef8522e9012501f01ff0ef842ae406, /*  888 */
128'h0141640260a200043023e11925019b5f, /*  889 */
128'h4a63945fe0efec060028e42a11018082, /*  890 */
128'h610560e245015ca78b23000087970005, /*  891 */
128'h1028002c4601e42a7159bfe5452d8082, /*  892 */
128'hec190005041bb25fe0efeca6f486f0a2, /*  893 */
128'h0005041bcb4ff0efe4be1028083c65a2, /*  894 */
128'h70a68522cbd8575277a2e9916586e41d, /*  895 */
128'hcb998bc100b5c7838082616564e67406, /*  896 */
128'h4791b7c5c8c8965fe0ef0004c50374a2, /*  897 */
128'he506e42afca67175bfd94415fcf41ee3, /*  898 */
128'h002c460184ae00050023f4cef8cae122, /*  899 */
128'h77e2ecbe081ce5212501ab9fe0ef1828, /*  900 */
128'h040991634996c2be4bdc02f009138426, /*  901 */
128'h071b5227470300008717e50567a24501, /*  902 */
128'h156300e780a303a0071300e780230307, /*  903 */
128'h00078023078d00e7812302f007130e94, /*  904 */
128'h45858082614979a6794674e6640a60aa, /*  905 */
128'hf0ef18284581fd4d2501f75fe0ef1828, /*  906 */
128'he0ef0007c50365c677e2f55d2501e6cf, /*  907 */
128'hf9512501f4ffe0ef18284581c2aa8bdf, /*  908 */
128'h65c677e2e1052501e46ff0ef18284581, /*  909 */
128'h458101350e632501897fe0ef0007c503, /*  910 */
128'h12e367a24711dd612501a86ff0ef1828, /*  911 */
128'h4781f48fe0ef1828100cb7614509f6e5, /*  912 */
128'he705fc97470397361094930102079713, /*  913 */
128'h662236fd86a285be04e460630037871b, /*  914 */
128'h0023fff7c793e989963a930102069713, /*  915 */
128'h059bfff5871bb7e12785bf199c3d0126, /*  916 */
128'h0023fc974703972a1088930117020007, /*  917 */
128'h0204169367220789bdf54545b7e900e6, /*  918 */
128'hfee78fa3240507850007470397369281, /*  919 */
128'hfc06f04af426f8227139b721fe9465e3, /*  920 */
128'h091bfa8fe0ef84ae842ae456e852ec4e, /*  921 */
128'h0007891bcf8900b44783000917630005, /*  922 */
128'h6aa26a4269e2790274a2854a744270e2, /*  923 */
128'h8b8900a4478300977763481880826121, /*  924 */
128'h4818445ce4bd00042623445884bae391, /*  925 */
128'h05230207e79300a44783c81cfcf778e3, /*  926 */
128'h4c50d3e51ff7f793445c4481bf7d00f4, /*  927 */
128'h0407f7930304099300a44783fc960ee3, /*  928 */
128'h341040ef0017c50385ce4685601cc385, /*  929 */
128'h00f40523fbf7f79300a44783ed512501, /*  930 */
128'h2ef040ef85ce0017c50386264685601c, /*  931 */
128'h999b002547836008bf59cc44ed352501, /*  932 */
128'h563b0336d6bbfff4869b377dc7290097, /*  933 */
128'h27814c0c8ff9413007bb02c6ed630337, /*  934 */
128'h445c0499ea634a855a7dd1c19c9dc45c, /*  935 */
128'hc79fe0ef6008d7b51ff4f793c45c9fa5, /*  936 */
128'he595484cbfb19ca90094d49bcd112501, /*  937 */
128'h478900f5976347850005059b802ff0ef, /*  938 */
128'h478500f5976357fdbded490900f405a3, /*  939 */
128'h4783b765cc0cc84cb5ed490500f405a3, /*  940 */
128'h0005059bfcbfe0efcb818b89600800a4, /*  941 */
128'h88e30005059bc3ffe0efbf6984cee599, /*  942 */
128'h445cfaf5fae34f9c601cfabafee3fd45, /*  943 */
128'h7139b7bdc45c013787bb413484bbcc0c, /*  944 */
128'h0828002c4601842ac52de42ef822fc06, /*  945 */
128'he01c852265a267e2e1152501fdafe0ef, /*  946 */
128'hcd996c0ce5292501968ff0eff01c101c, /*  947 */
128'ha02d000430234515e7898bc100b5c783, /*  948 */
128'h458167e2c448e24fe0ef0007c50367e2, /*  949 */
128'h2501cadfe0ef00f414230067d7838522, /*  950 */
128'h80826121744270e2f971fcf50be34791, /*  951 */
128'he0221141b7c1fcf501e34791bfdd4525, /*  952 */
128'h00043023e1192501daefe0ef842ae406, /*  953 */
128'he84aec26f022717980820141640260a2, /*  954 */
128'he8890005049bd8cfe0ef892e842af406, /*  955 */
128'h0005049bc4ffe0ef8522458100091f63, /*  956 */
128'h30238082614564e269428526740270a2, /*  957 */
128'h136347912501b34ff0ef852245810224, /*  958 */
128'h4581c58fe0ef852285ca00042a2302f5, /*  959 */
128'h2a2300f5166347912501f77fe0ef8522, /*  960 */
128'he42aeca67159bf6584aad16dbf7d0004, /*  961 */
128'hecefe0eff486f0a21028002c460184ae, /*  962 */
128'hf0efe4be1028083c65a2e00d0005041b, /*  963 */
128'h85a6c489cf816786e8010005041b85ef, /*  964 */
128'h616564e6740670a68522c00fe0ef1028, /*  965 */
128'he42af85a8432f0a27159bfcd44198082, /*  966 */
128'he8caeca6f486e0d28522002c46018b2e, /*  967 */
128'h0a1be70fe0efec66f062f45efc56e4ce, /*  968 */
128'h871b481c01842c836000000a1c630005, /*  969 */
128'h8552740670a600fb202302f76263ffec, /*  970 */
128'h7c027ba27b427ae26a0669a6694664e6, /*  971 */
128'h02fb9f63478500044b83808261656ce2, /*  972 */
128'ha49fe0ef852285ca4a8559fd44814909, /*  973 */
128'h4c1c2485e11109550863093508632501, /*  974 */
128'h0017e793c80400544783fef963e32905, /*  975 */
128'h10000ab7504cb74d009b202300f402a3, /*  976 */
128'h852200099e631afd4c09448149814901, /*  977 */
128'h091385cee9212501d04fe0ef0015899b, /*  978 */
128'h470300194783038b9163200009930344, /*  979 */
128'h39f909092485e3918fd90087979b0009, /*  980 */
128'haa2fe0efe02e854ab745fc0c94e33cfd, /*  981 */
128'h39f109112485e1116582015575332501, /*  982 */
128'h1101bfad8a2abfbd4a09b7494a05b7c5, /*  983 */
128'h049bbb8fe0ef842ae04aec06e426e822, /*  984 */
128'h60e20007849bcb9100b44783e4910005, /*  985 */
128'h00a447838082610564a2690285266442, /*  986 */
128'he793fed772e348144458cf390027f713, /*  987 */
128'hf0ef484cef01600800f40523c8180207, /*  988 */
128'h84aa00a405a3c53900042a232501a5af, /*  989 */
128'h146357fd0005091b941fe0ef4c0cbf7d, /*  990 */
128'he0ef167d100006374c0cb7dd450502f9, /*  991 */
128'h2501a1eff0ef85ca6008f9792501b25f, /*  992 */
128'h6008fcf900e345094785b769449db7e1, /*  993 */
128'hdba50407f79300a44783fcf96ae34d1c, /*  994 */
128'h40ef030405930017c50346854c50601c, /*  995 */
128'h0523fbf7f79300a44783f55d250171e0, /*  996 */
128'he5061008002c4605e42a7175b7b100f4, /*  997 */
128'h65a2e9052501c94fe0eff8cafca6e122, /*  998 */
128'h6786e1052501e27fe0efe0be1008081c, /*  999 */
128'hc59975e2eb890207f79300b7c7834519, /* 1000 */
128'h640a60aa451dcb810014f79300b5c483, /* 1001 */
128'he0ef00094503790280826149794674e6, /* 1002 */
128'h01492783c89d88c1cc0d0005041baccf, /* 1003 */
128'h952fe0ef00a8100c02800613fc878de3, /* 1004 */
128'h4581f1612501941fe0efcaa200a84589, /* 1005 */
128'hfaf518e34791d94d2501838ff0ef00a8, /* 1006 */
128'he0ef7502e411f15525019e3fe0ef1008, /* 1007 */
128'h250191eff0ef85a27502bf612501f12f, /* 1008 */
128'hf1221028002c4605e42a7171b7edf551, /* 1009 */
128'hf4def8dafcd6e152e54ee94aed26f506, /* 1010 */
128'h12630005041bbc4fe0efe8eaece6f0e2, /* 1011 */
128'h041bd53fe0efe4be1028083c65a21c04, /* 1012 */
128'h441967a61af4156347911c0407630005, /* 1013 */
128'h4581752218079d630207f79300b7c783, /* 1014 */
128'h75224785180480630005049bb33fe0ef, /* 1015 */
128'he0ef16f48863440557fd16f48c634409, /* 1016 */
128'hd91b85a67422160412630005041ba8cf, /* 1017 */
128'h2000061303440b13f60fe0ef85220104, /* 1018 */
128'h0593462d886fe0ef855a00050c1b4581, /* 1019 */
128'h999b0ff97a9347c187afe0ef855a0200, /* 1020 */
128'h07930109d99b02f40fa30109191b0104, /* 1021 */
128'hfa1304f4062302e00b930109591b0210, /* 1022 */
128'h06a30089591b0089d99b046007930ff4, /* 1023 */
128'h05a30404052303740a230200061304f4, /* 1024 */
128'h04a305540423053407a3054407230404, /* 1025 */
128'h0aa37722ff7fd0ef0544051385da0524, /* 1026 */
128'h571400d6166357d200074603468d0574, /* 1027 */
128'hd79b0107969b06f40723478100f69363, /* 1028 */
128'hd79b0106d69b0107979b06f404230107, /* 1029 */
128'h04a306d407a30087d79b0086d69b0107, /* 1030 */
128'he0ef1028040b99634c8500274b8306f4, /* 1031 */
128'h85a3752247416786e8350005041bf5ff, /* 1032 */
128'h8b230460071300e78c230210071300e7, /* 1033 */
128'h8da301478d2300e78ca300078ba30007, /* 1034 */
128'h00f50223478501278aa301578a230137, /* 1035 */
128'h001c0d1b7522a82d0005041bd50fe0ef, /* 1036 */
128'h0005041b8d4fe0ef0195022303852823, /* 1037 */
128'hf53fd0ef3bfd855a458120000613ec09, /* 1038 */
128'he0ef85a67522441db7498c6a0ffbfb93, /* 1039 */
128'h6a0a69aa694a64ea740a70aa8522f2bf, /* 1040 */
128'h8082614d6d466ce67c067ba67b467ae6, /* 1041 */
128'h843284aee42aeca6f0a27159b7c54421, /* 1042 */
128'he13125019c2fe0eff48610284605002c, /* 1043 */
128'he9152501b55fe0efe4be1028083c65a2, /* 1044 */
128'h6706e39d0207f79300b7c783451967a6, /* 1045 */
128'h027474138c658cbd752200b74783c30d, /* 1046 */
128'hc94fe0ef00f502234785008705a38c3d, /* 1047 */
128'he42a71718082616564e6740670a62501, /* 1048 */
128'he0efed26f122f5060088002c4605e02e, /* 1049 */
128'h008865a26786120795630005079b95cf, /* 1050 */
128'h99630005079bae7fe0eff0be083cf4be, /* 1051 */
128'h116302077713479900b7c70377861007, /* 1052 */
128'h102805ad46550e058d63479165e61007, /* 1053 */
128'he33fd0ef10a8008c02800613e3ffd0ef, /* 1054 */
128'h10a865820c054c6347adefdfd0ef850a, /* 1055 */
128'h0ce792634711cbf10005079ba9dfe0ef, /* 1056 */
128'h464d648aebdd0005079bdcbfe0ef10a8, /* 1057 */
128'h02814783df7fd0ef00d4851302a10593, /* 1058 */
128'h00f40223478500f485a30207e7936406, /* 1059 */
128'h06f7076357d64736cbb58bc100b4c783, /* 1060 */
128'h85220005059bf25fd0ef85a600044503, /* 1061 */
128'hd0ef8522c1bd47890005059bca4fe0ef, /* 1062 */
128'h468302e007936706efa90005079bfbbf, /* 1063 */
128'h06f707230107969b57d602f69c630557, /* 1064 */
128'h0107d79b0107979b06f704230107d79b, /* 1065 */
128'h06f704a30086d69b0106d69b0087d79b, /* 1066 */
128'he18fe0ef008800f7022306d707a34785, /* 1067 */
128'h0005079bb48fe0ef6506e7910005079b, /* 1068 */
128'hbfcd47a18082614d853e64ea740a70aa, /* 1069 */
128'hec861028002c4605842ee42ae8a2711d, /* 1070 */
128'he4be1028083c65a2e929250180afe0ef, /* 1071 */
128'h00b7c783451967a6e129250199dfe0ef, /* 1072 */
128'h752200645703cb856786eb950207f793, /* 1073 */
128'h0044570300e78ba30087571b00e78b23, /* 1074 */
128'h0223478500e78ca30087571b00e78c23, /* 1075 */
128'h80826125644660e62501acefe0ef00f5, /* 1076 */
128'h4601002c893284aee42ae0cae4a6711d, /* 1077 */
128'he0510005041bf95fd0efec86e8a20828, /* 1078 */
128'he5592501c9efe0efd20208284581c4b9, /* 1079 */
128'h462d75c2e93d2501b97fe0ef08284585, /* 1080 */
128'h0200061346ad00b48713c8dfd0ef8526, /* 1081 */
128'h17820007869bfff6879bce8900070023, /* 1082 */
128'h0a63fec783e3177d0007c78397a69381, /* 1083 */
128'he0150005041be63fd0ef510c65620209, /* 1084 */
128'h00e684630005468304300793470d6562, /* 1085 */
128'h2023c15fd0ef953e0347879302700793, /* 1086 */
128'h80826125690664a6644660e6852200a9, /* 1087 */
128'hb7d5842abf550004802300f515634791, /* 1088 */
128'hd0efec86e8a21028002c4605e42a711d, /* 1089 */
128'h478100010c236522e4710005041beddf, /* 1090 */
128'h0613eb2900074703972a930102079713, /* 1091 */
128'h041bbccfe0efda0210284581ebb10200, /* 1092 */
128'h15632501ac3fe0ef10284585e0450005, /* 1093 */
128'hd0ef082c462dc7e56506018147831005, /* 1094 */
128'h0460071300e78c23021007136786bb1f, /* 1095 */
128'h2785a0e900e78ca300078ba300078b23, /* 1096 */
128'h928102071693fff7871bb77d87bab745, /* 1097 */
128'h432d48e54701fec686e30006c68396aa, /* 1098 */
128'h030596930017061b0006c58300e506b3, /* 1099 */
128'h0108ec63030858131842f9f6881b92c1, /* 1100 */
128'h8e1bada585930000759792c116c23681, /* 1101 */
128'hfeb045e34185d59b0185959ba8310006, /* 1102 */
128'hc803058580826125644660e685224419, /* 1103 */
128'hfe6702e3b7ddffc81be3000805630005, /* 1104 */
128'he9e30007069b00d58023070595ba082c, /* 1105 */
128'h869b020006134729938102061793f8f6, /* 1106 */
128'h13e30e5007930181470300d779630007, /* 1107 */
128'hb7c5078500c6802396be0834b77df0f7, /* 1108 */
128'he0ef00f502234785752200f500235795, /* 1109 */
128'h478302f51b634791b7710005041b8b2f, /* 1110 */
128'hf8350005041ba19fe0ef1028d3c10181, /* 1111 */
128'h462d6506ab7fd0ef4581020006136506, /* 1112 */
128'hbdd100e785a347216786a8dfd0ef082c, /* 1113 */
128'h0585230305452e0305052e83bf81842a, /* 1114 */
128'h02938f2ae44ae826ec22110105c52883, /* 1115 */
128'h8f9300005f97887687f2869a86460405, /* 1116 */
128'h000fa38300b647338dfd00c6c5b3636f, /* 1117 */
128'h9db9007585bb0fc1008fa403000f2583, /* 1118 */
128'h0078159b0105883b004f2703ff4fa383, /* 1119 */
128'h00f805bb0077073b0105e8330198581b, /* 1120 */
128'h9e39008f23838e358e6d00f6c6339f31, /* 1121 */
128'h873b008383bb8e590146561b00c6171b, /* 1122 */
128'h00cf24038ef900b7c6b300d383bb00c5, /* 1123 */
128'he6b30116969b00f6d39b007686bb8ebd, /* 1124 */
128'h0007061b00d703bbffcfa4039fa100d3, /* 1125 */
128'h00a7579b9f3d8f2d9fa1007777338f2d, /* 1126 */
128'h0003869b0005881b0f418f5d0167171b, /* 1127 */
128'h678f0f1300005f17f45f17e300e387bb, /* 1128 */
128'h67828293000052975b0f8f9300005f97, /* 1129 */
128'h4383000fa58300b6c7338df100d7c5b3, /* 1130 */
128'h93aa038a000f47039db9002f4403001f, /* 1131 */
128'h004fa7039db9942a040a4318972a070a, /* 1132 */
128'ha70301b8581b9e390058159b0105883b, /* 1133 */
128'h00b7c6339f3100f805bb0105e8330003, /* 1134 */
128'h561b0096139b008fa7039e398e3d8e75, /* 1135 */
128'h9f3500c583bb00c3e63340189eb90176, /* 1136 */
128'h0fc18eadffff44838efd0075c6b30f11, /* 1137 */
128'h9fb900e6941b94aa048affcfa7039eb9, /* 1138 */
128'hc7339fb900d3843b8ec140980126d69b, /* 1139 */
128'h171b00c7579b9f3d007747338f6d0083, /* 1140 */
128'h0004069b0003861b0005881b8f5d0147, /* 1141 */
128'h598f8f9300005f97f25f1ee300e407bb, /* 1142 */
128'ha7030102c40350e383930000539782fe, /* 1143 */
128'h400000c5c4b3942a040a00d7c5b30003, /* 1144 */
128'h94aa048a0043a4039f210112c4839f25, /* 1145 */
128'h0048171b0122c4830107083b40809e21, /* 1146 */
128'h073b0083a4039e210107683301c8581b, /* 1147 */
128'h159b40809e2d9ea194aa8db9048a00f8, /* 1148 */
128'h05bb03c18e4d0156561b0132c90300b6, /* 1149 */
128'h090a8ead00e7c6b3ffc3a4839c3500c7, /* 1150 */
128'h24830106d69b9fa50106941b992a9ea1, /* 1151 */
128'h9fa58f2d0007081b00d5843b8ec10009, /* 1152 */
128'h02918f5d0177171b0097579b9f3d8f21, /* 1153 */
128'hf45f17e300e407bb0004069b0005861b, /* 1154 */
128'h45b38f5dfff647134902829300005297, /* 1155 */
128'h9f2d022fc403021fc3830002a70300d7, /* 1156 */
128'h040a418c95aa058a93aa038a020fc583, /* 1157 */
128'h0068171b0107083b0042a5839f2d942a, /* 1158 */
128'h073b0107683301a8581b0003a5839e2d, /* 1159 */
128'ha5839e2d8e3d8e59fff6c6139db100f8, /* 1160 */
128'he633400c9ead0166561b00a6139b0082, /* 1161 */
128'hfff7c593023fc4839ead00c703bb00c3, /* 1162 */
128'h048a9db5ffc2a4038db902c10075e5b3, /* 1163 */
128'h40809fa18dd50115d59b94aa00f5969b, /* 1164 */
128'h9fa18f4dfff747130007081b00b385bb, /* 1165 */
128'h8f5d0157171b00b7579b9f3d00774733, /* 1166 */
128'h1de300e587bb0005869b0003861b0f91, /* 1167 */
128'h00d306bb00fe07bb010e883b6462f3ff, /* 1168 */
128'h64c2cd70cd34c97c0505282300c8863b, /* 1169 */
128'hf84afc26e0a2715d653c808261056922, /* 1170 */
128'h03f7f413ec56f052e486e45ee85af44e, /* 1171 */
128'h0b9304000b13e53c893289ae84aa97b2, /* 1172 */
128'h74639381178200078a1b408b07bb0400, /* 1173 */
128'h85ce020ada93020a1a9300090a1b00f9, /* 1174 */
128'h09334a7020ef0144043b865600848533, /* 1175 */
128'h97824401852660bc0174176399d64159, /* 1176 */
128'h6ae27a0279a2794274e2640660a6b7c9, /* 1177 */
128'hf793f0227179653c808261616ba26b42, /* 1178 */
128'h00178513e84af406e44eec26842a03f7, /* 1179 */
128'h449d0400099300e7802397a2f8000713, /* 1180 */
128'h95224581920116020006091b40a9863b, /* 1181 */
128'h603cfc1c078e643c0124f5633f3020ef, /* 1182 */
128'h64e2740270a2fd24fde3450197828522, /* 1183 */
128'h14878793000077978082614569a26942, /* 1184 */
128'h1407879300007797e93c04053423639c, /* 1185 */
128'h8082e13cb807879300000797ed3c639c, /* 1186 */
128'h3e5020efec06850a4641050505931101, /* 1187 */
128'h85930000659734e68693000076974701, /* 1188 */
128'h070506890007c78300e107b345415765, /* 1189 */
128'hc78397ae000646038bbd962e0047d613, /* 1190 */
128'h60e2fca71de3fef68fa3fec68f230007, /* 1191 */
128'he1227175808261053105051300007517, /* 1192 */
128'h85a26622f71ff0efe42ee5060808842a, /* 1193 */
128'hf0ef0808f01ff0ef0808e85ff0ef0808, /* 1194 */
128'h711c46a1595880826149640a60aaf83f, /* 1195 */
128'hcf980200071300d71763469100d70d63, /* 1196 */
128'h11018082556dbfe50007ac2380824501, /* 1197 */
128'h026384ae842a420007b7ec06e426e822, /* 1198 */
128'h65970880061323e686930000569702f5, /* 1199 */
128'h30ef4ea50513000065174da585930000, /* 1200 */
128'h11018082610564a2644260e2fc241d30, /* 1201 */
128'h026384ae420007b7ec06e4266100e822, /* 1202 */
128'h659702f00613216686930000569702f4, /* 1203 */
128'h30ef4aa505130000651749a585930000, /* 1204 */
128'h11018082610564a2644260e2e0041930, /* 1205 */
128'h026384ae420007b7ec06e4266100e822, /* 1206 */
128'h6597036006131e6686930000569702f4, /* 1207 */
128'h30ef46a505130000651745a585930000, /* 1208 */
128'h11018082610564a2644260e2e4041530, /* 1209 */
128'h8263842e420007b7ec06e8226104e426, /* 1210 */
128'h659703e0061300e686930000769702f4, /* 1211 */
128'h30ef42a505130000651741a585930000, /* 1212 */
128'h610564a2644260e2e880900114021130, /* 1213 */
128'h420007b7ec06e8226104e42611018082, /* 1214 */
128'h0613fc2686930000769702f48263842e, /* 1215 */
128'h0513000065173d658593000065970450, /* 1216 */
128'h644260e2ec80900114020cf030ef3e65, /* 1217 */
128'hec06e4266100e82211018082610564a2, /* 1218 */
128'h86930000569702f4026384ae420007b7, /* 1219 */
128'h6517392585930000659704c0061312e6, /* 1220 */
128'h644260e2f00408b030ef3a2505130000, /* 1221 */
128'hec06e4266100e82211018082610564a2, /* 1222 */
128'h86930000569702f4026384ae420007b7, /* 1223 */
128'h65173525859300006597053006130fe6, /* 1224 */
128'h644260e2f40404b030ef362505130000, /* 1225 */
128'hf82200053983ec4e71398082610564a2, /* 1226 */
128'h8436893284ae420007b7fc06f04af426, /* 1227 */
128'h05a006130c4686930000569702f98463, /* 1228 */
128'h31850513000065173085859300006597, /* 1229 */
128'h8b0588090014141b67227fe030efe43a, /* 1230 */
128'h64330034949b8c59004979130029191b, /* 1231 */
128'h74a2744270e20289b8238c4588a10124, /* 1232 */
128'h47057100e02211418082612169e27902, /* 1233 */
128'h8522f7dff0efe4064581852246054681, /* 1234 */
128'h45814605468547058522f35ff0ef4581, /* 1235 */
128'h640260a2d97ff0ef45816008f67ff0ef, /* 1236 */
128'h46814705e022e4061141808201414501, /* 1237 */
128'hf0ef842a45810405302302053c234605, /* 1238 */
128'h470545818522ef1ff0ef45818522f39f, /* 1239 */
128'h458160a264026008f23ff0ef46054685, /* 1240 */
128'hec06e8226104e4261101d4dff06f0141, /* 1241 */
128'h86930000569702f48263842e420007b7, /* 1242 */
128'h6517222585930000659706100613fee6, /* 1243 */
128'hfc809041144271a030ef232505130000, /* 1244 */
128'h6104e42611018082610564a2644260e2, /* 1245 */
128'h569702f48263842e420007b7ec06e822, /* 1246 */
128'h85930000659706800613fba686930000, /* 1247 */
128'h14526d6030ef1ee50513000065171de5, /* 1248 */
128'h11018082610564a2644260e2e0a09051, /* 1249 */
128'h026384ae420007b7ec06e4266100e822, /* 1250 */
128'h659706f00613f86686930000569702f4, /* 1251 */
128'h30ef1aa505130000651719a585930000, /* 1252 */
128'h11018082610564a2644260e2e4246920, /* 1253 */
128'h420007b7ec06e426e82200053903e04a, /* 1254 */
128'hf50686930000569702f9026384ae842a, /* 1255 */
128'h00006517154585930000659707600613, /* 1256 */
128'h60e2c84404993c2364c030ef16450513, /* 1257 */
128'h7100f0a2715980826105690264a26442, /* 1258 */
128'hf45ef85afc56e0d2e4cef486e8caeca6, /* 1259 */
128'h84b2892e0005d783020408a3ec66f062, /* 1260 */
128'h6f6020ef00c9051345814611d01ce030, /* 1261 */
128'h00043983bf7ff0ef458560080e049c63, /* 1262 */
128'h0049278316f99a6304043a03420007b7, /* 1263 */
128'h4485e391448d8b89c7090017f7134481, /* 1264 */
128'h008a2783000a09638cdd03243c234c1c, /* 1265 */
128'h4605468147050144e493160786638b85, /* 1266 */
128'hbe3ff0ef85224581d73ff0ef85224581, /* 1267 */
128'h5583c55ff0ef00989a37852200892583, /* 1268 */
128'h852285a6c8bff0ef681a0a1385220009, /* 1269 */
128'h46854705cffff0ef85224581cc7ff0ef, /* 1270 */
128'h8593000f45b7d31ff0ef852245814605, /* 1271 */
128'hcdbff0ef85224585e9bff0ef85222405, /* 1272 */
128'he593e7ac8c9300005c9785220d89b583, /* 1273 */
128'h030a8a9300006a97ebbff0ef25810015, /* 1274 */
128'h740670a6efe9485c040b0b1300006b17, /* 1275 */
128'h7c027ba27b427ae26a0669a6694664e6, /* 1276 */
128'hf0efe024852244cc8082616545016ce2, /* 1277 */
128'h9be38b85449cdf5ff0ef8522488cdb9f, /* 1278 */
128'h63900107e683654100043883603cee07, /* 1279 */
128'hf005051300ff0e374311470147814581, /* 1280 */
128'h070500371f1b00064803ec0689e36e89, /* 1281 */
128'h036316fd060527810107e7b301e8183b, /* 1282 */
128'h010767330187971b0187d81bf2e50067, /* 1283 */
128'h010767330087d79b01c878330087981b, /* 1284 */
128'h938183751782170200be873b8fd98fe9, /* 1285 */
128'h00005697b765470147812585e31c9746, /* 1286 */
128'hf60585930000659714900613d6c68693, /* 1287 */
128'he493bd85458030eff705051300006517, /* 1288 */
128'h000b9d633bfd42000c378bd2bd6100c4, /* 1289 */
128'hf605051300006517d505859300005597, /* 1290 */
128'h86e60189096300043903b711702000ef, /* 1291 */
128'h07093483418030ef855a85d60f200613, /* 1292 */
128'h020937031404806324818cfd4981485c, /* 1293 */
128'hf9200793c7817c1c00f76f630c893783, /* 1294 */
128'hf0ef85224581b71ff0ef85224581cc5c, /* 1295 */
128'h7913852201442903c39d0044f793b29f, /* 1296 */
128'h85cad45ff0ef85ca290100896913ff39, /* 1297 */
128'h0084f79368a000eff005051300006517, /* 1298 */
128'h00496913ff397913852201442903c39d, /* 1299 */
128'h05130000651785cad1bff0ef85ca2901, /* 1300 */
128'h00043983cfb50014f793660000efefe5, /* 1301 */
128'hcb8686930000569701898c6303843903, /* 1302 */
128'hcba97c1c368030ef855a85d609c00613, /* 1303 */
128'h9f630037f693470d02043c2300492783, /* 1304 */
128'h4591480d468100c907930189871308e6, /* 1305 */
128'h01068763c3900086161bff8705136310, /* 1306 */
128'h0791872a2685c3988f518361ff873703, /* 1307 */
128'hc85c0027e793485ccbb5603cfeb690e3, /* 1308 */
128'h39036004cc9d49858889c85c9bf9485c, /* 1309 */
128'h0613c52686930000569701848c630404, /* 1310 */
128'h0963040430232ea030ef855a85d60ca0, /* 1311 */
128'hb4bff0ef8522ef8d8b85008927830009, /* 1312 */
128'hc43ff0ef8522484cc85c9bf54985485c, /* 1313 */
128'hdbd98b85bd85677020ef4505d8098ce3, /* 1314 */
128'hb1bff0ef8522b77100f926230009b783, /* 1315 */
128'hdcd5010964830009398397a667a1bf41, /* 1316 */
128'h20efe43e002c4621854e639c00878913, /* 1317 */
128'h08b041635535b7dd87ca14e109a13c20, /* 1318 */
128'he44ef406e84aec26f022048005137179, /* 1319 */
128'h85a2c41d5551842a1dc030ef892e84b2, /* 1320 */
128'h85aa89aa7b3010efbc05051300005517, /* 1321 */
128'h9d63508000efdce50513000065178622, /* 1322 */
128'h64e2740270a2557d1f6030ef85220009, /* 1323 */
128'h2423e01c420007b78082614569a26942, /* 1324 */
128'h4501c45c4789c7890024f793f4040124, /* 1325 */
128'h8082b7f9c45c4785d8f145018885bfe9, /* 1326 */
128'h07b7050ef73ff06f4200053745814609, /* 1327 */
128'he0221141711c80822501638897aa4200, /* 1328 */
128'h0000569702f40263420007b7e4066380, /* 1329 */
128'hcb0585930000659734c00613b5c68693, /* 1330 */
128'h4505703c1a8030efcc05051300006517, /* 1331 */
128'he822110180820141640260a2557de391, /* 1332 */
128'h644285a2501010efe42eec064501842a, /* 1333 */
128'h051371797a00006f6105468560e26622, /* 1334 */
128'h30efe052e44ee84aec26f022f4062000, /* 1335 */
128'h1ea030efd24505130000651784aa0e20, /* 1336 */
128'h842a4bf010ef4501479010ef0001b503, /* 1337 */
128'h638cd0a5051300006517681c224010ef, /* 1338 */
128'hd08505130000651706f44583402000ef, /* 1339 */
128'hd59bd125051300006517546c3f2000ef, /* 1340 */
128'h06c4458358303dc000ef91c115c20085, /* 1341 */
128'h0106569b0086571bd085051300006517, /* 1342 */
128'h0186561b0ff6f6930ff777130ff67793, /* 1343 */
128'h00efcfa50513000065175c0c3b2000ef, /* 1344 */
128'h6597c789c845859300006597545c3a40, /* 1345 */
128'h00efcea5051300006517c72585930000, /* 1346 */
128'h744813c030efcf650513000065173840, /* 1347 */
128'h19c42783daffb0ef2f85859300006597, /* 1348 */
128'h00006617e789c4e6061300006617584c, /* 1349 */
128'h346000efcd45051300006517fac60613, /* 1350 */
128'h0a1300006a174401ed9ff0ef85264581, /* 1351 */
128'h779320000913cd69899300006997cd6a, /* 1352 */
128'h87b3318000ef8552e7810004059b01f4, /* 1353 */
128'h819100f5f6130405854e0007c5830084, /* 1354 */
128'h2805051300006517fd241de3302000ef, /* 1355 */
128'h6a0269a2694264e2740270a22f2000ef, /* 1356 */
128'hb6830083b7830103b703808261454501, /* 1357 */
128'h00d7fe6393811782278540f707b30003, /* 1358 */
128'h0103b78300a7002300f3b82300170793, /* 1359 */
128'h0083b703808245018082000780234505, /* 1360 */
128'h0003b7038f999201020596130103b783, /* 1361 */
128'h9d9dfff7059b00c6f5638e9dfff70693, /* 1362 */
128'h002300b6e6630103b7030007869b4781, /* 1363 */
128'h06b300d3b823001706938082852e0007, /* 1364 */
128'h4301bfd900d7002307850006c68300f5, /* 1365 */
128'h06100693430540a0053be68100055663, /* 1366 */
128'h385986ba4e250ff6f81304100693c219, /* 1367 */
128'h04ae6a630ff5761302b8f53b0005089b, /* 1368 */
128'hd53bfec68fa306850ff676130306061b, /* 1369 */
128'h0300059340e0063b8536fcb8ffe302b8, /* 1370 */
128'h02d007930003076302f6e96300a606bb, /* 1371 */
128'h0015559b9d1900050023050500f50023, /* 1372 */
128'h808200b7ea630006879bfff5081b4681, /* 1373 */
128'h07bbb7d1feb50fa30505bf4500c8063b, /* 1374 */
128'h0007c30300d7063397ba9381178240f8, /* 1375 */
128'hb7e10117802300660023068500064883, /* 1376 */
128'he8d2eccef4a6f8a2597d011cf0ca7119, /* 1377 */
128'hf02ef42afc3e843684b2e0dafc86e4d6, /* 1378 */
128'h591303000a9306c00a1302500993f82a, /* 1379 */
128'h079bc52d8f1d0004c50377a277420209, /* 1380 */
128'h0135086304d7ff639381178276820017, /* 1381 */
128'h0014c503bfe1e71ff0ef020103930485, /* 1382 */
128'h0004c783035510634781048905450f63, /* 1383 */
128'h00f6f36346a50ff7f793fd07879bcb9d, /* 1384 */
128'h06d50f630640069304890014c5034781, /* 1385 */
128'h0630079304d50f630580069302a6eb63, /* 1386 */
128'h69e6790674a6744670e6f55d08f50963, /* 1387 */
128'hc503808261090007051b6b066aa66a46, /* 1388 */
128'h6c6306e50e6307300713b74d048d0024, /* 1389 */
128'h003800840b13f6e51ee30700071300a7, /* 1390 */
128'h071302e5006307500713a00d46014685, /* 1391 */
128'h003800840b13fa850613f6e510e30780, /* 1392 */
128'h0b13f8b50693a81145c1001636134685, /* 1393 */
128'hf0ef400845a946010016b69300380084, /* 1394 */
128'hdd1ff0ef0028020103930005059be31f, /* 1395 */
128'hf0ef00840b130201039300044503a809, /* 1396 */
128'h01247433600000840b13b5fd845ad89f, /* 1397 */
128'h8522020103930005059b501010ef8522, /* 1398 */
128'he0c2fc3ef83aec061034f436715db7f1, /* 1399 */
128'h715d8082616160e2e8dff0efe436e4c6, /* 1400 */
128'hf83aec06100005931014862ef436f032, /* 1401 */
128'h616160e2e69ff0efe436e4c6e0c2fc3e, /* 1402 */
128'h05931234862afe36fa32f62e710d8082, /* 1403 */
128'heec6eac2e6bee2baea22ee0608081000, /* 1404 */
128'h8522157020ef0808842ae3fff0efe436, /* 1405 */
128'h0087b303679c691c80826135645260f2, /* 1406 */
128'h04b7ec63479d80824501830200030363, /* 1407 */
128'h431c9736002597136b06869300004697, /* 1408 */
128'h2483795c878297b6e426e822ec061101, /* 1409 */
128'h54330e7010ef908114827540f55c08c5, /* 1410 */
128'h8082610545016442e90064a260e20294, /* 1411 */
128'h95aa058e05e135f1bfe1617cbff17d5c, /* 1412 */
128'he02211418082557d8082557db7f1659c, /* 1413 */
128'h679c681c00055e63ff5ff0ef842ae406, /* 1414 */
128'h014160a264028522000307630207b303, /* 1415 */
128'h8082557d80820141640260a245018302, /* 1416 */
128'h6487879300004797150200a7eb6347ad, /* 1417 */
128'h8c8505130000651780826108953e8175, /* 1418 */
128'h47a1715d83020007b303679c691c8082, /* 1419 */
128'he42e078517824785d23e47d502f11023, /* 1420 */
128'hcc3ed402e486100c200007930030e83e, /* 1421 */
128'h400407374d148082616160a6fd3ff0ef, /* 1422 */
128'h01f1041322813823dc01011308e6e063, /* 1423 */
128'h1a05348322113c232291342385a29801, /* 1424 */
128'h0d630a0447830a04c703e909fadff0ef, /* 1425 */
128'h34832301340323813083fb60051300f7, /* 1426 */
128'h0dd447830dd4c7038082240101132281, /* 1427 */
128'hfcf71be30c0447830c04c703fef711e3, /* 1428 */
128'h05934611fcf715e30e0447830e04c703, /* 1429 */
128'hbf654501fd4559b010ef0d4485130d44, /* 1430 */
128'hf4063e800513842af022717980824501, /* 1431 */
128'hc40200011023858a4601852271c020ef, /* 1432 */
128'h20ef7d000513e509842af21ff0efc202, /* 1433 */
128'h4785717980826145740270a285226fe0, /* 1434 */
128'h842ac402c23ef406f022478500f11023, /* 1435 */
128'hf80686934bdc008006b74538691cc195, /* 1436 */
128'h400007378fd98f75600006b78ff58ff9, /* 1437 */
128'he119ec9ff0ef8522858a4601c43e8fd9, /* 1438 */
128'h47b5711d80826145740270a2c43c47b2, /* 1439 */
128'hfc4ee0ca07c55783c23e47d500f11023, /* 1440 */
128'he8a26a056989fdf949370107979bf852, /* 1441 */
128'h4495c43e842e8b2af456ec86f05ae4a6, /* 1442 */
128'h858a4601e00a0a13e009899308090913, /* 1443 */
128'hc7891005f79345b2ed15e71ff0ef855a, /* 1444 */
128'h5517c7950125f7b3054795630135f7b3, /* 1445 */
128'h60e6fba00513d4dff0ef722505130000, /* 1446 */
128'h61257b027aa27a4279e2690664a66446, /* 1447 */
128'h00805863fff40a9bfe04c5e334fd8082, /* 1448 */
128'h45018456b74d8456608020ef3e800513, /* 1449 */
128'hd07ff0ef6f45051300005517fc8047e3, /* 1450 */
128'h47c17139e7a919c52783bf6df9200513, /* 1451 */
128'hfc06f822858a460147d5c42e00f11023, /* 1452 */
128'h1b842783c11ddddff0efc23e842af426, /* 1453 */
128'hdc7ff0ef8522858a46014495cb918b89, /* 1454 */
128'h8082612174a2744270e2f8ed34fdc901, /* 1455 */
128'hec86e0cae4a6711d80824501bfd54501, /* 1456 */
128'h270347c906d7f66384b6892a4785e8a2, /* 1457 */
128'hd432cf3108c92783260102f1102302c9, /* 1458 */
128'hd23a854a100c47850030cc3ee42e4755, /* 1459 */
128'hf0634785e529842ad6fff0efc83eca26, /* 1460 */
128'h854a100c47f5460102f1102347b10497, /* 1461 */
128'h051300005517c11dd4fff0efd23ed402, /* 1462 */
128'h690664a6644660e68522c41ff0ef64e5, /* 1463 */
128'h841bb74d02f6063bbf6147c580826125, /* 1464 */
128'hf426f822fc067139b7c54401b7d50004, /* 1465 */
128'h8a2e4148842ace05e456e852ec4ef04a, /* 1466 */
128'h00b44583c11d892a4a4010ef8ab684b2, /* 1467 */
128'h014485b3681000054d638b3fa0ef8522, /* 1468 */
128'hbd7ff0ef604505130000551700b67a63, /* 1469 */
128'hf96decdff0ef854a08c92583a0894481, /* 1470 */
128'h844e0089f3630207e4030109378389a6, /* 1471 */
128'hfc851ae3f01ff0ef854a85d6865286a2, /* 1472 */
128'h9aa2028784339a22408989b308c96783, /* 1473 */
128'h69e274a279028526744270e2fc0999e3, /* 1474 */
128'h0106161b0086969b808261216aa26a42, /* 1475 */
128'h8e5500f11023030006b78e5547997139, /* 1476 */
128'h440dc432c23e84aafc06f426f82247f5, /* 1477 */
128'h3e800593e919c4dff0ef8526858a4601, /* 1478 */
128'h8082612174a2744270e2d8bff0ef8526, /* 1479 */
128'hbffc07b7db0101134d18bfcdfc79347d, /* 1480 */
128'h3c2324813023241134239fb923213823, /* 1481 */
128'h1ce7f36349013ffc0737233134232291, /* 1482 */
128'h892ac03ff0ef84aa85a2980101f10413, /* 1483 */
128'h20ef20000513e7991a04b7831e051a63, /* 1484 */
128'h06131e0505631a04b5031aa4b0237920, /* 1485 */
128'h6d6347210c04478313d010ef85a22000, /* 1486 */
128'h53b897ba078a1ee70713000047171cf7, /* 1487 */
128'h278300e7fd63cc981ff78793400407b7, /* 1488 */
128'h73630147d69307a68007071367050d44, /* 1489 */
128'h06f48f2309b449830a044783f8dc00d7, /* 1490 */
128'h4783c7890e244783e7810019f9938b85, /* 1491 */
128'h8b890a04478300098a6308f480a30b34, /* 1492 */
128'h07130e24478306f48fa309c44783c789, /* 1493 */
128'h05130a844783fcdc07c60c8486130914, /* 1494 */
128'h00074583fff74783e0fc07c6468109d4, /* 1495 */
128'h97aeffe745839fad0105959b0087979b, /* 1496 */
128'h02f585b30e04458300098c634685c391, /* 1497 */
128'h0621070de21c07ce02b787b30dd44783, /* 1498 */
128'h08d4470308e4478304098f63fce514e3, /* 1499 */
128'h08c447039fb90087171b0107979b4685, /* 1500 */
128'h87b30dd4478302f707330e04470397ba, /* 1501 */
128'h979b08a4470308b44783f8fc07ce02e7, /* 1502 */
128'h0087171b089447039fb90107171b0187, /* 1503 */
128'h07a6c319f4fc54d89fb9088447039fb9, /* 1504 */
128'h8bfd09c44783c7898b850a044783f4fc, /* 1505 */
128'hf0ef852645850af006134685c6b5e391, /* 1506 */
128'h979b0e0447830af407a34785e141e0bf, /* 1507 */
128'h278300098663c79954dc08f4aa2300a7, /* 1508 */
128'h87bb0dd447030e044783f8dc07a60d44, /* 1509 */
128'h80230a74478308f4ac2300a7979b02e7, /* 1510 */
128'h23813483854a240134032481308308f4, /* 1511 */
128'h47838082250101132281398323013903, /* 1512 */
128'h0057d79b00a7d71b50fcf3dd8b850af4, /* 1513 */
128'h08f4aa2302f707bb278527058bfd8b7d, /* 1514 */
128'hb0235f0020efdd4d1a04b503892ab75d, /* 1515 */
128'hdc010113b7655929b7755951bf451a04, /* 1516 */
128'h23213023229134232281382322113c23, /* 1517 */
128'hed8554a9468104b7ec6306f584634789, /* 1518 */
128'h84aad3fff0ef892a45850b900613842e, /* 1519 */
128'h01f10413ed91258199f5ffe4059be11d, /* 1520 */
128'h0b944783e9159a7ff0ef854a85a29801, /* 1521 */
128'h85262301340323813083df400493e399, /* 1522 */
128'h879b8082240101132281348322013903, /* 1523 */
128'h84aab7554685fef760e354a94705ffc5, /* 1524 */
128'h4783f022f406e44ee84aec267179bfd9, /* 1525 */
128'h8edd892e9be10079f6930ff5f9930815, /* 1526 */
128'h57b5c519cc1ff0ef84aa45850b300613, /* 1527 */
128'hf0ef852685ca00091c6300f51e63842a, /* 1528 */
128'h8522013505a317a010ef8526842a86df, /* 1529 */
128'h01138082614569a2694264e2740270a2, /* 1530 */
128'h3023289134232881382328113c23d601, /* 1531 */
128'h3023275134232741382327313c232921, /* 1532 */
128'h3023259134232581382325713c232761, /* 1533 */
128'h07b74d180ac7ed63478923b13c2325a1, /* 1534 */
128'hbfe787933ffc07b79f3dbff7879bbffc, /* 1535 */
128'heb6320250513000055178a2e8b3284aa, /* 1536 */
128'h00005517e7b90016f79307e4c68300e7, /* 1537 */
128'h30838522f8400413f8eff0ef22450513, /* 1538 */
128'h39832801390328813483290134032981, /* 1539 */
128'h3b8326013b0326813a8327013a032781, /* 1540 */
128'h3d8324013d0324813c8325013c032581, /* 1541 */
128'h000055170984a70380822a0101132381, /* 1542 */
128'hf99302f109930045aa83db451fc50513, /* 1543 */
128'h0005ac83e79102eaf7bb060a8063fe09, /* 1544 */
128'hf0ef1fa5051300005517cb8902ecf7bb, /* 1545 */
128'he3994b8502eadabb54dcb7615429f14f, /* 1546 */
128'h47818956866200ca05138c0a009c9c9b, /* 1547 */
128'h02e878bb0017859b0005280343114e05, /* 1548 */
128'hed6ff0ef1f4505130000551700088d63, /* 1549 */
128'h202302e858bbb7f14b814a814c81b7c9, /* 1550 */
128'h8b850107c78397d2078e020800630116, /* 1551 */
128'h893b0ffbfb9300fbebb300be17bbcb89, /* 1552 */
128'h000b8963fa6596e387ae061105210128, /* 1553 */
128'h85ceee068de31d650513000055178a89, /* 1554 */
128'h09f9c603ee051ae3842af8aff0ef8526, /* 1555 */
128'hc7839e3d0087979b0106161b09e9c783, /* 1556 */
128'h05130000551785ca01267a63963e09d9, /* 1557 */
128'h0a79c683008a4783b5c9e50ff0ef1ce5, /* 1558 */
128'hc3990fe6f9138b89c71989360017f713, /* 1559 */
128'h078e0017861b4591450547810016e913, /* 1560 */
128'h00c517bbc39d8b850017579b4b9897d2, /* 1561 */
128'hd79b8b050189191b0187979b0027571b, /* 1562 */
128'h0ff979130127e933c70d4189591b4187, /* 1563 */
128'h8b850a69c78302d90263fcb614e387b2, /* 1564 */
128'hb5a939c020ef1865051300005517ef89, /* 1565 */
128'h8b8509b9c783bfd100f97933fff7c793, /* 1566 */
128'h547ddb8ff0ef1b65051300005517cb89, /* 1567 */
128'h4685e3958b850af9c783e20b05e3b535, /* 1568 */
128'h4785e579a21ff0ef852645850af00613, /* 1569 */
128'h08f4aa2300a7979b0e09c7830af987a3, /* 1570 */
128'hf88d061b00dcd6bb003d169b4d914d01, /* 1571 */
128'h9edff0ef852645850ff676130ff6f693, /* 1572 */
128'h003a169b4c8dfdbd1fe32d05e9458a2a, /* 1573 */
128'h0ff676130ff6f693f8ca061b00dad6bb, /* 1574 */
128'hff9a10e32a05e92d9c5ff0ef85264585, /* 1575 */
128'h26834c818ad209b00d934d6108f00a13, /* 1576 */
128'h85260ff6f6930196d6bb45858656000c, /* 1577 */
128'h90e30ffafa932ca12a85e139999ff0ef, /* 1578 */
128'h86defdba18e30c110ffa7a132a0dffac, /* 1579 */
128'h4785ed19971ff0ef8526458509c00613, /* 1580 */
128'h0613468501279b630a79c783d4fb0ee3, /* 1581 */
128'h86cab381842a953ff0ef8526458509b0, /* 1582 */
128'hdd79842a941ff0ef852645850a700613, /* 1583 */
128'he0ef842ae406e0221141b325842ab335, /* 1584 */
128'h07630187b303679c681c00055e63ffdf, /* 1585 */
128'h60a245058302014160a2640285220003, /* 1586 */
128'hf04af822fc06f4267139808201416402, /* 1587 */
128'h04f592635529478500f5866384aa4791, /* 1588 */
128'h4955842e07c4d78300f1102303700793, /* 1589 */
128'hf0efc43ec24a8526858a46010107979b, /* 1590 */
128'h1f634791c24a00f110234799ed19d44f, /* 1591 */
128'hd26ff0ef8526858a4601c43e478900f4, /* 1592 */
128'h14e3478580826121790274a2744270e2, /* 1593 */
128'h0007869b4f5c6918e215b7cdc402fef4, /* 1594 */
128'h0007069b0007859b4f1887ae00d5f363, /* 1595 */
128'h02c50823dd0c0007859b87ba00d5f363, /* 1596 */
128'h711910000737691c80828082c18ff06f, /* 1597 */
128'he8d2eccef0caf4a6fc86f8a2070d4b9c, /* 1598 */
128'h842ac17c8fd9f466f862fc5ee0dae4d6, /* 1599 */
128'h2423eb8d6b9c679c681cc509f07ff0ef, /* 1600 */
128'h0493b98ff0effb650513000055170204, /* 1601 */
128'h6a4669e674a679068526744670e6f850, /* 1602 */
128'h541c808261097ca27c427be26b066aa6, /* 1603 */
128'h47851af42c23478df93ff0eff3e54481, /* 1604 */
128'h0513b8eff0ef852202042c2302f40823, /* 1605 */
128'h97826b9c679c8522681c43b010ef7d00, /* 1606 */
128'h1a04282318042e2308842783f94584aa, /* 1607 */
128'h4601b5eff0ef8522d85c478508f42223, /* 1608 */
128'h84aacdaff0ef8522f13ff0ef85224581, /* 1609 */
128'h102347a1000505a346d000ef8522f149, /* 1610 */
128'h1aa007138ff94bdc00ff8737681c00f1, /* 1611 */
128'hc43a8522858a460147d50aa00713e399, /* 1612 */
128'h0aa0079300c14703e911be0ff0efc23e, /* 1613 */
128'h09933e900913cc1c800207b700f71563, /* 1614 */
128'h0c3700ff8bb74b0502900a934a550370, /* 1615 */
128'h013110238522858a460140000cb78002, /* 1616 */
128'h10234c18681ce13db9eff0efc402c252, /* 1617 */
128'h01871563c43e0177f7b3c25a4bdc0151, /* 1618 */
128'hb76ff0ef8522858a4601c43e0197e7b3, /* 1619 */
128'h051306090863397d0007ca6347b2ed1d, /* 1620 */
128'h8563800207374c14bf4534b010ef3e80, /* 1621 */
128'h8b8541e7d79bc43ccc188001073700e6, /* 1622 */
128'h0793b55d18f40ca3478506041e23d45c, /* 1623 */
128'h85224581becff0ef852202f51f63f920, /* 1624 */
128'h0c2347850007d663443ced09c1cff0ef, /* 1625 */
128'h5517d965c04ff0ef85224585bfd118f4, /* 1626 */
128'hb595fa1004939fcff0efe32505130000, /* 1627 */
128'heb4aef26f706f3227161551cb58584aa, /* 1628 */
128'heaeaeee6f2e2f6defadafed6e352e74e, /* 1629 */
128'hc783219010ef45018baae3b54401e6ee, /* 1630 */
128'h4789e7b5180b8ca3198bc783c7b1199b, /* 1631 */
128'hc482c2be855e008c479d460104f11023, /* 1632 */
128'h8b851b8ba78312050ae3842aaa2ff0ef, /* 1633 */
128'h842aa88ff0ef855e008c46014495cf81, /* 1634 */
128'h855ea031020ba423f4fd34fd10050de3, /* 1635 */
128'h64fa741a70ba8522d55d842ad99ff0ef, /* 1636 */
128'h6cf67c167bb67b567af66a1a69ba695a, /* 1637 */
128'h180b8c23048ba7838082615d6db66d56, /* 1638 */
128'h187010ef4501afeff0ef855e0407c163, /* 1639 */
128'hf0ef855e45853e800913908102051493, /* 1640 */
128'h85260007cc63048ba783f155842ab1ef, /* 1641 */
128'h1f1010ef0640051308a96fe3163010ef, /* 1642 */
128'hd79b048ba78300fbac23400007b7bfe9, /* 1643 */
128'hbf0506fb9e23478502fba6238b8541e7, /* 1644 */
128'h071b40010737a0292007071b40010737, /* 1645 */
128'h00003a178a1d0036571b00ebac234007, /* 1646 */
128'h1086260396529752060a8b3d7f4a0a13, /* 1647 */
128'hd61b02c7073b018ba88345050f874703, /* 1648 */
128'h04cba823180bae231a0ba8238a0500c7, /* 1649 */
128'h183b8b3d0107d71b08eba22308eba423, /* 1650 */
128'ha703090ba8231408dd63090ba62300e5, /* 1651 */
128'h8f7d003f07370107979b14070f6302cb, /* 1652 */
128'h00d797b32689078546a18fd90106d79b, /* 1653 */
128'h0c0bb4230c0bb0230a0bbc23030787b3, /* 1654 */
128'h0afbb8230e0bb0230c0bbc230c0bb823, /* 1655 */
128'h090ba70308fba6230107d46320000793, /* 1656 */
128'ha783c21508fba82300e7f46320000793, /* 1657 */
128'h46010107979b471100e78e63577d04cb, /* 1658 */
128'h8f6ff0efc282c4be04e11023855e008c, /* 1659 */
128'h979b4601495507cbd78304f11023479d, /* 1660 */
128'h842a8d8ff0efc4bec2ca855e008c0107, /* 1661 */
128'h08fb80a357fd08fbaa234785e4051ce3, /* 1662 */
128'h00ef855ee40510e3842ac94ff0ef855e, /* 1663 */
128'h15e3842aff3fe0ef855e00b545831130, /* 1664 */
128'h2789100007b754075963018ba703e205, /* 1665 */
128'h07cbd78306f110230370079304fba023, /* 1666 */
128'hf0efd4bed2ca855e0107979b108c4601, /* 1667 */
128'h033007930bf104934905d2caed05874f, /* 1668 */
128'h0a854991d48206f11023988102091a93, /* 1669 */
128'hf0efd05aec56e826855e108c08104b21, /* 1670 */
128'h0737bb75842afe0996e339fdc529844f, /* 1671 */
128'hbd9140040737bda940030737bd894002, /* 1672 */
128'hb54508bba82300b515bb89bd0165d59b, /* 1673 */
128'h8fd901e6d71b8ff90027979b17716705, /* 1674 */
128'h05374098bd798a9d938100f6d69b1782, /* 1675 */
128'h8fd50087161b0187179b0187569b00ff, /* 1676 */
128'h8ef1f00706138fd167410087569b8e69, /* 1677 */
128'h169b0187559b40d804fbaa2327818fd5, /* 1678 */
128'h8ecd0087571b8de90087159b8ecd0187, /* 1679 */
128'h0d638b3d0187d71b04ebac238f558f71, /* 1680 */
128'hac238001073708d70e634689c7010927, /* 1681 */
128'h0737040ba7830007596302d7971300eb, /* 1682 */
128'h800107b7018ba70304fba0238fd92000, /* 1683 */
128'ha903639c21c787930000579708f71363, /* 1684 */
128'h00003497044ba783f0be0ff10c13040b, /* 1685 */
128'h9a93478500f97933fe0c7c9360c48493, /* 1686 */
128'h00e797bb478540980a8583f979130207, /* 1687 */
128'h87930000379704a1ebc5278100f977b3, /* 1688 */
128'he0efa7a5051300005517fef493e35ee7, /* 1689 */
128'ha007071b80011737b949df400413e15f, /* 1690 */
128'hb785800207370007456303079713b7bd, /* 1691 */
128'h01000ab70ff104934905bfa980030737, /* 1692 */
128'h0209886339fd09053ac5499598811902, /* 1693 */
128'h040007931030c33e47d508f110234799, /* 1694 */
128'heb7fe0efdc3ef84af426c556855e010c, /* 1695 */
128'h674144dcfbe18b8583a54cdce6051de3, /* 1696 */
128'h8fd58ff90087d79b0087969bf0070713, /* 1697 */
128'h0087e793040ba783f20750e302e79713, /* 1698 */
128'h0b1b06010993017d8b37bf0104fba023, /* 1699 */
128'h01a7f7b300f977b30009ad0340dc840b, /* 1700 */
128'h00fd0d6345a1400007b712078e632781, /* 1701 */
128'h05b3100005b700fd08634591200007b7, /* 1702 */
128'h19638daa8bfff0ef855e0015b59340bd, /* 1703 */
128'h2000073700ed0d6347a1400007370e05, /* 1704 */
128'h379340fd0d33100007b700ed08634791, /* 1705 */
128'h4705409cd41fe0ef855e02fbaa23001d, /* 1706 */
128'h102347994d850ae79d63470d00e78663, /* 1707 */
128'he7b317c12d81810007b7d33e47d50af1, /* 1708 */
128'he166855e110c040007930110d53e00fd, /* 1709 */
128'h8bbd010cc783e541dcffe0efc93ee556, /* 1710 */
128'h088ba583efd91afba823409c09b79063, /* 1711 */
128'h460118fbae2308bba2230017b79317ed, /* 1712 */
128'hd7830af1102303700793895ff0ef855e, /* 1713 */
128'hd33a855e110c0107979b4601475507cb, /* 1714 */
128'h7d1347b56702ed05d7ffe0efd53ee03a, /* 1715 */
128'h07134791d5028dead33a0af11023fe0c, /* 1716 */
128'hc93ae556e16ae43e855e110c01100400, /* 1717 */
128'hf3f537fd670267a2c521d51fe0efe03a, /* 1718 */
128'hae23096ba2231afba823017d85b74785, /* 1719 */
128'h099181dff0ef855e840585934601180b, /* 1720 */
128'hf6f762e34581472db575def98be310bc, /* 1721 */
128'h66c1bf91118725839752837902079713, /* 1722 */
128'h000d2783f006869300ff0537040d0593, /* 1723 */
128'h0087961b8f510187971b0187d61b0d11, /* 1724 */
128'hfefd2e238fd98ff58f510087d79b8e69, /* 1725 */
128'h8bbd00c7579b46a5008da703fda59ee3, /* 1726 */
128'h04d61c63800306b7018ba60300f6f863, /* 1727 */
128'h1487a78397b6078a2e06869300003697, /* 1728 */
128'h17fd67c100cda68308fbae230087171b, /* 1729 */
128'h0126d71bc78d27818fd18ff90186d61b, /* 1730 */
128'hd69b02e6073b3e800613c30503f77713, /* 1731 */
128'h0afba02302d606bb02f757bb8a8d0106, /* 1732 */
128'h19cba7831afbaa231b0ba7830adba223, /* 1733 */
128'h855e08fba82308fba62320000793c799, /* 1734 */
128'h08cba70300050623000515234a0000ef, /* 1735 */
128'hccc68693aaa78793ccccd6b7aaaab7b7, /* 1736 */
128'h00f037b3068600d036b327818ef98ff9, /* 1737 */
128'h00d036b38ef90f068693f0f0f6b79fb5, /* 1738 */
128'h36b38ef9f0068693ff0106b79fb5068a, /* 1739 */
128'h37338f750207161376c19fb5068e00d0, /* 1740 */
128'hed1092010a8bb783d11c9fb9071200e0, /* 1741 */
128'h06fbc603074bd68307abd70302c7d7b3, /* 1742 */
128'h362302450513756585930000459784aa, /* 1743 */
128'hc603077bc883070ba683a8dfe0effef5, /* 1744 */
128'hf7930ff6f8130106d71b0086d79b06cb, /* 1745 */
128'h8593000045970186d69b0ff777130ff7, /* 1746 */
128'h4597074ba603a59fe0ef04d485137365, /* 1747 */
128'h561b0106569b06248513732585930000, /* 1748 */
128'h00d010ef8526a39fe0ef8a3d8abd0146, /* 1749 */
128'ha0232785100007b7b0cd02fba4234785, /* 1750 */
128'h07b700f778631a0bb603400407b704fb, /* 1751 */
128'h00004517e611b5f1e225ecf769e34004, /* 1752 */
128'ha0230016879b700006b7b1296a450513, /* 1753 */
128'hf5931abba42303f7f5930c46478304fb, /* 1754 */
128'ha0230216869bc58900c7f593cd910027, /* 1755 */
128'h8b8504dba0230106e693040ba68304db, /* 1756 */
128'h07b704fba02300c7e793040ba783d7dd, /* 1757 */
128'ha583044ba783040ba983e6f769e34004, /* 1758 */
128'hdaaff0ef2981855e00f9f9b34601088b, /* 1759 */
128'h0b1300003b174a851784849300003497, /* 1760 */
128'h97bb409c1c0c8c9300003c974c2d18eb, /* 1761 */
128'hff6498e304a1eb99278100f9f7b300fa, /* 1762 */
128'h3917bd2197bfe0ef5e05051300004517, /* 1763 */
128'h409c10000db720000d3715a909130000, /* 1764 */
128'h40dc04f719630017b79317ed00494703, /* 1765 */
128'h4683c3a127818ff900f9f7b300092703, /* 1766 */
128'he0ef855e0fb6f69345850b7006130089, /* 1767 */
128'he0ef855e45850b7006134681c90ddbbf, /* 1768 */
128'ha223180bae231a0ba823088ba783dabf, /* 1769 */
128'h10e30931941fe0ef855e035baa2308fb, /* 1770 */
128'h89634721400006b700092783bfa5fb99, /* 1771 */
128'h0017b71341b787b301a78663471100d7, /* 1772 */
128'he0ef855e408c913fe0ef855e02ebaa23, /* 1773 */
128'h409ce79d0046f79300892683f14dfeff, /* 1774 */
128'h0017b79317ed088ba583ef8d1afba823, /* 1775 */
128'hc9aff0ef855e460118fbae2308bba223, /* 1776 */
128'h06130ff6f693bb35f53d9d9fe0ef855e, /* 1777 */
128'h4581bfa1d171d13fe0ef855e45850b70, /* 1778 */
128'h118725839752837902079713fcfc65e3, /* 1779 */
128'h851300ec4641ef2ff06ffa100413bf6d, /* 1780 */
128'h07cbd78304f11023478d6ce000ef06cb, /* 1781 */
128'hc2be47d5855ec4be0107979b008c4601, /* 1782 */
128'hd663018ba783ec051163842a943fe0ef, /* 1783 */
128'h04f1102347a506fb9e2304e157830007, /* 1784 */
128'h0107979b008c460107cbd783c2be479d, /* 1785 */
128'h4636e8051763842a90ffe0efc4be855e, /* 1786 */
128'ha02304cbae23018ba50345e646d647c6, /* 1787 */
128'h1c634000073706bba42306dba22306fb, /* 1788 */
128'h450d0007081b377d8b3d01a6571bf0e5, /* 1789 */
128'h8379eea50513000035171702ef056863, /* 1790 */
128'h557d80824501c56c8702972a4318972a, /* 1791 */
128'h00005797808218b50d238082557d8082, /* 1792 */
128'he406e02247851141ef9d439cda878793, /* 1793 */
128'h852212a000efd8f7292300005717842a, /* 1794 */
128'h0513fc5ff0ef852200055563ac0fe0ef, /* 1795 */
128'h4501640260a20dc000ef13e000ef02c0, /* 1796 */
128'hd6070713000057178082450180820141, /* 1797 */
128'h0000451785aa114102e790636394631c, /* 1798 */
128'h853e478160a2f3cfe0efe40651450513, /* 1799 */
128'hbfd187b600a604630fc7a60380820141, /* 1800 */
128'hfbdff0efe42eec06110141488082853e, /* 1801 */
128'h0815470302b7006365a210354703c105, /* 1802 */
128'he97fe06f610560e200f70c630ff00793, /* 1803 */
128'hf8400513bfe545018082610560e25535, /* 1804 */
128'hf7dff0ef84aee822ec06e4261101bfcd, /* 1805 */
128'he0800f840413e501ce0ff0ef842acd09, /* 1806 */
128'h5797bfd555358082610564a2644260e2, /* 1807 */
128'h8082c3980015071b4388b02787930000, /* 1808 */
128'h4388aea787930000579780820f850513, /* 1809 */
128'h6380e822c94787930000579711018082, /* 1810 */
128'h64a2644260e20094176384beec06e426, /* 1811 */
128'ha8cff0ef8522c78119a4478380826105, /* 1812 */
128'he79ce39cc647879300005797b7d56000, /* 1813 */
128'h00005797e5088082aa07a02300005797, /* 1814 */
128'h8082e308e518e11ce7886798c4c78793, /* 1815 */
128'h6080e8a2c344849300005497e4a6711d, /* 1816 */
128'he06ae466e862ec5ef05af456f852fc4e, /* 1817 */
128'h4a973faa0a1300004a1789aae0caec86, /* 1818 */
128'h4b973fab0b1300004b173faa8a930000, /* 1819 */
128'h8c9300004c9700050c1b3fab8b930000, /* 1820 */
128'h690664a660e66446029415634d299dec, /* 1821 */
128'h6d026ca26c426be27b027aa27a4279e2, /* 1822 */
128'h541cdb8fe06f61255485051300004517, /* 1823 */
128'h681c89560007c36389524c1cc7914901, /* 1824 */
128'h00090663d9afe0ef638c855a0fc42603, /* 1825 */
128'h85e200978e63601cd8efe0ef855e85ca, /* 1826 */
128'h05130000451701a98863d80fe0ef8566, /* 1827 */
128'hec06e8221101b7716000334010ef9665, /* 1828 */
128'h4d5ccfad44014d1cc1414401e04ae426, /* 1829 */
128'h892ec7ad639cc7bd651ccbad511ccbbd, /* 1830 */
128'hcd21842a20a010ef45051c00059384aa, /* 1831 */
128'h10f502a347850ef52c234799c57c57fd, /* 1832 */
128'hf797e65ff0ef0405282303253023e904, /* 1833 */
128'h87930000179716f43c238fa78793ffff, /* 1834 */
128'h34232b8787930000179718f430232c87, /* 1835 */
128'h00230247c78385220ea42e23681c18f4, /* 1836 */
128'h690264a2644260e28522e99ff0ef10f4, /* 1837 */
128'h88068693000056971c60106f80826105, /* 1838 */
128'h97360017671302d786b365186294611c, /* 1839 */
128'h00f7553b93ed836d8f3d0127d713e118, /* 1840 */
128'h5517808225018d5d00f717bb40f007bb, /* 1841 */
128'he022e4061141fc3ff06faaa505130000, /* 1842 */
128'h8d410105151bfe9ff0ef842afefff0ef, /* 1843 */
128'he022e4061141808201412501640260a2, /* 1844 */
128'h9001fd1ff0ef14020005041bfdbff0ef, /* 1845 */
128'h058587aa80820141640260a28d411502, /* 1846 */
128'h47818082fb75fee78fa30785fff5c703, /* 1847 */
128'h00f506b30007470300f5873300c78c63, /* 1848 */
128'h0007c70387aa8082f76d00e680230785, /* 1849 */
128'h8fa30785fff5c7030585eb0900178693, /* 1850 */
128'h8082e21987aab7d587b68082fb75fee7, /* 1851 */
128'h0585963efb7d001786930007c70387b6, /* 1852 */
128'hfec799e3d375fee78fa30785fff5c703, /* 1853 */
128'hfff5c783000547030585808200078023, /* 1854 */
128'h0505e3994187d79b0187979b40f707bb, /* 1855 */
128'ha015478100e6146347018082853ef37d, /* 1856 */
128'h0007c78300e587b30007c68300e507b3, /* 1857 */
128'h0705e3994187d79b0187979b40f687bb, /* 1858 */
128'h9363000547830ff5f5938082853efee1, /* 1859 */
128'hf59380824501bfcd0505c399808200b7, /* 1860 */
128'h0505dffd808200b79363000547830ff5, /* 1861 */
128'h808240a78533e7010007c70387aabfcd, /* 1862 */
128'hf0efec06842ae42ee8221101bfcd0785, /* 1863 */
128'h8663000547830ff5f593952265a2fe5f, /* 1864 */
128'h6105644260e24501fe857be3157d00b7, /* 1865 */
128'he7010007c70300b7856387aa95aa8082, /* 1866 */
128'h00f507334781b7fd0785808240a78533, /* 1867 */
128'h0705fed60ee38082853eea9900074683, /* 1868 */
128'h4781bfd5872eb7d50785fa7d00074603, /* 1869 */
128'h0863a021872eca890007468300f50733, /* 1870 */
128'h07858082853efa7d00074603070500d6, /* 1871 */
128'hfee68fe380824501eb1900054703b7c5, /* 1872 */
128'hbfd587aeb7e50505fafd0007c6830785, /* 1873 */
128'h5797e519842a84aeec06e426e8221101, /* 1874 */
128'hf0ef85a68522cc1163808aa787930000, /* 1875 */
128'hb72300005797ef8100044783942afa1f, /* 1876 */
128'h8082610564a2644260e2852244018807, /* 1877 */
128'hc78100054783c519f9fff0ef852285a6, /* 1878 */
128'hbfd986a7b12300005797050500050023, /* 1879 */
128'h8526842ac891e822ec066104e4261101, /* 1880 */
128'h60e2e008050500050023c501f73ff0ef, /* 1881 */
128'h00054783c11d8082610564a285266442, /* 1882 */
128'he3110017c703ce810007c68387aacf99, /* 1883 */
128'h4501b7e5078900d780a300e780238082, /* 1884 */
128'h0ff5f69347a1eb0587aa007577138082, /* 1885 */
128'h469d00c508b387aaffed8f5537fd0722, /* 1886 */
128'h87335761003657930106ee6340f88833, /* 1887 */
128'h808200c79763963e963a97aa078e02e7, /* 1888 */
128'hb7f5feb78fa30785bfe9fee7bc2307a1, /* 1889 */
128'h4781eb9d872a8b9d00b567b304b50463, /* 1890 */
128'h00f506b30006b80300f586b3a811471d, /* 1891 */
128'h5793fed765e340f606b30106b02307a1, /* 1892 */
128'h0733963a95be078e02e7873357610036, /* 1893 */
128'hc80300f586b3808200f61363478100f5, /* 1894 */
128'h7179b7e501068023078500f706b30006, /* 1895 */
128'he02ee84af406e432ec26852e842af022, /* 1896 */
128'h64636582892ace1184aa6622dd3ff0ef, /* 1897 */
128'hf75ff0ef944a864a8522fff6091300c5, /* 1898 */
128'h614564e269428526740270a200040023, /* 1899 */
128'hf0ef00a5e963842ae406e02211418082, /* 1900 */
128'h86ae883280820141640260a28522f53f, /* 1901 */
128'h00f80733fef605e317fd4781fff64613, /* 1902 */
128'hb7e500b7002397220005c58300e685b3, /* 1903 */
128'h86b300e507b3a821478100e614634701, /* 1904 */
128'hd3f59f9507050006c6830007c78300e5, /* 1905 */
128'h00054783808200c51363962a8082853e, /* 1906 */
128'h852e842af0227179bfc50505feb78de3, /* 1907 */
128'h049bd19ff0ef892ee44ef406e84aec26, /* 1908 */
128'h87bb008509bbd0dff0ef8522c8990005, /* 1909 */
128'h64e2740270a2852244010097db634089, /* 1910 */
128'hf0ef852285ca86268082614569a26942, /* 1911 */
128'h14630ff5f593962abfe10405d17df83f, /* 1912 */
128'h0be300150793000547038082450100c5, /* 1913 */
128'h00c7ef630ff5f59347c1b7ed853efeb7, /* 1914 */
128'h0007c7038082853e4781e60187aa2601, /* 1915 */
128'hc39d00757793b7f5367d0785feb71ce3, /* 1916 */
128'h9de30007c68387aa00a7083b9f1d4721, /* 1917 */
128'h93011702fed819e30007869b0785fcb6, /* 1918 */
128'h0107179300b7e733008597938e19953a, /* 1919 */
128'h87aa27018edd00365713020796938fd9, /* 1920 */
128'h0785f8b71fe30007c703d24d8a1deb11, /* 1921 */
128'h00d80a63008785130007b803bfcd367d, /* 1922 */
128'hbfa5fef51be30785f8b712e30007c703, /* 1923 */
128'h079300054703e7c9419cb7f1377d87aa, /* 1924 */
128'h8793000027970015470306f71e630300, /* 1925 */
128'h071bc6898a850006c68300e786b32a67, /* 1926 */
128'h470304d71763078006930ff777130207, /* 1927 */
128'h47c1cf950447f7930007c78397ba0025, /* 1928 */
128'h478302f71f630300079300054703c19c, /* 1929 */
128'h00074703973e25e70713000027170015, /* 1930 */
128'h078007130ff7f7930207879bc7098b05, /* 1931 */
128'h47a98082c19c47a1a809050900e79c63, /* 1932 */
128'h842ee82211018082fae78fe34741bfed, /* 1933 */
128'h468100c16583f61ff0efc632ec06006c, /* 1934 */
128'h0007079b000547032108081300002817, /* 1935 */
128'h00089863044678930006460300f80633, /* 1936 */
128'h00467893808261058536644260e2ec05, /* 1937 */
128'h02d586b3feb7f4e3fd07879b00088b63, /* 1938 */
128'hf793fe07079bc6098a09b7d196be0505, /* 1939 */
128'hf8227139b7e1e008b7cdfc97879b0ff7, /* 1940 */
128'h84b2842ae42e00063023f04afc06f426, /* 1941 */
128'h74a2744270e25529e90165a2b03ff0ef, /* 1942 */
128'hf0ef8522082c892a862e808261217902, /* 1943 */
128'h8f81cb010007c703fe8782e367e2f5df, /* 1944 */
128'h4501e088fcf718e347a9fd279be30785, /* 1945 */
128'hf06f00e6846302d0071300054683b7e9, /* 1946 */
128'h053360a2f23ff0efe40605051141f2df, /* 1947 */
128'hf0ef842ee406e02211418082014140a0, /* 1948 */
128'h02d704630007c70304b00693601cf0df, /* 1949 */
128'h640260a202d70e630470069300e6ea63, /* 1950 */
128'h06b0069302d7076304d0069380820141, /* 1951 */
128'h9fe3052a069007130017c683fed716e3, /* 1952 */
128'h078d00e69863042007130027c683fce6, /* 1953 */
128'h1101bfd50789bff1052a052ab7e9e01c, /* 1954 */
128'h6583e0dff0efc632ec06006c842ee822, /* 1955 */
128'h000547030bc8081300002817468100c1, /* 1956 */
128'h044678930006460300f806330007079b, /* 1957 */
128'h808261058536644260e2ec0500089863, /* 1958 */
128'hfeb7f4e3fd07879b00088b6300467893, /* 1959 */
128'h079bc6098a09b7d196be050502d586b3, /* 1960 */
128'hb7e1e008b7cdfc97879b0ff7f793fe07, /* 1961 */
128'h0693601cf87ff0ef842ee406e0221141, /* 1962 */
128'h069300e6ea6302d704630007c70304b0, /* 1963 */
128'h069380820141640260a202d70e630470, /* 1964 */
128'hc683fed716e306b0069302d7076304d0, /* 1965 */
128'h0027c683fce69fe3052a069007130017, /* 1966 */
128'h052ab7e9e01c078d00e6986304200713, /* 1967 */
128'h842ae406e0221141bfd50789bff1052a, /* 1968 */
128'h2797fff5c70300a405b3951ff0efe589, /* 1969 */
128'h00074703973efff58513fe2787930000, /* 1970 */
128'h157d80820141557d640260a2e7198b11, /* 1971 */
128'h8b1100074703973e00054703fea47ae3, /* 1972 */
128'hf06f014105054581462960a26402f77d, /* 1973 */
128'h8d5d05220085579bfa5ff06f4581d7df, /* 1974 */
128'h87930000479780820141914115421141, /* 1975 */
128'hf06f95be9201160291811582639c4767, /* 1976 */
128'h853ee31900054703462946a54781a93f, /* 1977 */
128'h02f607bb00b6e763fd07059b27018082, /* 1978 */
128'he406e0221141b7c50505fd07879b9fb9, /* 1979 */
128'h55bb45a900b7f86347a500a04563842e, /* 1980 */
128'h640202a4753b4529fe7ff0ef357d02b4, /* 1981 */
128'h081007935020006f03050513014160a2, /* 1982 */
128'h3f23000047173ef73f230000471707e2, /* 1983 */
128'h3f04041300004417e822110180823ef7, /* 1984 */
128'ha05ff0efec06600885aa84ae862ee426, /* 1985 */
128'h8082610564a26442e00c95a660e2600c, /* 1986 */
128'h00004497e4263c678793000047971101, /* 1987 */
128'h0513000045176380e82260903b448493, /* 1988 */
128'h85a26088b5bfd0ef85a29c11ec0697e5, /* 1989 */
128'h051300004517862286aa608ce2dfc0ef, /* 1990 */
128'hd0ef9825051300004517b41fd0ef9765, /* 1991 */
128'h5e63809f90efef85051300000517b35f, /* 1992 */
128'h0000451740a005b364a260e264420005, /* 1993 */
128'h64a260e26442b0dfd06f610597450513, /* 1994 */
128'ha0ef8432e406e022114166a0006f6105, /* 1995 */
128'h0141640260a28522547d00850363822f, /* 1996 */
128'he64e01258413f2227169808245018082, /* 1997 */
128'hf76ff0ef892eea4aee26f606852289aa, /* 1998 */
128'h95260505f6aff0ef852600a404b30505, /* 1999 */
128'h04e7ee631ff00793fff5071be93ff0ef, /* 2000 */
128'h84aaf48ff0ef85222ca7ac2300004797, /* 2001 */
128'h07939526f3aff0ef6e85051300003517, /* 2002 */
128'h3517842af2aff0ef852204a7f2630ff0, /* 2003 */
128'h451700a405b3f1cff0ef6ca505130000, /* 2004 */
128'h64f2741270b2a5dfd0ef8e2505130000, /* 2005 */
128'h00004717200007938082615569b26952, /* 2006 */
128'hf0ef850a458110000613b75526f72e23, /* 2007 */
128'hde0ff0ef850a6865859300003597855f, /* 2008 */
128'h0000459700f7096302f0079301294703, /* 2009 */
128'hf0ef850a85a2df4ff0ef850a8b458593, /* 2010 */
128'h4517858a43902367879300004797decf, /* 2011 */
128'h07e2081007939edfd0ef89a505130000, /* 2012 */
128'h3f230000471720f73f23000047174511, /* 2013 */
128'h4501fea79d2300004797d87ff0ef20f7, /* 2014 */
128'h45974611fea7972300004797d79ff0ef, /* 2015 */
128'h47174785eafff0ef854efe2585930000, /* 2016 */
128'he426ec06e8221101b7911cf71f230000, /* 2017 */
128'h84ae450d892a08c7df638432478de04a, /* 2018 */
128'h451708a7956325010004d783d39ff0ef, /* 2019 */
128'h25010024d783d23ff0ef1ae555030000, /* 2020 */
128'hda9ff0ef00448513ffc4059b06a79a63, /* 2021 */
128'h4517f6a79d2300004797d07ff0ef4511, /* 2022 */
128'h000047974611cf3ff0ef17e555030000, /* 2023 */
128'hf0ef854af5c5859300004597f6a79323, /* 2024 */
128'h1545d58300004597256000ef4535e29f, /* 2025 */
128'h4797240000ef02000513d19ff0ef4515, /* 2026 */
128'h0000471727850007d78313e787930000, /* 2027 */
128'h278d439c124787930000479712f71823, /* 2028 */
128'h8d7fd0ef7a450513000035170087cf63, /* 2029 */
128'h60e2d47ff06f6105690264a260e26442, /* 2030 */
128'hf022f406717980826105690264a26442, /* 2031 */
128'h0f230115c70300e10fa346890105c703, /* 2032 */
128'h02f70a63478d00d70e6301e1570300e1, /* 2033 */
128'hd06f6145784505130000351770a27402, /* 2034 */
128'hd0efe42e75c5051300003517842a885f, /* 2035 */
128'hd8bff06f614570a265a274028522875f, /* 2036 */
128'h0113ebfff06f614505c170a241907402, /* 2037 */
128'h842a232130232291342322813823dc01, /* 2038 */
128'h22113c230028218006134581893284ae, /* 2039 */
128'he802c44a08282040061385a6e52ff0ef, /* 2040 */
128'h23813083f63ff0ef8522002ce90ff0ef, /* 2041 */
128'h24010113220139032281348323013403, /* 2042 */
128'h45974611cb8103a7d783000047978082, /* 2043 */
128'he40611418082cf1ff06fe22585930000, /* 2044 */
128'ha70300e57763878e1041e703504000ef, /* 2045 */
128'h1007e78310a7a22310e1a02327051001, /* 2046 */
128'h4501808201418d5d91011782150260a2, /* 2047 */
128'hfc1ff0ef84aae426e822ec0611018082, /* 2048 */
128'h150202f407b33e800793440000ef842a, /* 2049 */
128'h610564a28d0502a7d533644260e29101, /* 2050 */
128'h00ef842af95ff0efe022e40611418082, /* 2051 */
128'h60a202f407b324078793000f47b74140, /* 2052 */
128'h1101808202a7d5330141910115026402, /* 2053 */
128'h892af63ff0ef84aae04ae426e822ec06, /* 2054 */
128'h24040413000f443702a485333e2000ef, /* 2055 */
128'hfe856ee3f45ff0ef0405944a02855433, /* 2056 */
128'he426110180826105690264a2644260e2, /* 2057 */
128'h68048493842ae04aec06e822009894b7, /* 2058 */
128'hf0ef41240433854a89260084f3638922, /* 2059 */
128'h80826105690264a2644260e2f47dfa1f, /* 2060 */
128'h410007b7808200054503808200b50023, /* 2061 */
128'h4783410007378082020575130147c503, /* 2062 */
128'h07b7808200a70023dfe50207f7930147, /* 2063 */
128'h476d00e78623f8000713000782234100, /* 2064 */
128'h071300e78623470d0007822300e78023, /* 2065 */
128'h808200e788230200071300e78423fc70, /* 2066 */
128'h60a2e50900044503842ae406e0221141, /* 2067 */
128'h2797b7f50405fa5ff0ef808201416402, /* 2068 */
128'h97aa973e811100f57713f1a787930000, /* 2069 */
128'h00f5802300e580a30007c78300074703, /* 2070 */
128'hf0efec068121842a002ce82211018082, /* 2071 */
128'hf0ef00914503f65ff0ef00814503fd1f, /* 2072 */
128'h00814503fb7ff0ef0ff47513002cf5df, /* 2073 */
128'h644260e2f43ff0ef00914503f4bff0ef, /* 2074 */
128'h892af406e84aec26f022717980826105, /* 2075 */
128'hf0ef0ff57513002c0089553b54e14461, /* 2076 */
128'h00914503f13ff0ef346100814503f81f, /* 2077 */
128'h694264e2740270a2fe9410e3f0bff0ef, /* 2078 */
128'h892af406e84aec26f022717980826145, /* 2079 */
128'h0ff57513002c0089553354e103800413, /* 2080 */
128'h4503ed1ff0ef346100814503f3fff0ef, /* 2081 */
128'h64e2740270a2fe9410e3ec9ff0ef0091, /* 2082 */
128'hf13ff0efec06002c1101808261456942, /* 2083 */
128'he9fff0ef00914503ea7ff0ef00814503, /* 2084 */
128'h439cfe278793000047978082610560e2, /* 2085 */
128'h842e892aec4efc06f04af426f8227139, /* 2086 */
128'hb0efd8a505130000451702b7856384b2, /* 2087 */
128'h70e2faa7ab2300004797c10d2501f08f, /* 2088 */
128'h471757fd8082612169e2790274a27442, /* 2089 */
128'h0000451785ca86260074f8f72d230000, /* 2090 */
128'h00004797c50d2501fe3fa0efd5450513, /* 2091 */
128'h0000351785a6049675634632f8a7a023, /* 2092 */
128'h2123000047174785cdefd0ef3fc50513, /* 2093 */
128'h099b00c4591be05ff0ef4521b775f6f7, /* 2094 */
128'h993e003979133f678793000037970009, /* 2095 */
128'hbf5d2f4010ef854ede7ff0ef00094503, /* 2096 */
128'he0221141bf95f287a323000047979c25, /* 2097 */
128'hd0efe4063cc5051300003517842a85aa, /* 2098 */
128'h8322f14025730ff0000f0000100fc84f, /* 2099 */
128'h83020141d7c585930000259760a26402, /* 2100 */
128'h000045170b4585930000359746051141, /* 2101 */
128'hc9112501d47fa0efe022e406ee450513, /* 2102 */
128'hd06f014160a264023b05051300003517, /* 2103 */
128'h4605c28fd0ef3be5051300003517c34f, /* 2104 */
128'hc6850513000045173d05859300003597, /* 2105 */
128'h3c85051300003517c5112501d69fa0ef, /* 2106 */
128'h0517bf8fd0ef2465051300003517b7e1, /* 2107 */
128'h4797e607ab2300004797e98505130000, /* 2108 */
128'h00054863842a8bcf90efe607a5230000, /* 2109 */
128'h408005b3cf81439ce5c7879300004797, /* 2110 */
128'hd06f014121c505130000351760a26402, /* 2111 */
128'h2501b72fb0efbfe5051300004517bb4f, /* 2112 */
128'h35974605bfb93765051300003517c511, /* 2113 */
128'hc5112501c87fa0ef4501fea585930000, /* 2114 */
128'hee1ff0ef8522b7813705051300003517, /* 2115 */
128'hd69ff0efe40625011141900200000023, /* 2116 */
128'h80824501808224050513000f4537a001, /* 2117 */
128'h00756513157d631cdd07071300004717, /* 2118 */
128'h953e055e10d00513e308953600178693, /* 2119 */
128'he4328532ec06e822110102b506338082, /* 2120 */
128'h936ff0ef45816622c509842afd1ff0ef, /* 2121 */
128'h35171141808280826105644260e28522, /* 2122 */
128'h42000537afafd0efe40630a505130000, /* 2123 */
128'h8082450180820141450160a2eadfc0ef, /* 2124 */
128'h808202f5553347a9b000257380824501, /* 2125 */
128'h05130000351785aa862e86b287361141, /* 2126 */
128'ha001cbbff0ef4505abefd0efe4062f65, /* 2127 */
128'h07b3f57ff0efe406952e842ae0221141, /* 2128 */
128'h4505808201418d7d640260a295224080, /* 2129 */
128'hec26f022717980824505808245058082, /* 2130 */
128'h740270a20096186300c684bb842ef406, /* 2131 */
128'hc0efe432852285b280826145450164e2, /* 2132 */
128'h80824509bff92605200404136622dfff, /* 2133 */
128'h45018082808280828082450980824509, /* 2134 */
128'he822ec061101bbbff06f808245018082, /* 2135 */
128'h00d5043300d584b3003796934781e426, /* 2136 */
128'h80826105450164a2644260e200c79863, /* 2137 */
128'h35176090600c02e80363609800043803, /* 2138 */
128'h351785a286269fcfd0ef26a505130000, /* 2139 */
128'hbf5d0785a0019ecfd0ef282505130000, /* 2140 */
128'he0a2282505130000351784aafc26715d, /* 2141 */
128'h892ee45ee486e85aec56f052f44ef84a, /* 2142 */
128'h3a9727298993000039979c0fd0ef4401, /* 2143 */
128'h4a41282b0b1300003b1727aa8a930000, /* 2144 */
128'hd0ef855685de00040b9b9a0fd0ef854e, /* 2145 */
128'h986fd0ef854e03271863470187a6994f, /* 2146 */
128'h03259963458187a697efd0ef855a85de, /* 2147 */
128'hd0ef2aa5051300003517fd4417e30405, /* 2148 */
128'hc299863e8a85008706b3a0a94501964f, /* 2149 */
128'h8733bf6d07a107056394e390fff7c613, /* 2150 */
128'h0b63fff7c693c31986be8b0563900085, /* 2151 */
128'h926fd0ef2145051300003517058e02d6, /* 2152 */
128'h60a6557d91afd0ef2405051300003517, /* 2153 */
128'h6ba26b426ae27a0279a2794274e26406, /* 2154 */
128'hfc56e0d27159b75107a1058580826161, /* 2155 */
128'hf45ef85ae4ceeca6020005138aaa6a05, /* 2156 */
128'h8b2ee46ee86aec66e8caf0a2f486f062, /* 2157 */
128'h3c179c4a0a134981b53ff0ef44818bb2, /* 2158 */
128'h0cb300fa8db30034979351ac0c130000, /* 2159 */
128'hd0ef212505130000351703749b6300fb, /* 2160 */
128'h7c027ba26a0669a6694670a674068a4f, /* 2161 */
128'h85567b4264e685da86266da26d426ce2, /* 2162 */
128'he0ef842abe7fe0efe47ff06f61657ae2, /* 2163 */
128'hf7b3bd5fe0ef892abdbfe0ef8d2abe1f, /* 2164 */
128'h643300a96533010d1d1b0105151b0344, /* 2165 */
128'hb02300acb0238d4191011402150201a4, /* 2166 */
128'h0039f7930985ac1ff0ef4521ef8100ad, /* 2167 */
128'h7139b7ad0485ab1ff0ef0007c50397e2, /* 2168 */
128'h89aaec4ef04af426f822fc06e032e42e, /* 2169 */
128'hb73fe0ef892ab79fe0ef842ab7ffe0ef, /* 2170 */
128'h8d450109179b0105151bb6dfe0ef84aa, /* 2171 */
128'h47818d5d9101178265a2660215028fc1, /* 2172 */
128'h744200c79c63974e00e5883300379713, /* 2173 */
128'hf06f6121863e69e2854e790274a270e2, /* 2174 */
128'h8f2900083703e3148ea907856314d8df, /* 2175 */
128'hf822fc06e032e42e7139b7f100e83023, /* 2176 */
128'he0ef842ab07fe0ef89aaec4ef04af426, /* 2177 */
128'h151baf5fe0ef84aaafbfe0ef892ab01f, /* 2178 */
128'h65a2660215028fc18d450109179b0105, /* 2179 */
128'h00e588330037971347818d5d91011782, /* 2180 */
128'h854e790274a270e2744200c79c63974e, /* 2181 */
128'h8e8907856314d15ff06f6121863e69e2, /* 2182 */
128'h7139b7f100e830238f0900083703e314, /* 2183 */
128'h89aaec4ef04af426f822fc06e032e42e, /* 2184 */
128'ha83fe0ef892aa89fe0ef842aa8ffe0ef, /* 2185 */
128'h8d450109179b0105151ba7dfe0ef84aa, /* 2186 */
128'h47818d5d9101178265a2660215028fc1, /* 2187 */
128'h744200c79c63974e00e5883300379713, /* 2188 */
128'hf06f6121863e69e2854e790274a270e2, /* 2189 */
128'h00083703e31402a686b307856314c9df, /* 2190 */
128'he032e42e7139b7e100e8302302a70733, /* 2191 */
128'ha13fe0ef89aaec4ef04af426f822fc06, /* 2192 */
128'he0ef84aaa07fe0ef892aa0dfe0ef842a, /* 2193 */
128'h15028fc18d450109179b0105151ba01f, /* 2194 */
128'h0037971347818d5d9101178265a26602, /* 2195 */
128'h74a270e2744200c79c63974e00e58833, /* 2196 */
128'he111c21ff06f6121863e69e2854e7902, /* 2197 */
128'h00083703e31402a6d6b3078563144505, /* 2198 */
128'he032e42e7139b7d100e8302302a75733, /* 2199 */
128'h993fe0ef89aaec4ef04af426f822fc06, /* 2200 */
128'he0ef84aa987fe0ef892a98dfe0ef842a, /* 2201 */
128'h15028fc18d450109179b0105151b981f, /* 2202 */
128'h0037971347818d5d9101178265a26602, /* 2203 */
128'h74a270e2744200c79c63974e00e58833, /* 2204 */
128'h6314ba1ff06f6121863e69e2854e7902, /* 2205 */
128'h00e830238f4900083703e3148ec90785, /* 2206 */
128'hf04af426f822fc06e032e42e7139b7f1, /* 2207 */
128'h892a915fe0ef842a91bfe0ef89aaec4e, /* 2208 */
128'h179b0105151b909fe0ef84aa90ffe0ef, /* 2209 */
128'h9101178265a2660215028fc18d450109, /* 2210 */
128'h9c63974e00e588330037971347818d5d, /* 2211 */
128'h863e69e2854e790274a270e2744200c7, /* 2212 */
128'h3703e3148ee907856314b29ff06f6121, /* 2213 */
128'he032e42e7139b7f100e830238f690008, /* 2214 */
128'h8a3fe0ef89aaec4ef04af426f822fc06, /* 2215 */
128'he0ef84aa897fe0ef892a89dfe0ef842a, /* 2216 */
128'h14828fc18cc90109179b0105151b891f, /* 2217 */
128'h0037169347018fc59081178265a26602, /* 2218 */
128'h74a270e2744200c71c6396ae00d98833, /* 2219 */
128'h0533ab1ff06f6121863a69e2854e7902, /* 2220 */
128'he8ca7159bfc9070500a83023e28800f7, /* 2221 */
128'he0d2e4cef0a2d765051300003517892a, /* 2222 */
128'h89aeec66eca6f486f062f45ef85afc56, /* 2223 */
128'hd60a0a1300003a17caffc0ef44018b32, /* 2224 */
128'hd70c0c1300003c17d68b8b9300003b97, /* 2225 */
128'h85a2fff44493c8dfc0ef855204000a93, /* 2226 */
128'h14fd460140900cb3c7ffc0ef8885855e, /* 2227 */
128'h85520566186397ce00f905b300361793, /* 2228 */
128'h6622c59fc0ef856285a2c61fc0efe432, /* 2229 */
128'h1be32405e12984aaa17ff0ef854a85ce, /* 2230 */
128'h70a6c39fc0efd7e5051300003517fb54, /* 2231 */
128'h7b427ae26a0669a664e6694685267406, /* 2232 */
128'h876600167693808261656ce27c027ba2, /* 2233 */
128'hbfc154fdbf590605e198e3988726c291, /* 2234 */
128'hf0a2ca2505130000351784aaeca67159, /* 2235 */
128'hec66f062f45ef85afc56e0d2e4cee8ca, /* 2236 */
128'h3997bd9fc0ef44018ab2892ee86af486, /* 2237 */
128'h3b97f8ab0b1300003b17c8a989930000, /* 2238 */
128'h3c97c82c0c1300003c17f8ab8b930000, /* 2239 */
128'hba7fc0ef854e04000a13c8ac8c930000, /* 2240 */
128'hc0ef856285a2000bbd03cba500147793, /* 2241 */
128'h00f485b300361793fffd45134601b95f, /* 2242 */
128'h85a2b79fc0efe432854e05561c6397ca, /* 2243 */
128'h92fff0ef852685ca6622b71fc0ef8566, /* 2244 */
128'h051300003517fb441ae32405e5298d2a, /* 2245 */
128'h694664e6856a740670a6b51fc0efc965, /* 2246 */
128'h6d426ce27c027ba27b427ae26a0669a6, /* 2247 */
128'h876a00167693bf49000b3d0380826165, /* 2248 */
128'hb7e15d7db7790605e198e398872ac291, /* 2249 */
128'he4a6bb25051300003517842ae8a2711d, /* 2250 */
128'hfc4eec86e862ec5ef05af456f852e0ca, /* 2251 */
128'h091300003917aedfc0ef4c018ab284ae, /* 2252 */
128'h8b9300003b97ba6b0b1300003b17b9e9, /* 2253 */
128'h000c099bacbfc0ef854a10000a13baeb, /* 2254 */
128'h008c1793010c1713abffc0ef855a85ce, /* 2255 */
128'h020c17138fd9018c17130187e7b38fd9, /* 2256 */
128'h17138fd9030c17138fd9028c17138fd9, /* 2257 */
128'h972600e406b30036171346018fd9038c, /* 2258 */
128'h855e85cea7bfc0efe432854a05561763, /* 2259 */
128'h89aa831ff0ef852285a66622a73fc0ef, /* 2260 */
128'hb985051300003517f94c19e30c05e91d, /* 2261 */
128'h79e2690664a6854e644660e6a53fc0ef, /* 2262 */
128'he31c808261256c426be27b027aa27a42, /* 2263 */
128'h84aaf4a67119bff159fdb74d0605e29c, /* 2264 */
128'he8d2eccef0caf8a2ac85051300003517, /* 2265 */
128'hec6efc86f06af466f862fc5ee0dae4d6, /* 2266 */
128'h0a1300003a179fdfc0ef44018b32892e, /* 2267 */
128'h498507f00b93ab6c8c9300003c97aaea, /* 2268 */
128'h08000a93ab4d0d1300003d1703f00c13, /* 2269 */
128'h873b9c9fc0ef856685a29d1fc0ef8552, /* 2270 */
128'h003617934601008995b300e99733408b, /* 2271 */
128'hc0efe432855205661a6397ca00f486b3, /* 2272 */
128'h852685ca662299dfc0ef856a85a29a5f, /* 2273 */
128'h3517fb541be32405e1398daaf5aff0ef, /* 2274 */
128'h856e744670e697dfc0efac2505130000, /* 2275 */
128'h7c427be26b066aa66a4669e6790674a6, /* 2276 */
128'he38c008c6663808261096de27d027ca2, /* 2277 */
128'hb7f15dfdbfe5e298e398bf610605e28c, /* 2278 */
128'hf8a29e2505130000351784aaf4a67119, /* 2279 */
128'hf466f862fc5ee0dae4d6e8d2eccef0ca, /* 2280 */
128'h917fc0ef44018b32892eec6efc86f06a, /* 2281 */
128'h9d0c8c9300003c979c8a0a1300003a17, /* 2282 */
128'h0d1300003d1703f00c13498507f00b93, /* 2283 */
128'h856685a28ebfc0ef855208000a939ced, /* 2284 */
128'h008996b300f997b3408b87bb8e3fc0ef, /* 2285 */
128'h85b3003617134601fff6c693fff7c793, /* 2286 */
128'h8b7fc0efe432855205661a63974a00e4, /* 2287 */
128'hf0ef852685ca66228affc0ef856a85a2, /* 2288 */
128'h00003517fb5417e32405e1398daae6cf, /* 2289 */
128'h74a6856e744670e688ffc0ef9d450513, /* 2290 */
128'h7ca27c427be26b066aa66a4669e67906, /* 2291 */
128'he194e314008c6663808261096de27d02, /* 2292 */
128'h7119b7f15dfdbfe5e19ce31cbf610605, /* 2293 */
128'hf0caf8a28f4505130000351784aaf4a6, /* 2294 */
128'hf06af466f862fc5ee0dae4d6e8d2ecce, /* 2295 */
128'h3997829fc0ef44018a32892eec6efc86, /* 2296 */
128'h0a938e2c0c1300003c178da989930000, /* 2297 */
128'h00003c9703f00b9308100b134d0507f0, /* 2298 */
128'hc0ef856285a2ffcfc0ef854e8dcc8c93, /* 2299 */
128'h173300fd17b3408b07bb408a873bff4f, /* 2300 */
128'h008d16b300fd17b30024079b8f5d00ed, /* 2301 */
128'h003616934601fff7c893fff743138fd5, /* 2302 */
128'hc0efe432854e05461c6396ca00d48533, /* 2303 */
128'h852685ca6622facfc0ef856685a2fb4f, /* 2304 */
128'h1be3080007932405ed298daad6aff0ef, /* 2305 */
128'h70e6f88fc0ef8ce5051300003517f8f4, /* 2306 */
128'h6b066aa66a4669e6790674a6856e7446, /* 2307 */
128'h7813808261096de27d027ca27c427be2, /* 2308 */
128'he28c85c60008036385be008bea630016, /* 2309 */
128'hbfc5859afe080be385bab7610605e10c, /* 2310 */
128'h051300002517892af0ca7119bf755dfd, /* 2311 */
128'hfc86ec6ef06af466fc5ee8d2ecce7de5, /* 2312 */
128'h4b81e03289aef862e0dae4d6f4a6f8a2, /* 2313 */
128'h00002c977c4a0a1300002a17f12fc0ef, /* 2314 */
128'h47854da17d4d0d1300002d177ccc8c93, /* 2315 */
128'hee6fc0ef85524401003b949b01779c33, /* 2316 */
128'hfffc4a93edafc0ef856685da00848b3b, /* 2317 */
128'h1063974e00e908330036171367824601, /* 2318 */
128'hc0ef856a85daebcfc0efe432855206f6, /* 2319 */
128'he9318b2ac72ff0ef854a85ce6622eb4f, /* 2320 */
128'h90e3040007932b85fbb41be38c562405, /* 2321 */
128'h70e6e88fc0ef7ce5051300002517fafb, /* 2322 */
128'h6b066aa66a4669e6790674a6855a7446, /* 2323 */
128'h7513808261096de27d027ca27c427be2, /* 2324 */
128'h060500b83023e30c85d6e11185e20016, /* 2325 */
128'h892af4cef8cafca67175b7e95b7db749, /* 2326 */
128'he4dee8daecd6f0d269850200051384ae, /* 2327 */
128'h8acae032f46ee122e506f86afc66e0e2, /* 2328 */
128'h0c1300003c174b014a098ba68a6ff0ef, /* 2329 */
128'ha60d0d1300003d179c4989934ca12f6c, /* 2330 */
128'h866e04fd966396d6003d969367824d81, /* 2331 */
128'h8bca4785ed4d842abb6ff0ef854a85a6, /* 2332 */
128'hc0ef742505130000251702fa18638aa6, /* 2333 */
128'h7a0679a6794674e6640a60aa8522dd4f, /* 2334 */
128'h61497da27d427ce26c066ba66b466ae6, /* 2335 */
128'he0ef842a916fe0efec36b7754a058082, /* 2336 */
128'h67a2904fe0efe42a90afe0efe82a910f, /* 2337 */
128'h15028c510106161b8d5d0105151b6642, /* 2338 */
128'h24a7bc23000037978d4166e291011402, /* 2339 */
128'h00fb86330006c683018786b34781e288, /* 2340 */
128'hf7b3ff9795e300d600230ff6f6930785, /* 2341 */
128'h001b079bfcffe0ef4521ef910ba1033d, /* 2342 */
128'hfbbfe0ef0007c50397ea8b8d00078b1b, /* 2343 */
128'hf4cef8cafca67175bfb1547dbf050d85, /* 2344 */
128'he8daecd6f0d269850200051384ae892a, /* 2345 */
128'he032f46ee122e506f86afc66e0e2e4de, /* 2346 */
128'h00003c174b014a098ba6f85fe0ef8aca, /* 2347 */
128'h0d1300003d179c4989934ca11dcc0c13, /* 2348 */
128'h04fd966396d6003d969367824d8193ed, /* 2349 */
128'h4785ed4d842aa94ff0ef854a85a6866e, /* 2350 */
128'h620505130000251702fa18638aa68bca, /* 2351 */
128'h79a6794674e6640a60aa8522cb2fc0ef, /* 2352 */
128'h7da27d427ce26c066ba66b466ae67a06, /* 2353 */
128'h842aff5fd0efec36b7754a0580826149, /* 2354 */
128'hfe3fd0efe42afe9fd0efe82afeffd0ef, /* 2355 */
128'h8c510106161b8d5d0105151b664267a2, /* 2356 */
128'hbf23000037978d4166e2910114021502, /* 2357 */
128'h86330006d683018786b34781e28812a7, /* 2358 */
128'hff9795e300d6102392c116c2078900fb, /* 2359 */
128'h079beadfe0ef4521ef910ba1033df7b3, /* 2360 */
128'he0ef0007c50397ea8b8d00078b1b001b, /* 2361 */
128'h711980826505bfb1547dbf050d85e99f, /* 2362 */
128'h892e962af0caf8a2fff5861389b2ecce, /* 2363 */
128'he8d2f4a655c505130000251785aa842a, /* 2364 */
128'hfc86ec6ef06af466f862fc5ee0dae4d6, /* 2365 */
128'h44854a81e03e00395793bd0fc0efe436, /* 2366 */
128'h550b8b9300002b97550b0b1300002b17, /* 2367 */
128'h550c8c9300002c97550c0c1300002c17, /* 2368 */
128'h558d8d9300002d97558d0d1300002d17, /* 2369 */
128'h000025170299f863058a0a1300003a17, /* 2370 */
128'h74a68556744670e6b7efc0ef54c50513, /* 2371 */
128'h7ca27c427be26b066aa66a4669e67906, /* 2372 */
128'hb56fc0ef855a85a6808261096de27d02, /* 2373 */
128'hc0ef8562b4afc0ef855e85ce00098663, /* 2374 */
128'hf0ef85226582b3cfc0ef856a85e6b44f, /* 2375 */
128'h6722010a2783b2cfc0ef856ee129952f, /* 2376 */
128'h051300002517c985000a358302f74c63, /* 2377 */
128'h561300195593008a3783b10fc0ef4ce5, /* 2378 */
128'h4b850513000025179782852295a20049, /* 2379 */
128'h2705051300002517b7d14a89af2fc0ef, /* 2380 */
128'h0513000025177179bf890485ae2fc0ef, /* 2381 */
128'hc45fe0efe44ee84aec26f022f4064a65, /* 2382 */
128'hab6fc0ef4a4505130000251704000593, /* 2383 */
128'h00002517aaafc0ef4c05051300002517, /* 2384 */
128'h2205051300002517a9efc0ef4e450513, /* 2385 */
128'h95b3497901f499934441a90fc0ef4485, /* 2386 */
128'he73ff0ef240501358533460546850084, /* 2387 */
128'h614569a2694264e2740270a2ff2417e3, /* 2388 */
128'h46814881470100c5131b460580828082, /* 2389 */
128'h000780234000081387f245a901f61e13, /* 2390 */
128'h802397aa0007802397aa0007802397aa, /* 2391 */
128'h02b71d632705fe0813e397aa387d0007, /* 2392 */
128'h86b33e800513c00026f38e15c0202673, /* 2393 */
128'h45bb02c747334000059302a687334116, /* 2394 */
128'h05130000251702a7473302a767b302b3, /* 2395 */
128'h28f3c02026f3fac710e39f0fc06f47e5, /* 2396 */
128'h4505f7bff0ef4501e4061141bf51c000, /* 2397 */
128'hf69ff0ef4511f6fff0ef4509f75ff0ef, /* 2398 */
128'h1502bff1f5dff0ef4541f63ff0ef4521, /* 2399 */
128'h6388440007b78082e388440007b79101, /* 2400 */
128'h25016b880007b823440007b780822501, /* 2401 */
128'h0085979b808225017b88440007b78082, /* 2402 */
128'h2581f788440007b78d510106161b8d5d, /* 2403 */
128'h079300b76f630007871b440006374781, /* 2404 */
128'hffe537fdc3198b097a98440006b73e80, /* 2405 */
128'h670397360027971380827388440007b7, /* 2406 */
128'h4785e406e0221141bfc1f61807850007, /* 2407 */
128'hfedff0ef0045551b35fd00b7d763842a, /* 2408 */
128'h00044503943e3ee7879300002797883d, /* 2409 */
128'h004007b7711da45fe06f014160a26402, /* 2410 */
128'h0189571b3006869300a7893b6685e0ca, /* 2411 */
128'h0034e4a6e8a20587e7938f550089179b, /* 2412 */
128'hc43aec86c63e4589454d84ae842a4601, /* 2413 */
128'h458946010034f47ff0eff456f852fc4e, /* 2414 */
128'h4589460189aa0034f39ff0ef454d8a2a, /* 2415 */
128'h02f8073b46a158614781f2bff0ef454d, /* 2416 */
128'h00b6002300ea55b30387071b963e0810, /* 2417 */
128'h963e083000b6002300e9d5b300f48633, /* 2418 */
128'h45a1fcd799e3078500e6002300e55733, /* 2419 */
128'hc0ef45a5051300001517f37ff0ef854a, /* 2420 */
128'h07bb4a2144ca8a9300001a974981864f, /* 2421 */
128'h4589ff07c50397ba9381101817820134, /* 2422 */
128'hff4991e383afc0ef8556f07ff0ef2985, /* 2423 */
128'h854a45a182afc0effb85051300002517, /* 2424 */
128'h816fc0ef40c5051300001517ee9ff0ef, /* 2425 */
128'h013407bb4a213fea8a9300001a974981, /* 2426 */
128'hf0ef298545890007c50397a693811782, /* 2427 */
128'h00002517ff4992e3feffb0ef8556ebbf, /* 2428 */
128'he9dff0ef45a1854afdffb0eff6c50513, /* 2429 */
128'h19974481fcbfb0ef3c05051300001517, /* 2430 */
128'h10181782009407bb49213b2989930000, /* 2431 */
128'he6dff0ef24854589ff87c50397ba9381, /* 2432 */
128'h051300002517ff2491e3fa1fb0ef854e, /* 2433 */
128'h79e2690664a6644660e6f91fb0eff1e5, /* 2434 */
128'hfc4ee0cae4a6711d808261257aa27a42, /* 2435 */
128'h8b2e89aaf852e8a2ec86ec5ef05af456, /* 2436 */
128'h0004841b44000bb7ff860a9b44818932, /* 2437 */
128'hf0ef002c055464630164053b00998a33, /* 2438 */
128'hd0ef002c9201855216024089063be3df, /* 2439 */
128'h2b174ac131ca0a1300001a174401da3f, /* 2440 */
128'h64a6644660e603246763eaab0b130000, /* 2441 */
128'h808261256be27b027aa27a4279e26906, /* 2442 */
128'hb02304a1df3ff0ef00c4541b85d22421, /* 2443 */
128'hb0ef8552db1ff0ef852245a1bf69008b, /* 2444 */
128'hc50397ce93811782009407bb4481ee5f, /* 2445 */
128'hec7fb0ef8552d93ff0ef248545890007, /* 2446 */
128'h1141bf692441ebdfb0ef855aff5492e3, /* 2447 */
128'h0517ea9fb0efe406cf85051300002517, /* 2448 */
128'h60a200055c63b7df70eff2a505130000, /* 2449 */
128'hb06f0141cec505130000251740a005b3, /* 2450 */
128'h0513000025179e7fe06f014160a2e85f, /* 2451 */
128'hf04af426f822fc067139feefe06f1fe5, /* 2452 */
128'h00002517fa6fe0efe05ae456e852ec4e, /* 2453 */
128'h2917440009b74401fccfe0ef13c50513, /* 2454 */
128'h639097ce00341793449513a909130000, /* 2455 */
128'hfe9416e3e2bfb0ef0405854a0004059b, /* 2456 */
128'h04b723ab0b1300002b174901be0f80ef, /* 2457 */
128'h0a1300002a17116a8a9300002a974400, /* 2458 */
128'h090585560007c783016907b34991126a, /* 2459 */
128'hde7fb0ef8622240125816080608ce09c, /* 2460 */
128'h1be3dd9fb0ef25818552688c0004b823, /* 2461 */
128'h02f7646347190054579b0ff47413fd39, /* 2462 */
128'h97ba439c97ba078a6b07071300000717, /* 2463 */
128'h8522da9fb0ef0e650513000025178782, /* 2464 */
128'hb0ef0e25051300002517a001941fe0ef, /* 2465 */
128'h051300002517b7f5edbff0ef8522d95f, /* 2466 */
128'h00002517bfe9aa3ff0efd81fb0ef0de5, /* 2467 */
128'h2517b7e1c60f80efd6ffb0ef0dc50513, /* 2468 */
128'hbf5db7bff0efd5dfb0ef0da505130000, /* 2469 */
128'h00000000000000000000000000000000, /* 2470 */
128'h00000000000000000000000000000000, /* 2471 */
128'h00000000000000000000000000000000, /* 2472 */
128'h00000000000000000000000000000000, /* 2473 */
128'h00000000000000000000000000000000, /* 2474 */
128'h00000000000000000000000000000000, /* 2475 */
128'h00000000000000000000000000000000, /* 2476 */
128'h00000000000000000000000000000000, /* 2477 */
128'h00000000000000000000000000000000, /* 2478 */
128'h00000000000000000000000000000000, /* 2479 */
128'h08082828282828080808080808080808, /* 2480 */
128'h08080808080808080808080808080808, /* 2481 */
128'h101010101010101010101010101010a0, /* 2482 */
128'h10101010101004040404040404040404, /* 2483 */
128'h01010101010101010141414141414110, /* 2484 */
128'h10101010100101010101010101010101, /* 2485 */
128'h02020202020202020242424242424210, /* 2486 */
128'h08101010100202020202020202020202, /* 2487 */
128'h00000000000000000000000000000000, /* 2488 */
128'h00000000000000000000000000000000, /* 2489 */
128'h101010101010101010101010101010a0, /* 2490 */
128'h10101010101010101010101010101010, /* 2491 */
128'h01010101010101010101010101010101, /* 2492 */
128'h02010101010101011001010101010101, /* 2493 */
128'h02020202020202020202020202020202, /* 2494 */
128'h02020202020202021002020202020202, /* 2495 */
128'hc1bdceee242070dbe8c7b756d76aa478, /* 2496 */
128'hfd469501a83046134787c62af57c0faf, /* 2497 */
128'h895cd7beffff5bb18b44f7af698098d8, /* 2498 */
128'h49b40821a679438efd9871936b901122, /* 2499 */
128'he9b6c7aa265e5a51c040b340f61e2562, /* 2500 */
128'he7d3fbc8d8a1e68102441453d62f105d, /* 2501 */
128'h455a14edf4d50d87c33707d621e1cde6, /* 2502 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /* 2503 */
128'hfde5380c6d9d61228771f681fffa3942, /* 2504 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /* 2505 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /* 2506 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /* 2507 */
128'hfc93a039ab9423a7432aff97f4292244, /* 2508 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /* 2509 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /* 2510 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /* 2511 */
128'h0c07020d08030e09040f0a05000b0601, /* 2512 */
128'h020f0c090603000d0a0704010e0b0805, /* 2513 */
128'h09020b040d060f08010a030c050e0700, /* 2514 */
128'h6c5f7465735f64735f63736972776f6c, /* 2515 */
128'h6e67696c615f64730000000000006465, /* 2516 */
128'h645f6b6c635f64730000000000000000, /* 2517 */
128'h69747465735f64730000000000007669, /* 2518 */
128'h735f646d635f6473000000000000676e, /* 2519 */
128'h74657365725f64730000000074726174, /* 2520 */
128'h6e636b6c625f64730000000000000000, /* 2521 */
128'h69736b6c625f64730000000000000074, /* 2522 */
128'h6f656d69745f6473000000000000657a, /* 2523 */
128'h655f7172695f64730000000000007475, /* 2524 */
128'h5f63736972776f6c000000000000006e, /* 2525 */
128'h00000000646d635f74726174735f6473, /* 2526 */
128'h746e695f746961775f63736972776f6c, /* 2527 */
128'h000000000067616c665f747075727265, /* 2528 */
128'h00007172695f64735f63736972776f6c, /* 2529 */
128'h695f646d635f64735f63736972776f6c, /* 2530 */
128'h5f63736972776f6c0000000000007172, /* 2531 */
128'h007172695f646e655f617461645f6473, /* 2532 */
128'h0000000087fe9e880000000087feb160, /* 2533 */
128'h004c4b40004c4b400030000020000000, /* 2534 */
128'h6d6d5f6472616f62000000020000ffff, /* 2535 */
128'h0000000087fe4eaa0064637465675f63, /* 2536 */
128'h0000000087fe4d180000000087fe4aba, /* 2537 */
128'h00000000000000000000000000000000, /* 2538 */
128'hffffb994ffffb990ffffb990ffffb96c, /* 2539 */
128'hffffb998ffffb998ffffb998ffffb998, /* 2540 */
128'hffffc9baffffc9b4ffffc9aeffffc80a, /* 2541 */
128'h0000000087feb4880000000087feb478, /* 2542 */
128'h0000000087feb4b00000000087feb498, /* 2543 */
128'h0000000087feb4e00000000087feb4c8, /* 2544 */
128'h0000000087feb5100000000087feb4f8, /* 2545 */
128'h0000000087feb5400000000087feb528, /* 2546 */
128'h0000000087feb5700000000087feb558, /* 2547 */
128'h40040300400402004004010040040000, /* 2548 */
128'h40050000400405004004040140040400, /* 2549 */
128'h30000000000000030000000040050100, /* 2550 */
128'h60000000000000053000000000000001, /* 2551 */
128'h70000000000000027000000000000004, /* 2552 */
128'h00000001400000007000000000000000, /* 2553 */
128'h00000005000000012000000000000006, /* 2554 */
128'h20000000000000020000000040000000, /* 2555 */
128'h00000000100000000000000100000000, /* 2556 */
128'h1e19140f0d0c0a000000000000000000, /* 2557 */
128'h000186a00000271050463c37322d2823, /* 2558 */
128'h017d7840017d784000989680000f4240, /* 2559 */
128'h031975000319750002faf080018cba80, /* 2560 */
128'h02faf08005f5e10002faf080017d7840, /* 2561 */
128'h00000020000000000bebc2000c65d400, /* 2562 */
128'h00000200000001000000008000000040, /* 2563 */
128'h00002000000010000000080000000400, /* 2564 */
128'h0000c000000080000000600000004000, /* 2565 */
128'h37363534333231300002000000010000, /* 2566 */
128'h2043534952776f4c4645444342413938, /* 2567 */
128'h746f6f622d7520646573696d696e696d, /* 2568 */
128'h00000000647261432d445320726f6620, /* 2569 */
128'hfffff974fffff98afffff976fffff962, /* 2570 */
128'h00000000fffff9aefffff974fffff99c, /* 2571 */
128'he00600003800000039080000edfe0dd0, /* 2572 */
128'h00000000100000001100000028000000, /* 2573 */
128'h0000000000000000a806000059010000, /* 2574 */
128'h00000000010000000000000000000000, /* 2575 */
128'h02000000000000000400000003000000, /* 2576 */
128'h020000000f0000000400000003000000, /* 2577 */
128'h2c6874651b0000001400000003000000, /* 2578 */
128'h007665642d657261622d656e61697261, /* 2579 */
128'h2c687465260000001000000003000000, /* 2580 */
128'h0100000000657261622d656e61697261, /* 2581 */
128'h1a0000000300000000006e65736f6863, /* 2582 */
128'h303140747261752f636f732f2c000000, /* 2583 */
128'h0000003030323531313a303030303030, /* 2584 */
128'h00000000737570630100000002000000, /* 2585 */
128'h01000000000000000400000003000000, /* 2586 */
128'h000000000f0000000400000003000000, /* 2587 */
128'h40787d01380000000400000003000000, /* 2588 */
128'h03000000000000304075706301000000, /* 2589 */
128'h0300000080f0fa024b00000004000000, /* 2590 */
128'h03000000007570635b00000004000000, /* 2591 */
128'h03000000000000006700000004000000, /* 2592 */
128'h0000000079616b6f6b00000005000000, /* 2593 */
128'h7a6874651b0000001300000003000000, /* 2594 */
128'h0000766373697200656e61697261202c, /* 2595 */
128'h34367672720000000b00000003000000, /* 2596 */
128'h0b000000030000000000636466616d69, /* 2597 */
128'h0000393376732c76637369727c000000, /* 2598 */
128'h01000000850000000000000003000000, /* 2599 */
128'h6f72746e6f632d747075727265746e69, /* 2600 */
128'h04000000030000000000000072656c6c, /* 2601 */
128'h0000000003000000010000008f000000, /* 2602 */
128'h1b0000000f00000003000000a0000000, /* 2603 */
128'h000063746e692d7570632c7663736972, /* 2604 */
128'h01000000b50000000400000003000000, /* 2605 */
128'h01000000bb0000000400000003000000, /* 2606 */
128'h01000000020000000200000002000000, /* 2607 */
128'h0030303030303030384079726f6d656d, /* 2608 */
128'h6f6d656d5b0000000700000003000000, /* 2609 */
128'h67000000100000000300000000007972, /* 2610 */
128'h00000008000000000000008000000000, /* 2611 */
128'h0300000000636f730100000002000000, /* 2612 */
128'h03000000020000000000000004000000, /* 2613 */
128'h03000000020000000f00000004000000, /* 2614 */
128'h616972612c6874651b0000001f000000, /* 2615 */
128'h706d697300636f732d657261622d656e, /* 2616 */
128'h000000000300000000007375622d656c, /* 2617 */
128'h303240746e696c6301000000c3000000, /* 2618 */
128'h0d000000030000000000003030303030, /* 2619 */
128'h30746e696c632c76637369721b000000, /* 2620 */
128'hca000000100000000300000000000000, /* 2621 */
128'h07000000010000000300000001000000, /* 2622 */
128'h00000000670000001000000003000000, /* 2623 */
128'h0300000000000c000000000000000002, /* 2624 */
128'h006c6f72746e6f63de00000008000000, /* 2625 */
128'h7075727265746e690100000002000000, /* 2626 */
128'h3030634072656c6c6f72746e6f632d74, /* 2627 */
128'h04000000030000000000000030303030, /* 2628 */
128'h04000000030000000000000000000000, /* 2629 */
128'h0c00000003000000010000008f000000, /* 2630 */
128'h003063696c702c76637369721b000000, /* 2631 */
128'h03000000a00000000000000003000000, /* 2632 */
128'h0b00000001000000ca00000010000000, /* 2633 */
128'h10000000030000000900000001000000, /* 2634 */
128'h000000000000000c0000000067000000, /* 2635 */
128'he8000000040000000300000000000004, /* 2636 */
128'hfb000000040000000300000007000000, /* 2637 */
128'hb5000000040000000300000003000000, /* 2638 */
128'hbb000000040000000300000002000000, /* 2639 */
128'h75626564010000000200000002000000, /* 2640 */
128'h0000304072656c6c6f72746e6f632d67, /* 2641 */
128'h637369721b0000001000000003000000, /* 2642 */
128'h03000000003331302d67756265642c76, /* 2643 */
128'hffff000001000000ca00000008000000, /* 2644 */
128'h00000000670000001000000003000000, /* 2645 */
128'h03000000001000000000000000000000, /* 2646 */
128'h006c6f72746e6f63de00000008000000, /* 2647 */
128'h30303140747261750100000002000000, /* 2648 */
128'h08000000030000000000003030303030, /* 2649 */
128'h03000000003035373631736e1b000000, /* 2650 */
128'h00000010000000006700000010000000, /* 2651 */
128'h04000000030000000010000000000000, /* 2652 */
128'h040000000300000080f0fa024b000000, /* 2653 */
128'h040000000300000000c2010006010000, /* 2654 */
128'h04000000030000000200000014010000, /* 2655 */
128'h04000000030000000100000025010000, /* 2656 */
128'h04000000030000000200000030010000, /* 2657 */
128'h0100000002000000040000003a010000, /* 2658 */
128'h3030303240636d6d2d63736972776f6c, /* 2659 */
128'h10000000030000000000000030303030, /* 2660 */
128'h00000000000000200000000067000000, /* 2661 */
128'h14010000040000000300000000000100, /* 2662 */
128'h25010000040000000300000002000000, /* 2663 */
128'h1b0000000c0000000300000002000000, /* 2664 */
128'h0200000000636d6d2d63736972776f6c, /* 2665 */
128'h406874652d63736972776f6c01000000, /* 2666 */
128'h03000000000000003030303030303033, /* 2667 */
128'h2d63736972776f6c1b0000000c000000, /* 2668 */
128'h5b000000080000000300000000687465, /* 2669 */
128'h0400000003000000006b726f7774656e, /* 2670 */
128'h04000000030000000200000014010000, /* 2671 */
128'h06000000030000000300000025010000, /* 2672 */
128'h0300000000007fe3023e180047010000, /* 2673 */
128'h00000030000000006700000010000000, /* 2674 */
128'h01000000020000000080000000000000, /* 2675 */
128'h303440646e7277682d63736972776f6c, /* 2676 */
128'h0e000000030000000000303030303030, /* 2677 */
128'h6e7277682d63736972776f6c1b000000, /* 2678 */
128'h67000000100000000300000000000064, /* 2679 */
128'h00100000000000000000004000000000, /* 2680 */
128'h09000000020000000200000002000000, /* 2681 */
128'h2300736c6c65632d7373657264646123, /* 2682 */
128'h61706d6f6300736c6c65632d657a6973, /* 2683 */
128'h6f647473006c65646f6d00656c626974, /* 2684 */
128'h65736162656d697400687461702d7475, /* 2685 */
128'h6b636f6c630079636e6575716572662d, /* 2686 */
128'h63697665640079636e6575716572662d, /* 2687 */
128'h75746174730067657200657079745f65, /* 2688 */
128'h2d756d6d006173692c76637369720073, /* 2689 */
128'h230074696c70732d626c740065707974, /* 2690 */
128'h00736c6c65632d747075727265746e69, /* 2691 */
128'h6f72746e6f632d747075727265746e69, /* 2692 */
128'h646e6168702c78756e696c0072656c6c, /* 2693 */
128'h727265746e69007365676e617200656c, /* 2694 */
128'h6572006465646e657478652d73747075, /* 2695 */
128'h616d2c76637369720073656d616e2d67, /* 2696 */
128'h766373697200797469726f6972702d78, /* 2697 */
128'h70732d746e6572727563007665646e2c, /* 2698 */
128'h61702d747075727265746e6900646565, /* 2699 */
128'h0073747075727265746e6900746e6572, /* 2700 */
128'h6f692d6765720074666968732d676572, /* 2701 */
128'h63616d2d6c61636f6c0068746469772d, /* 2702 */
128'h0000000000000000737365726464612d, /* 2703 */
128'h0000000000203a642520656369766544, /* 2704 */
128'h00203a6425206563697665642073250a, /* 2705 */
128'h00000000203a6425206563697665440a, /* 2706 */
128'h000a656369766564206e776f6e6b6e75, /* 2707 */
128'h00000a2973252c73252870756b6f6f6c, /* 2708 */
128'h7265206c616e7265746e692070636864, /* 2709 */
128'h00000000000000000a7025202c726f72, /* 2710 */
128'h5145525f5043484420676e69646e6553, /* 2711 */
128'h4b434120504348440000000a54534555, /* 2712 */
128'h696c432050434844000000000000000a, /* 2713 */
128'h203a7373657264644120504920746e65, /* 2714 */
128'h0000000a64252e64252e64252e642520, /* 2715 */
128'h73657264644120504920726576726553, /* 2716 */
128'h0a64252e64252e64252e642520203a73, /* 2717 */
128'h6120726574756f520000000000000000, /* 2718 */
128'h252e64252e642520203a737365726464, /* 2719 */
128'h6b73616d2074654e0000000a64252e64, /* 2720 */
128'h64252e642520203a7373657264646120, /* 2721 */
128'h697420657361654c000a64252e64252e, /* 2722 */
128'h7364253a6d64253a686425203d20656d, /* 2723 */
128'h3d206e69616d6f44000000000000000a, /* 2724 */
128'h4820746e65696c4300000a2273252220, /* 2725 */
128'h000a22732522203d20656d616e74736f, /* 2726 */
128'h000000000a44455050494b53204b4341, /* 2727 */
128'h000000000000000a4b414e2050434844, /* 2728 */
128'h73657264646120646574736575716552, /* 2729 */
128'h0000000000000a646573756665722073, /* 2730 */
128'h000000000000000a732520726f727245, /* 2731 */
128'h6e6f6974706f2064656c646e61686e75, /* 2732 */
128'h656c646e61686e55000000000a642520, /* 2733 */
128'h64252065646f63706f20504348442064, /* 2734 */
128'h20676e69646e6553000000000000000a, /* 2735 */
128'h000a595245564f435349445f50434844, /* 2736 */
128'h00000000000a29732528726f72726570, /* 2737 */
128'h3a2043414d2073250000000030687465, /* 2738 */
128'h3a583230253a583230253a5832302520, /* 2739 */
128'h000a583230253a583230253a58323025, /* 2740 */
128'h484420646e65732074276e646c756f43, /* 2741 */
128'h206e6f20595245564f43534944205043, /* 2742 */
128'h00000a7325203a732520656369766564, /* 2743 */
128'h5043484420726f6620676e6974696157, /* 2744 */
128'h2020202020202020000a524546464f5f, /* 2745 */
128'h00000000000063250000000000000020, /* 2746 */
128'h0000005832302520000000000000002e, /* 2747 */
128'h00000000732573250000000000000a0a, /* 2748 */
128'h00000000007325203a646c697542202c, /* 2749 */
128'h73257a4820756c250000000000007325, /* 2750 */
128'h0000000000756c250000000000000000, /* 2751 */
128'h0073257a4863252000000000646c252e, /* 2752 */
128'h00000000007325736574794220756c25, /* 2753 */
128'h00003a786c3830250073254269632520, /* 2754 */
128'h000a73252020202000786c6c2a302520, /* 2755 */
128'h000000203a5d64255b6e6f6974636553, /* 2756 */
128'h727265207974696e6173207264646170, /* 2757 */
128'h2c7825286e666c6500000a702520726f, /* 2758 */
128'h000000000a3b29782578302c78257830, /* 2759 */
128'h782578302c302c7825287465736d656d, /* 2760 */
128'h464f5f4f4c43414d00000000000a3b29, /* 2761 */
128'h464f5f494843414d0000000054455346, /* 2762 */
128'h46464f5f524c50540000000054455346, /* 2763 */
128'h46464f5f534346540000000000544553, /* 2764 */
128'h4c5254434f49444d0000000000544553, /* 2765 */
128'h46464f5f534346520054455346464f5f, /* 2766 */
128'h5346464f5f5253520000000000544553, /* 2767 */
128'h46464f5f444142520000000000005445, /* 2768 */
128'h46464f5f524c50520000000000544553, /* 2769 */
128'h000000003f3f3f3f0000000000544553, /* 2770 */
128'h000064252b54455346464f5f524c5052, /* 2771 */
128'h6f746f72502050490000000000000047, /* 2772 */
128'h00000000000000000a50495049203d20, /* 2773 */
128'h6f746f72502050490000000000000054, /* 2774 */
128'h6f746f7250205049000a504745203d20, /* 2775 */
128'h6165682074736574000a505550203d20, /* 2776 */
128'h6e6f6320747365740000000a3a726564, /* 2777 */
128'h6f746f7250205049000a3a73746e6574, /* 2778 */
128'h6f746f7250205049000a504449203d20, /* 2779 */
128'h6f746f725020504900000a5054203d20, /* 2780 */
128'h00000000000000000a50434344203d20, /* 2781 */
128'h6f746f72502050490000000000000036, /* 2782 */
128'h00000000000000000a50565352203d20, /* 2783 */
128'h000a455247203d206f746f7250205049, /* 2784 */
128'h000a505345203d206f746f7250205049, /* 2785 */
128'h00000a4841203d206f746f7250205049, /* 2786 */
128'h000a50544d203d206f746f7250205049, /* 2787 */
128'h5054454542203d206f746f7250205049, /* 2788 */
128'h6f746f72502050490000000000000a48, /* 2789 */
128'h000000000000000a5041434e45203d20, /* 2790 */
128'h6f746f7250205049000000000000004d, /* 2791 */
128'h00000000000000000a504d4f43203d20, /* 2792 */
128'h0a50544353203d206f746f7250205049, /* 2793 */
128'h6f746f72502050490000000000000000, /* 2794 */
128'h00000000000a4554494c504455203d20, /* 2795 */
128'h0a534c504d203d206f746f7250205049, /* 2796 */
128'h6f746f72502050490000000000000000, /* 2797 */
128'h6f746f7270205049000a574152203d20, /* 2798 */
128'h2820646574726f707075736e75203d20, /* 2799 */
128'h79745f6f746f7270000000000a297825, /* 2800 */
128'h0000000000000a78257830203d206570, /* 2801 */
128'h727265746e692064656c646e61686e75, /* 2802 */
128'h414d2070757465530000000a21747075, /* 2803 */
128'h4d454f2049505351000a726464612043, /* 2804 */
128'h0000000000000a7825203d205d64255b, /* 2805 */
128'h00000a786c253a786c25203d2043414d, /* 2806 */
128'h3025203d20737365726464612043414d, /* 2807 */
128'h3230253a783230253a783230253a7832, /* 2808 */
128'h0000000a2e783230253a783230253a78, /* 2809 */
128'h00007f7c5d5b3f3e3d3c3b3a2c2b2a22, /* 2810 */
128'h007f7c5d5b3f3e3d3c3b3a2e2c2b2a22, /* 2811 */
128'h66656463626139383736353433323130, /* 2812 */
128'h72776f6c2f6372730000000000000000, /* 2813 */
128'h00000000000000632e636d6d5f637369, /* 2814 */
128'h61625f6473203d3d20657361625f6473, /* 2815 */
128'h5f63736972776f6c00726464615f6573, /* 2816 */
128'h000a74756f656d6974207325203a6473, /* 2817 */
128'h616d202c6465766f6d65722064726143, /* 2818 */
128'h6425206f74206465676e616863206b73, /* 2819 */
128'h736e692064726143000000000000000a, /* 2820 */
128'h6e616863206b73616d202c6465747265, /* 2821 */
128'h0000000000000a6425206f7420646567, /* 2822 */
128'h25207461206465746165726320636d6d, /* 2823 */
128'h0000000a7825203d2074736f68202c78, /* 2824 */
128'h0000000000006f4e0000000000736559, /* 2825 */
128'h002020203a434d4d0000000052444420, /* 2826 */
128'h00000000000a7325203a656369766544, /* 2827 */
128'h3a4449207265727574636166756e614d, /* 2828 */
128'h0a7825203a4d454f000000000a782520, /* 2829 */
128'h6325203a656d614e0000000000000000, /* 2830 */
128'h0000000000000a206325632563256325, /* 2831 */
128'h00000a6425203a646565705320737542, /* 2832 */
128'h25203a79746963617061432068676948, /* 2833 */
128'h79746963617061430000000000000a73, /* 2834 */
128'h7464695720737542000000000000203a, /* 2835 */
128'h000000000a73257469622d6425203a68, /* 2836 */
128'h0000007825782520000000203a78250a, /* 2837 */
128'h00000000000064735f63736972776f6c, /* 2838 */
128'h0000000065646f6d206e776f6e6b6e55, /* 2839 */
128'h7830203a726f72724520737574617453, /* 2840 */
128'h2074756f656d69540000000a58383025, /* 2841 */
128'h616572206472616320676e6974696177, /* 2842 */
128'h6c69616620636d6d00000000000a7964, /* 2843 */
128'h6d6320706f747320646e6573206f7420, /* 2844 */
128'h6f6c62203a434d4d0000000000000a64, /* 2845 */
128'h20786c257830207265626d756e206b63, /* 2846 */
128'h6c2578302878616d2073646565637865, /* 2847 */
128'h203d3e20434d4d6500000000000a2978, /* 2848 */
128'h726f6620646572697571657220342e34, /* 2849 */
128'h642072657375206465636e61686e6520, /* 2850 */
128'h000000000000000a6165726120617461, /* 2851 */
128'h757320746f6e2073656f642064726143, /* 2852 */
128'h696e6f697469747261702074726f7070, /* 2853 */
128'h656f64206472614300000000000a676e, /* 2854 */
128'h20434820656e6966656420746f6e2073, /* 2855 */
128'h00000a657a69732070756f7267205057, /* 2856 */
128'h636e61686e6520617461642072657355, /* 2857 */
128'h5720434820746f6e2061657261206465, /* 2858 */
128'h696c6120657a69732070756f72672050, /* 2859 */
128'h72617020692550470000000a64656e67, /* 2860 */
128'h505720434820746f6e206e6f69746974, /* 2861 */
128'h67696c6120657a69732070756f726720, /* 2862 */
128'h656f642064726143000000000a64656e, /* 2863 */
128'h6e652074726f7070757320746f6e2073, /* 2864 */
128'h657475626972747461206465636e6168, /* 2865 */
128'h6e65206c61746f54000000000000000a, /* 2866 */
128'h6563786520657a6973206465636e6168, /* 2867 */
128'h20752528206d756d6978616d20736465, /* 2868 */
128'h656f64206472614300000a297525203e, /* 2869 */
128'h6f682074726f7070757320746f6e2073, /* 2870 */
128'h61702064656c6c6f72746e6f63207473, /* 2871 */
128'h6572206574697277206e6f6974697472, /* 2872 */
128'h6e6974746573207974696c696261696c, /* 2873 */
128'h726c61206472614300000000000a7367, /* 2874 */
128'h64656e6f697469747261702079646165, /* 2875 */
128'h206f6e203a434d4d000000000000000a, /* 2876 */
128'h0000000a746e65736572702064726163, /* 2877 */
128'h73657220746f6e206469642064726143, /* 2878 */
128'h20656761746c6f76206f7420646e6f70, /* 2879 */
128'h00000000000000000a217463656c6573, /* 2880 */
128'h7463656c6573206f7420656c62616e75, /* 2881 */
128'h00000000000000000a65646f6d206120, /* 2882 */
128'h646e756f66206473635f747865206f4e, /* 2883 */
128'h78363025206e614d0000000000000a21, /* 2884 */
128'h000000783430257834302520726e5320, /* 2885 */
128'h00000000632563256325632563256325, /* 2886 */
128'h6167656c20434d4d00000064252e6425, /* 2887 */
128'h636167654c2044530000000000007963, /* 2888 */
128'h6867694820434d4d0000000000000079, /* 2889 */
128'h0000297a484d36322820646565705320, /* 2890 */
128'h35282064656570532068676948204453, /* 2891 */
128'h6867694820434d4d000000297a484d30, /* 2892 */
128'h0000297a484d32352820646565705320, /* 2893 */
128'h7a484d32352820323552444420434d4d, /* 2894 */
128'h31524453205348550000000000000029, /* 2895 */
128'h00000000000000297a484d3532282032, /* 2896 */
128'h7a484d30352820353252445320534855, /* 2897 */
128'h35524453205348550000000000000029, /* 2898 */
128'h000000000000297a484d303031282030, /* 2899 */
128'h7a484d30352820303552444420534855, /* 2900 */
128'h31524453205348550000000000000029, /* 2901 */
128'h0000000000297a484d38303228203430, /* 2902 */
128'h0000297a484d30303228203030325348, /* 2903 */
128'h6f6e2064252065636976654420434d4d, /* 2904 */
128'h00000000000000000a646e756f662074, /* 2905 */
128'h00000000434d4d650000000000004453, /* 2906 */
128'h000000297325282000006425203a7325, /* 2907 */
128'h6e656c20656c69460000000000636d6d, /* 2908 */
128'h000000000000000a6425203d20687467, /* 2909 */
128'h0a7325203d202964252c70252835646d, /* 2910 */
128'h666c652064616f6c0000000000000000, /* 2911 */
128'h000a79726f6d656d20524444206f7420, /* 2912 */
128'h2064656c696166206461657220666c65, /* 2913 */
128'h000000646c252065646f632068746977, /* 2914 */
128'h6f6f7420687461702074736575716552, /* 2915 */
128'h00000000000a646c25202e676e6f6c20, /* 2916 */
128'h732522203a717277000000000000002f, /* 2917 */
128'h0a64253d657a69736b636f6c62202c22, /* 2918 */
128'h20657669656365520000000000000000, /* 2919 */
128'h0000000000000a2e646e6520656c6966, /* 2920 */
128'h656c6c6163207172775f656c646e6168, /* 2921 */
128'h206c6167656c6c4900000000000a2e64, /* 2922 */
128'h0a2e6e6f6974617265706f2050544654, /* 2923 */
128'h75716572206e656c0000000000000000, /* 2924 */
128'h6175746361202c5825203d2064657269, /* 2925 */
128'h000000005c2d2f7c000a7825203d206c, /* 2926 */
128'h20646564616f6c2065687420746f6f42, /* 2927 */
128'h6572646461207461206d6172676f7270, /* 2928 */
128'h000000000000000a2e2e2e7025207373, /* 2929 */
128'h445320746e756f6d206f74206c696146, /* 2930 */
128'h000000000000000a2172657669726420, /* 2931 */
128'h6e69206e69622e746f6f622064616f4c, /* 2932 */
128'h0000000000000a79726f6d656d206f74, /* 2933 */
128'h00000000000000006e69622e746f6f62, /* 2934 */
128'h62206e65706f206f742064656c696146, /* 2935 */
128'h206f74206c6961660000000a21746f6f, /* 2936 */
128'h000000000021656c69662065736f6c63, /* 2937 */
128'h6420746e756f6d75206f74206c696166, /* 2938 */
128'h20746f6f622d750a00000000216b7369, /* 2939 */
128'h67617473207473726966206465736162, /* 2940 */
128'h00000a726564616f6c20746f6f622065, /* 2941 */
128'h696166207325206e6f69747265737361, /* 2942 */
128'h696c202c732520656c6966202c64656c, /* 2943 */
128'h206e6f6974636e7566202c642520656e, /* 2944 */
128'h3a4552554c49414600000000000a7325, /* 2945 */
128'h74612078257830203d21207825783020, /* 2946 */
128'h00000a2e782578302074657366666f20, /* 2947 */
128'h7025203d203270202c7025203d203170, /* 2948 */
128'h2020202020202020000000000000000a, /* 2949 */
128'h08080808080808080000000000202020, /* 2950 */
128'h20676e69747465730000000000080808, /* 2951 */
128'h20676e69747365740000000000007525, /* 2952 */
128'h3a4552554c4941460000000000007525, /* 2953 */
128'h64612064616220656c626973736f7020, /* 2954 */
128'h666f20746120656e696c207373657264, /* 2955 */
128'h00000000000a2e782578302074657366, /* 2956 */
128'h7478656e206f7420676e697070696b53, /* 2957 */
128'h000000000000000a2e2e2e7473657420, /* 2958 */
128'h20202020200808080808080808080808, /* 2959 */
128'h08080808080808080808202020202020, /* 2960 */
128'h00000000000820080000000000000008, /* 2961 */
128'h78302073692065676e61722074736574, /* 2962 */
128'h00000000000a70257830206f74207025, /* 2963 */
128'h000000000075252f00752520706f6f4c, /* 2964 */
128'h6441206b637574530000000000000a3a, /* 2965 */
128'h0000203a732520200000007373657264, /* 2966 */
128'h00000a2e656e6f4400000000000a6b6f, /* 2967 */
128'h4d415244206c6174656d20657261420a, /* 2968 */
128'h65747365746d656d00000a7473657420, /* 2969 */
128'h20302e332e34206e6f69737265762072, /* 2970 */
128'h000000000000000a297469622d642528, /* 2971 */
128'h30322029432820746867697279706f43, /* 2972 */
128'h2073656c7261684320323130322d3130, /* 2973 */
128'h000000000000000a2e6e6f62617a6143, /* 2974 */
128'h74207265646e75206465736e6563694c, /* 2975 */
128'h50206c6172656e654720554e47206568, /* 2976 */
128'h65762065736e6563694c2063696c6275, /* 2977 */
128'h0a2e29796c6e6f282032206e6f697372, /* 2978 */
128'h5f676e696b726f770000000000000000, /* 2979 */
128'h20646c25202c424b6425203d20746573, /* 2980 */
128'h6c25202c736e6f697463757274736e69, /* 2981 */
128'h203d20495043202c73656c6379632064, /* 2982 */
128'h00000000000000000a646c252e646c25, /* 2983 */
128'h46454443424139383736353433323130, /* 2984 */
128'h6f57206f6c6c65480000000000000000, /* 2985 */
128'h205d64255b70777300000a0d21646c72, /* 2986 */
128'h73206863746977530000000a5825203d, /* 2987 */
128'h000a58252c5825203d20676e69747465, /* 2988 */
128'h5825203d2064656573206d6f646e6152, /* 2989 */
128'h0a746f6f62204453000000000000000a, /* 2990 */
128'h6f6f6220495053510000000000000000, /* 2991 */
128'h736574204d4152440000000000000a74, /* 2992 */
128'h6f6f6220505446540000000000000a74, /* 2993 */
128'h65742065686361430000000000000a74, /* 2994 */
128'h00000a0d7061727400000000000a7473, /* 2995 */
128'h00000002464c457fcccccccccccccccd, /* 2996 */
128'h1032547698badcfeefcdab8967452301, /* 2997 */
128'h5851f42d4c957f2d1000000020000000, /* 2998 */
128'haaaaaaaaaaaaaaaa5555555555555555, /* 2999 */
128'h00004b4d47545045000000030f060301, /* 3000 */
128'h000000004300000000000000004b4d47, /* 3001 */
128'h00000000ffffffff0000000000000000, /* 3002 */
128'h0000646d635f6473000000000c000000, /* 3003 */
128'h0000000087feb40800006772615f6473, /* 3004 */
128'h000000000000000000000000cc33aa55, /* 3005 */
128'h00000000000000000000000000000000, /* 3006 */
128'h00000000000000000000000000000000, /* 3007 */
128'h000000002f7c5c2d00000000ffffffff, /* 3008 */
128'hffffffff000000060000000087feb5c0, /* 3009 */
128'h0000000087fe70d20000000000000000, /* 3010 */
128'h00000000000000000000000000000094, /* 3011 */
128'h00000000000000000000000000000000, /* 3012 */
128'h00000000000000000000000000000000, /* 3013 */
128'h00000000000000000000000000000000, /* 3014 */
128'h00000000000000000000000000000000, /* 3015 */
128'h00000000000000000000000000000000, /* 3016 */
128'h00000000000000000000000000000000, /* 3017 */
128'h00000000000000000000000000000000, /* 3018 */
128'h00000000000000000000000000000000, /* 3019 */
128'h00000000000000000000000000000000, /* 3020 */
128'h00000000000000000000000000000000, /* 3021 */
128'h00000000000000000000000000000000, /* 3022 */
128'h00000000000000000000000000000000, /* 3023 */
128'h00000000000000000000000000000000, /* 3024 */
128'h00000000000000000000000000000000, /* 3025 */
128'h00000000000000000000000000000000, /* 3026 */
128'h00000000000000000000000000000000, /* 3027 */
128'h00000000000000000000000000000000, /* 3028 */
128'h00000000000000000000000000000000, /* 3029 */
128'h00000000000000000000000000000000, /* 3030 */
128'h00000000000000000000000000000000, /* 3031 */
128'h00000000000000000000000000000000, /* 3032 */
128'h00000000000000000000000000000000, /* 3033 */
128'h00000000000000000000000000000000, /* 3034 */
128'h00000000000000000000000000000000, /* 3035 */
128'h00000000000000000000000000000000, /* 3036 */
128'h00000000000000000000000000000000, /* 3037 */
128'h00000000000000000000000000000000, /* 3038 */
128'h00000000000000000000000000000000, /* 3039 */
128'h00000000000000000000000000000000, /* 3040 */
128'h00000000000000000000000000000000, /* 3041 */
128'h00000000000000000000000000000000, /* 3042 */
128'h00000000000000000000000000000000, /* 3043 */
128'h00000000000000000000000000000000, /* 3044 */
128'h00000000000000000000000000000000, /* 3045 */
128'h00000000000000000000000000000000, /* 3046 */
128'h00000000000000000000000000000000, /* 3047 */
128'h00000000000000000000000000000000, /* 3048 */
128'h00000000000000000000000000000000, /* 3049 */
128'h00000000000000000000000000000000, /* 3050 */
128'h00000000000000000000000000000000, /* 3051 */
128'h00000000000000000000000000000000, /* 3052 */
128'h00000000000000000000000000000000, /* 3053 */
128'h00000000000000000000000000000000, /* 3054 */
128'h00000000000000000000000000000000, /* 3055 */
128'h00000000000000000000000000000000, /* 3056 */
128'h00000000000000000000000000000000, /* 3057 */
128'h00000000000000000000000000000000, /* 3058 */
128'h00000000000000000000000000000000, /* 3059 */
128'h00000000000000000000000000000000, /* 3060 */
128'h00000000000000000000000000000000, /* 3061 */
128'h00000000000000000000000000000000, /* 3062 */
128'h00000000000000000000000000000000, /* 3063 */
128'h00000000000000000000000000000000, /* 3064 */
128'h00000000000000000000000000000000, /* 3065 */
128'h00000000000000000000000000000000, /* 3066 */
128'h00000000000000000000000000000000, /* 3067 */
128'h00000000000000000000000000000000, /* 3068 */
128'h00000000000000000000000000000000, /* 3069 */
128'h00000000000000000000000000000000, /* 3070 */
128'h00000000000000000000000000000000, /* 3071 */
128'h00000000000000000000000000000000, /* 3072 */
128'h00000000000000000000000000000000, /* 3073 */
128'h00000000000000000000000000000000, /* 3074 */
128'h00000000000000000000000000000000, /* 3075 */
128'h00000000000000000000000000000000, /* 3076 */
128'h00000000000000000000000000000000, /* 3077 */
128'h00000000000000000000000000000000, /* 3078 */
128'h00000000000000000000000000000000, /* 3079 */
128'h00000000000000000000000000000000, /* 3080 */
128'h00000000000000000000000000000000, /* 3081 */
128'h00000000000000000000000000000000, /* 3082 */
128'h00000000000000000000000000000000, /* 3083 */
128'h00000000000000000000000000000000, /* 3084 */
128'h00000000000000000000000000000000, /* 3085 */
128'h00000000000000000000000000000000, /* 3086 */
128'h00000000000000000000000000000000, /* 3087 */
128'h00000000000000000000000000000000, /* 3088 */
128'h00000000000000000000000000000000, /* 3089 */
128'h00000000000000000000000000000000, /* 3090 */
128'h00000000000000000000000000000000, /* 3091 */
128'h00000000000000000000000000000000, /* 3092 */
128'h00000000000000000000000000000000, /* 3093 */
128'h00000000000000000000000000000000, /* 3094 */
128'h00000000000000000000000000000000, /* 3095 */
128'h00000000000000000000000000000000, /* 3096 */
128'h00000000000000000000000000000000, /* 3097 */
128'h00000000000000000000000000000000, /* 3098 */
128'h00000000000000000000000000000000, /* 3099 */
128'h00000000000000000000000000000000, /* 3100 */
128'h00000000000000000000000000000000, /* 3101 */
128'h00000000000000000000000000000000, /* 3102 */
128'h00000000000000000000000000000000, /* 3103 */
128'h00000000000000000000000000000000, /* 3104 */
128'h00000000000000000000000000000000, /* 3105 */
128'h00000000000000000000000000000000, /* 3106 */
128'h00000000000000000000000000000000, /* 3107 */
128'h00000000000000000000000000000000, /* 3108 */
128'h00000000000000000000000000000000, /* 3109 */
128'h00000000000000000000000000000000, /* 3110 */
128'h00000000000000000000000000000000, /* 3111 */
128'h00000000000000000000000000000000, /* 3112 */
128'h00000000000000000000000000000000, /* 3113 */
128'h00000000000000000000000000000000, /* 3114 */
128'h00000000000000000000000000000000, /* 3115 */
128'h00000000000000000000000000000000, /* 3116 */
128'h00000000000000000000000000000000, /* 3117 */
128'h00000000000000000000000000000000, /* 3118 */
128'h00000000000000000000000000000000, /* 3119 */
128'h00000000000000000000000000000000, /* 3120 */
128'h00000000000000000000000000000000, /* 3121 */
128'h00000000000000000000000000000000, /* 3122 */
128'h00000000000000000000000000000000, /* 3123 */
128'h00000000000000000000000000000000, /* 3124 */
128'h00000000000000000000000000000000, /* 3125 */
128'h00000000000000000000000000000000, /* 3126 */
128'h00000000000000000000000000000000, /* 3127 */
128'h00000000000000000000000000000000, /* 3128 */
128'h00000000000000000000000000000000, /* 3129 */
128'h00000000000000000000000000000000, /* 3130 */
128'h00000000000000000000000000000000, /* 3131 */
128'h00000000000000000000000000000000, /* 3132 */
128'h00000000000000000000000000000000, /* 3133 */
128'h00000000000000000000000000000000, /* 3134 */
128'h00000000000000000000000000000000, /* 3135 */
128'h00000000000000000000000000000000, /* 3136 */
128'h00000000000000000000000000000000, /* 3137 */
128'h00000000000000000000000000000000, /* 3138 */
128'h00000000000000000000000000000000, /* 3139 */
128'h00000000000000000000000000000000, /* 3140 */
128'h00000000000000000000000000000000, /* 3141 */
128'h00000000000000000000000000000000, /* 3142 */
128'h00000000000000000000000000000000, /* 3143 */
128'h00000000000000000000000000000000, /* 3144 */
128'h00000000000000000000000000000000, /* 3145 */
128'h00000000000000000000000000000000, /* 3146 */
128'h00000000000000000000000000000000, /* 3147 */
128'h00000000000000000000000000000000, /* 3148 */
128'h00000000000000000000000000000000, /* 3149 */
128'h00000000000000000000000000000000, /* 3150 */
128'h00000000000000000000000000000000, /* 3151 */
128'h00000000000000000000000000000000, /* 3152 */
128'h00000000000000000000000000000000, /* 3153 */
128'h00000000000000000000000000000000, /* 3154 */
128'h00000000000000000000000000000000, /* 3155 */
128'h00000000000000000000000000000000, /* 3156 */
128'h00000000000000000000000000000000, /* 3157 */
128'h00000000000000000000000000000000, /* 3158 */
128'h00000000000000000000000000000000, /* 3159 */
128'h00000000000000000000000000000000, /* 3160 */
128'h00000000000000000000000000000000, /* 3161 */
128'h00000000000000000000000000000000, /* 3162 */
128'h00000000000000000000000000000000, /* 3163 */
128'h00000000000000000000000000000000, /* 3164 */
128'h00000000000000000000000000000000, /* 3165 */
128'h00000000000000000000000000000000, /* 3166 */
128'h00000000000000000000000000000000, /* 3167 */
128'h00000000000000000000000000000000, /* 3168 */
128'h00000000000000000000000000000000, /* 3169 */
128'h00000000000000000000000000000000, /* 3170 */
128'h00000000000000000000000000000000, /* 3171 */
128'h00000000000000000000000000000000, /* 3172 */
128'h00000000000000000000000000000000, /* 3173 */
128'h00000000000000000000000000000000, /* 3174 */
128'h00000000000000000000000000000000, /* 3175 */
128'h00000000000000000000000000000000, /* 3176 */
128'h00000000000000000000000000000000, /* 3177 */
128'h00000000000000000000000000000000, /* 3178 */
128'h00000000000000000000000000000000, /* 3179 */
128'h00000000000000000000000000000000, /* 3180 */
128'h00000000000000000000000000000000, /* 3181 */
128'h00000000000000000000000000000000, /* 3182 */
128'h00000000000000000000000000000000, /* 3183 */
128'h00000000000000000000000000000000, /* 3184 */
128'h00000000000000000000000000000000, /* 3185 */
128'h00000000000000000000000000000000, /* 3186 */
128'h00000000000000000000000000000000, /* 3187 */
128'h00000000000000000000000000000000, /* 3188 */
128'h00000000000000000000000000000000, /* 3189 */
128'h00000000000000000000000000000000, /* 3190 */
128'h00000000000000000000000000000000, /* 3191 */
128'h00000000000000000000000000000000, /* 3192 */
128'h00000000000000000000000000000000, /* 3193 */
128'h00000000000000000000000000000000, /* 3194 */
128'h00000000000000000000000000000000, /* 3195 */
128'h00000000000000000000000000000000, /* 3196 */
128'h00000000000000000000000000000000, /* 3197 */
128'h00000000000000000000000000000000, /* 3198 */
128'h00000000000000000000000000000000, /* 3199 */
128'h00000000000000000000000000000000, /* 3200 */
128'h00000000000000000000000000000000, /* 3201 */
128'h00000000000000000000000000000000, /* 3202 */
128'h00000000000000000000000000000000, /* 3203 */
128'h00000000000000000000000000000000, /* 3204 */
128'h00000000000000000000000000000000, /* 3205 */
128'h00000000000000000000000000000000, /* 3206 */
128'h00000000000000000000000000000000, /* 3207 */
128'h00000000000000000000000000000000, /* 3208 */
128'h00000000000000000000000000000000, /* 3209 */
128'h00000000000000000000000000000000, /* 3210 */
128'h00000000000000000000000000000000, /* 3211 */
128'h00000000000000000000000000000000, /* 3212 */
128'h00000000000000000000000000000000, /* 3213 */
128'h00000000000000000000000000000000, /* 3214 */
128'h00000000000000000000000000000000, /* 3215 */
128'h00000000000000000000000000000000, /* 3216 */
128'h00000000000000000000000000000000, /* 3217 */
128'h00000000000000000000000000000000, /* 3218 */
128'h00000000000000000000000000000000, /* 3219 */
128'h00000000000000000000000000000000, /* 3220 */
128'h00000000000000000000000000000000, /* 3221 */
128'h00000000000000000000000000000000, /* 3222 */
128'h00000000000000000000000000000000, /* 3223 */
128'h00000000000000000000000000000000, /* 3224 */
128'h00000000000000000000000000000000, /* 3225 */
128'h00000000000000000000000000000000, /* 3226 */
128'h00000000000000000000000000000000, /* 3227 */
128'h00000000000000000000000000000000, /* 3228 */
128'h00000000000000000000000000000000, /* 3229 */
128'h00000000000000000000000000000000, /* 3230 */
128'h00000000000000000000000000000000, /* 3231 */
128'h00000000000000000000000000000000, /* 3232 */
128'h00000000000000000000000000000000, /* 3233 */
128'h00000000000000000000000000000000, /* 3234 */
128'h00000000000000000000000000000000, /* 3235 */
128'h00000000000000000000000000000000, /* 3236 */
128'h00000000000000000000000000000000, /* 3237 */
128'h00000000000000000000000000000000, /* 3238 */
128'h00000000000000000000000000000000, /* 3239 */
128'h00000000000000000000000000000000, /* 3240 */
128'h00000000000000000000000000000000, /* 3241 */
128'h00000000000000000000000000000000, /* 3242 */
128'h00000000000000000000000000000000, /* 3243 */
128'h00000000000000000000000000000000, /* 3244 */
128'h00000000000000000000000000000000, /* 3245 */
128'h00000000000000000000000000000000, /* 3246 */
128'h00000000000000000000000000000000, /* 3247 */
128'h00000000000000000000000000000000, /* 3248 */
128'h00000000000000000000000000000000, /* 3249 */
128'h00000000000000000000000000000000, /* 3250 */
128'h00000000000000000000000000000000, /* 3251 */
128'h00000000000000000000000000000000, /* 3252 */
128'h00000000000000000000000000000000, /* 3253 */
128'h00000000000000000000000000000000, /* 3254 */
128'h00000000000000000000000000000000, /* 3255 */
128'h00000000000000000000000000000000, /* 3256 */
128'h00000000000000000000000000000000, /* 3257 */
128'h00000000000000000000000000000000, /* 3258 */
128'h00000000000000000000000000000000, /* 3259 */
128'h00000000000000000000000000000000, /* 3260 */
128'h00000000000000000000000000000000, /* 3261 */
128'h00000000000000000000000000000000, /* 3262 */
128'h00000000000000000000000000000000, /* 3263 */
128'h00000000000000000000000000000000, /* 3264 */
128'h00000000000000000000000000000000, /* 3265 */
128'h00000000000000000000000000000000, /* 3266 */
128'h00000000000000000000000000000000, /* 3267 */
128'h00000000000000000000000000000000, /* 3268 */
128'h00000000000000000000000000000000, /* 3269 */
128'h00000000000000000000000000000000, /* 3270 */
128'h00000000000000000000000000000000, /* 3271 */
128'h00000000000000000000000000000000, /* 3272 */
128'h00000000000000000000000000000000, /* 3273 */
128'h00000000000000000000000000000000, /* 3274 */
128'h00000000000000000000000000000000, /* 3275 */
128'h00000000000000000000000000000000, /* 3276 */
128'h00000000000000000000000000000000, /* 3277 */
128'h00000000000000000000000000000000, /* 3278 */
128'h00000000000000000000000000000000, /* 3279 */
128'h00000000000000000000000000000000, /* 3280 */
128'h00000000000000000000000000000000, /* 3281 */
128'h00000000000000000000000000000000, /* 3282 */
128'h00000000000000000000000000000000, /* 3283 */
128'h00000000000000000000000000000000, /* 3284 */
128'h00000000000000000000000000000000, /* 3285 */
128'h00000000000000000000000000000000, /* 3286 */
128'h00000000000000000000000000000000, /* 3287 */
128'h00000000000000000000000000000000, /* 3288 */
128'h00000000000000000000000000000000, /* 3289 */
128'h00000000000000000000000000000000, /* 3290 */
128'h00000000000000000000000000000000, /* 3291 */
128'h00000000000000000000000000000000, /* 3292 */
128'h00000000000000000000000000000000, /* 3293 */
128'h00000000000000000000000000000000, /* 3294 */
128'h00000000000000000000000000000000, /* 3295 */
128'h00000000000000000000000000000000, /* 3296 */
128'h00000000000000000000000000000000, /* 3297 */
128'h00000000000000000000000000000000, /* 3298 */
128'h00000000000000000000000000000000, /* 3299 */
128'h00000000000000000000000000000000, /* 3300 */
128'h00000000000000000000000000000000, /* 3301 */
128'h00000000000000000000000000000000, /* 3302 */
128'h00000000000000000000000000000000, /* 3303 */
128'h00000000000000000000000000000000, /* 3304 */
128'h00000000000000000000000000000000, /* 3305 */
128'h00000000000000000000000000000000, /* 3306 */
128'h00000000000000000000000000000000, /* 3307 */
128'h00000000000000000000000000000000, /* 3308 */
128'h00000000000000000000000000000000, /* 3309 */
128'h00000000000000000000000000000000, /* 3310 */
128'h00000000000000000000000000000000, /* 3311 */
128'h00000000000000000000000000000000, /* 3312 */
128'h00000000000000000000000000000000, /* 3313 */
128'h00000000000000000000000000000000, /* 3314 */
128'h00000000000000000000000000000000, /* 3315 */
128'h00000000000000000000000000000000, /* 3316 */
128'h00000000000000000000000000000000, /* 3317 */
128'h00000000000000000000000000000000, /* 3318 */
128'h00000000000000000000000000000000, /* 3319 */
128'h00000000000000000000000000000000, /* 3320 */
128'h00000000000000000000000000000000, /* 3321 */
128'h00000000000000000000000000000000, /* 3322 */
128'h00000000000000000000000000000000, /* 3323 */
128'h00000000000000000000000000000000, /* 3324 */
128'h00000000000000000000000000000000, /* 3325 */
128'h00000000000000000000000000000000, /* 3326 */
128'h00000000000000000000000000000000, /* 3327 */
128'h00000000000000000000000000000000, /* 3328 */
128'h00000000000000000000000000000000, /* 3329 */
128'h00000000000000000000000000000000, /* 3330 */
128'h00000000000000000000000000000000, /* 3331 */
128'h00000000000000000000000000000000, /* 3332 */
128'h00000000000000000000000000000000, /* 3333 */
128'h00000000000000000000000000000000, /* 3334 */
128'h00000000000000000000000000000000, /* 3335 */
128'h00000000000000000000000000000000, /* 3336 */
128'h00000000000000000000000000000000, /* 3337 */
128'h00000000000000000000000000000000, /* 3338 */
128'h00000000000000000000000000000000, /* 3339 */
128'h00000000000000000000000000000000, /* 3340 */
128'h00000000000000000000000000000000, /* 3341 */
128'h00000000000000000000000000000000, /* 3342 */
128'h00000000000000000000000000000000, /* 3343 */
128'h00000000000000000000000000000000, /* 3344 */
128'h00000000000000000000000000000000, /* 3345 */
128'h00000000000000000000000000000000, /* 3346 */
128'h00000000000000000000000000000000, /* 3347 */
128'h00000000000000000000000000000000, /* 3348 */
128'h00000000000000000000000000000000, /* 3349 */
128'h00000000000000000000000000000000, /* 3350 */
128'h00000000000000000000000000000000, /* 3351 */
128'h00000000000000000000000000000000, /* 3352 */
128'h00000000000000000000000000000000, /* 3353 */
128'h00000000000000000000000000000000, /* 3354 */
128'h00000000000000000000000000000000, /* 3355 */
128'h00000000000000000000000000000000, /* 3356 */
128'h00000000000000000000000000000000, /* 3357 */
128'h00000000000000000000000000000000, /* 3358 */
128'h00000000000000000000000000000000, /* 3359 */
128'h00000000000000000000000000000000, /* 3360 */
128'h00000000000000000000000000000000, /* 3361 */
128'h00000000000000000000000000000000, /* 3362 */
128'h00000000000000000000000000000000, /* 3363 */
128'h00000000000000000000000000000000, /* 3364 */
128'h00000000000000000000000000000000, /* 3365 */
128'h00000000000000000000000000000000, /* 3366 */
128'h00000000000000000000000000000000, /* 3367 */
128'h00000000000000000000000000000000, /* 3368 */
128'h00000000000000000000000000000000, /* 3369 */
128'h00000000000000000000000000000000, /* 3370 */
128'h00000000000000000000000000000000, /* 3371 */
128'h00000000000000000000000000000000, /* 3372 */
128'h00000000000000000000000000000000, /* 3373 */
128'h00000000000000000000000000000000, /* 3374 */
128'h00000000000000000000000000000000, /* 3375 */
128'h00000000000000000000000000000000, /* 3376 */
128'h00000000000000000000000000000000, /* 3377 */
128'h00000000000000000000000000000000, /* 3378 */
128'h00000000000000000000000000000000, /* 3379 */
128'h00000000000000000000000000000000, /* 3380 */
128'h00000000000000000000000000000000, /* 3381 */
128'h00000000000000000000000000000000, /* 3382 */
128'h00000000000000000000000000000000, /* 3383 */
128'h00000000000000000000000000000000, /* 3384 */
128'h00000000000000000000000000000000, /* 3385 */
128'h00000000000000000000000000000000, /* 3386 */
128'h00000000000000000000000000000000, /* 3387 */
128'h00000000000000000000000000000000, /* 3388 */
128'h00000000000000000000000000000000, /* 3389 */
128'h00000000000000000000000000000000, /* 3390 */
128'h00000000000000000000000000000000, /* 3391 */
128'h00000000000000000000000000000000, /* 3392 */
128'h00000000000000000000000000000000, /* 3393 */
128'h00000000000000000000000000000000, /* 3394 */
128'h00000000000000000000000000000000, /* 3395 */
128'h00000000000000000000000000000000, /* 3396 */
128'h00000000000000000000000000000000, /* 3397 */
128'h00000000000000000000000000000000, /* 3398 */
128'h00000000000000000000000000000000, /* 3399 */
128'h00000000000000000000000000000000, /* 3400 */
128'h00000000000000000000000000000000, /* 3401 */
128'h00000000000000000000000000000000, /* 3402 */
128'h00000000000000000000000000000000, /* 3403 */
128'h00000000000000000000000000000000, /* 3404 */
128'h00000000000000000000000000000000, /* 3405 */
128'h00000000000000000000000000000000, /* 3406 */
128'h00000000000000000000000000000000, /* 3407 */
128'h00000000000000000000000000000000, /* 3408 */
128'h00000000000000000000000000000000, /* 3409 */
128'h00000000000000000000000000000000, /* 3410 */
128'h00000000000000000000000000000000, /* 3411 */
128'h00000000000000000000000000000000, /* 3412 */
128'h00000000000000000000000000000000, /* 3413 */
128'h00000000000000000000000000000000, /* 3414 */
128'h00000000000000000000000000000000, /* 3415 */
128'h00000000000000000000000000000000, /* 3416 */
128'h00000000000000000000000000000000, /* 3417 */
128'h00000000000000000000000000000000, /* 3418 */
128'h00000000000000000000000000000000, /* 3419 */
128'h00000000000000000000000000000000, /* 3420 */
128'h00000000000000000000000000000000, /* 3421 */
128'h00000000000000000000000000000000, /* 3422 */
128'h00000000000000000000000000000000, /* 3423 */
128'h00000000000000000000000000000000, /* 3424 */
128'h00000000000000000000000000000000, /* 3425 */
128'h00000000000000000000000000000000, /* 3426 */
128'h00000000000000000000000000000000, /* 3427 */
128'h00000000000000000000000000000000, /* 3428 */
128'h00000000000000000000000000000000, /* 3429 */
128'h00000000000000000000000000000000, /* 3430 */
128'h00000000000000000000000000000000, /* 3431 */
128'h00000000000000000000000000000000, /* 3432 */
128'h00000000000000000000000000000000, /* 3433 */
128'h00000000000000000000000000000000, /* 3434 */
128'h00000000000000000000000000000000, /* 3435 */
128'h00000000000000000000000000000000, /* 3436 */
128'h00000000000000000000000000000000, /* 3437 */
128'h00000000000000000000000000000000, /* 3438 */
128'h00000000000000000000000000000000, /* 3439 */
128'h00000000000000000000000000000000, /* 3440 */
128'h00000000000000000000000000000000, /* 3441 */
128'h00000000000000000000000000000000, /* 3442 */
128'h00000000000000000000000000000000, /* 3443 */
128'h00000000000000000000000000000000, /* 3444 */
128'h00000000000000000000000000000000, /* 3445 */
128'h00000000000000000000000000000000, /* 3446 */
128'h00000000000000000000000000000000, /* 3447 */
128'h00000000000000000000000000000000, /* 3448 */
128'h00000000000000000000000000000000, /* 3449 */
128'h00000000000000000000000000000000, /* 3450 */
128'h00000000000000000000000000000000, /* 3451 */
128'h00000000000000000000000000000000, /* 3452 */
128'h00000000000000000000000000000000, /* 3453 */
128'h00000000000000000000000000000000, /* 3454 */
128'h00000000000000000000000000000000, /* 3455 */
128'h00000000000000000000000000000000, /* 3456 */
128'h00000000000000000000000000000000, /* 3457 */
128'h00000000000000000000000000000000, /* 3458 */
128'h00000000000000000000000000000000, /* 3459 */
128'h00000000000000000000000000000000, /* 3460 */
128'h00000000000000000000000000000000, /* 3461 */
128'h00000000000000000000000000000000, /* 3462 */
128'h00000000000000000000000000000000, /* 3463 */
128'h00000000000000000000000000000000, /* 3464 */
128'h00000000000000000000000000000000, /* 3465 */
128'h00000000000000000000000000000000, /* 3466 */
128'h00000000000000000000000000000000, /* 3467 */
128'h00000000000000000000000000000000, /* 3468 */
128'h00000000000000000000000000000000, /* 3469 */
128'h00000000000000000000000000000000, /* 3470 */
128'h00000000000000000000000000000000, /* 3471 */
128'h00000000000000000000000000000000, /* 3472 */
128'h00000000000000000000000000000000, /* 3473 */
128'h00000000000000000000000000000000, /* 3474 */
128'h00000000000000000000000000000000, /* 3475 */
128'h00000000000000000000000000000000, /* 3476 */
128'h00000000000000000000000000000000, /* 3477 */
128'h00000000000000000000000000000000, /* 3478 */
128'h00000000000000000000000000000000, /* 3479 */
128'h00000000000000000000000000000000, /* 3480 */
128'h00000000000000000000000000000000, /* 3481 */
128'h00000000000000000000000000000000, /* 3482 */
128'h00000000000000000000000000000000, /* 3483 */
128'h00000000000000000000000000000000, /* 3484 */
128'h00000000000000000000000000000000, /* 3485 */
128'h00000000000000000000000000000000, /* 3486 */
128'h00000000000000000000000000000000, /* 3487 */
128'h00000000000000000000000000000000, /* 3488 */
128'h00000000000000000000000000000000, /* 3489 */
128'h00000000000000000000000000000000, /* 3490 */
128'h00000000000000000000000000000000, /* 3491 */
128'h00000000000000000000000000000000, /* 3492 */
128'h00000000000000000000000000000000, /* 3493 */
128'h00000000000000000000000000000000, /* 3494 */
128'h00000000000000000000000000000000, /* 3495 */
128'h00000000000000000000000000000000, /* 3496 */
128'h00000000000000000000000000000000, /* 3497 */
128'h00000000000000000000000000000000, /* 3498 */
128'h00000000000000000000000000000000, /* 3499 */
128'h00000000000000000000000000000000, /* 3500 */
128'h00000000000000000000000000000000, /* 3501 */
128'h00000000000000000000000000000000, /* 3502 */
128'h00000000000000000000000000000000, /* 3503 */
128'h00000000000000000000000000000000, /* 3504 */
128'h00000000000000000000000000000000, /* 3505 */
128'h00000000000000000000000000000000, /* 3506 */
128'h00000000000000000000000000000000, /* 3507 */
128'h00000000000000000000000000000000, /* 3508 */
128'h00000000000000000000000000000000, /* 3509 */
128'h00000000000000000000000000000000, /* 3510 */
128'h00000000000000000000000000000000, /* 3511 */
128'h00000000000000000000000000000000, /* 3512 */
128'h00000000000000000000000000000000, /* 3513 */
128'h00000000000000000000000000000000, /* 3514 */
128'h00000000000000000000000000000000, /* 3515 */
128'h00000000000000000000000000000000, /* 3516 */
128'h00000000000000000000000000000000, /* 3517 */
128'h00000000000000000000000000000000, /* 3518 */
128'h00000000000000000000000000000000, /* 3519 */
128'h00000000000000000000000000000000, /* 3520 */
128'h00000000000000000000000000000000, /* 3521 */
128'h00000000000000000000000000000000, /* 3522 */
128'h00000000000000000000000000000000, /* 3523 */
128'h00000000000000000000000000000000, /* 3524 */
128'h00000000000000000000000000000000, /* 3525 */
128'h00000000000000000000000000000000, /* 3526 */
128'h00000000000000000000000000000000, /* 3527 */
128'h00000000000000000000000000000000, /* 3528 */
128'h00000000000000000000000000000000, /* 3529 */
128'h00000000000000000000000000000000, /* 3530 */
128'h00000000000000000000000000000000, /* 3531 */
128'h00000000000000000000000000000000, /* 3532 */
128'h00000000000000000000000000000000, /* 3533 */
128'h00000000000000000000000000000000, /* 3534 */
128'h00000000000000000000000000000000, /* 3535 */
128'h00000000000000000000000000000000, /* 3536 */
128'h00000000000000000000000000000000, /* 3537 */
128'h00000000000000000000000000000000, /* 3538 */
128'h00000000000000000000000000000000, /* 3539 */
128'h00000000000000000000000000000000, /* 3540 */
128'h00000000000000000000000000000000, /* 3541 */
128'h00000000000000000000000000000000, /* 3542 */
128'h00000000000000000000000000000000, /* 3543 */
128'h00000000000000000000000000000000, /* 3544 */
128'h00000000000000000000000000000000, /* 3545 */
128'h00000000000000000000000000000000, /* 3546 */
128'h00000000000000000000000000000000, /* 3547 */
128'h00000000000000000000000000000000, /* 3548 */
128'h00000000000000000000000000000000, /* 3549 */
128'h00000000000000000000000000000000, /* 3550 */
128'h00000000000000000000000000000000, /* 3551 */
128'h00000000000000000000000000000000, /* 3552 */
128'h00000000000000000000000000000000, /* 3553 */
128'h00000000000000000000000000000000, /* 3554 */
128'h00000000000000000000000000000000, /* 3555 */
128'h00000000000000000000000000000000, /* 3556 */
128'h00000000000000000000000000000000, /* 3557 */
128'h00000000000000000000000000000000, /* 3558 */
128'h00000000000000000000000000000000, /* 3559 */
128'h00000000000000000000000000000000, /* 3560 */
128'h00000000000000000000000000000000, /* 3561 */
128'h00000000000000000000000000000000, /* 3562 */
128'h00000000000000000000000000000000, /* 3563 */
128'h00000000000000000000000000000000, /* 3564 */
128'h00000000000000000000000000000000, /* 3565 */
128'h00000000000000000000000000000000, /* 3566 */
128'h00000000000000000000000000000000, /* 3567 */
128'h00000000000000000000000000000000, /* 3568 */
128'h00000000000000000000000000000000, /* 3569 */
128'h00000000000000000000000000000000, /* 3570 */
128'h00000000000000000000000000000000, /* 3571 */
128'h00000000000000000000000000000000, /* 3572 */
128'h00000000000000000000000000000000, /* 3573 */
128'h00000000000000000000000000000000, /* 3574 */
128'h00000000000000000000000000000000, /* 3575 */
128'h00000000000000000000000000000000, /* 3576 */
128'h00000000000000000000000000000000, /* 3577 */
128'h00000000000000000000000000000000, /* 3578 */
128'h00000000000000000000000000000000, /* 3579 */
128'h00000000000000000000000000000000, /* 3580 */
128'h00000000000000000000000000000000, /* 3581 */
128'h00000000000000000000000000000000, /* 3582 */
128'h00000000000000000000000000000000, /* 3583 */
128'h00000000000000000000000000000000, /* 3584 */
128'h00000000000000000000000000000000, /* 3585 */
128'h00000000000000000000000000000000, /* 3586 */
128'h00000000000000000000000000000000, /* 3587 */
128'h00000000000000000000000000000000, /* 3588 */
128'h00000000000000000000000000000000, /* 3589 */
128'h00000000000000000000000000000000, /* 3590 */
128'h00000000000000000000000000000000, /* 3591 */
128'h00000000000000000000000000000000, /* 3592 */
128'h00000000000000000000000000000000, /* 3593 */
128'h00000000000000000000000000000000, /* 3594 */
128'h00000000000000000000000000000000, /* 3595 */
128'h00000000000000000000000000000000, /* 3596 */
128'h00000000000000000000000000000000, /* 3597 */
128'h00000000000000000000000000000000, /* 3598 */
128'h00000000000000000000000000000000, /* 3599 */
128'h00000000000000000000000000000000, /* 3600 */
128'h00000000000000000000000000000000, /* 3601 */
128'h00000000000000000000000000000000, /* 3602 */
128'h00000000000000000000000000000000, /* 3603 */
128'h00000000000000000000000000000000, /* 3604 */
128'h00000000000000000000000000000000, /* 3605 */
128'h00000000000000000000000000000000, /* 3606 */
128'h00000000000000000000000000000000, /* 3607 */
128'h00000000000000000000000000000000, /* 3608 */
128'h00000000000000000000000000000000, /* 3609 */
128'h00000000000000000000000000000000, /* 3610 */
128'h00000000000000000000000000000000, /* 3611 */
128'h00000000000000000000000000000000, /* 3612 */
128'h00000000000000000000000000000000, /* 3613 */
128'h00000000000000000000000000000000, /* 3614 */
128'h00000000000000000000000000000000, /* 3615 */
128'h00000000000000000000000000000000, /* 3616 */
128'h00000000000000000000000000000000, /* 3617 */
128'h00000000000000000000000000000000, /* 3618 */
128'h00000000000000000000000000000000, /* 3619 */
128'h00000000000000000000000000000000, /* 3620 */
128'h00000000000000000000000000000000, /* 3621 */
128'h00000000000000000000000000000000, /* 3622 */
128'h00000000000000000000000000000000, /* 3623 */
128'h00000000000000000000000000000000, /* 3624 */
128'h00000000000000000000000000000000, /* 3625 */
128'h00000000000000000000000000000000, /* 3626 */
128'h00000000000000000000000000000000, /* 3627 */
128'h00000000000000000000000000000000, /* 3628 */
128'h00000000000000000000000000000000, /* 3629 */
128'h00000000000000000000000000000000, /* 3630 */
128'h00000000000000000000000000000000, /* 3631 */
128'h00000000000000000000000000000000, /* 3632 */
128'h00000000000000000000000000000000, /* 3633 */
128'h00000000000000000000000000000000, /* 3634 */
128'h00000000000000000000000000000000, /* 3635 */
128'h00000000000000000000000000000000, /* 3636 */
128'h00000000000000000000000000000000, /* 3637 */
128'h00000000000000000000000000000000, /* 3638 */
128'h00000000000000000000000000000000, /* 3639 */
128'h00000000000000000000000000000000, /* 3640 */
128'h00000000000000000000000000000000, /* 3641 */
128'h00000000000000000000000000000000, /* 3642 */
128'h00000000000000000000000000000000, /* 3643 */
128'h00000000000000000000000000000000, /* 3644 */
128'h00000000000000000000000000000000, /* 3645 */
128'h00000000000000000000000000000000, /* 3646 */
128'h00000000000000000000000000000000, /* 3647 */
128'h00000000000000000000000000000000, /* 3648 */
128'h00000000000000000000000000000000, /* 3649 */
128'h00000000000000000000000000000000, /* 3650 */
128'h00000000000000000000000000000000, /* 3651 */
128'h00000000000000000000000000000000, /* 3652 */
128'h00000000000000000000000000000000, /* 3653 */
128'h00000000000000000000000000000000, /* 3654 */
128'h00000000000000000000000000000000, /* 3655 */
128'h00000000000000000000000000000000, /* 3656 */
128'h00000000000000000000000000000000, /* 3657 */
128'h00000000000000000000000000000000, /* 3658 */
128'h00000000000000000000000000000000, /* 3659 */
128'h00000000000000000000000000000000, /* 3660 */
128'h00000000000000000000000000000000, /* 3661 */
128'h00000000000000000000000000000000, /* 3662 */
128'h00000000000000000000000000000000, /* 3663 */
128'h00000000000000000000000000000000, /* 3664 */
128'h00000000000000000000000000000000, /* 3665 */
128'h00000000000000000000000000000000, /* 3666 */
128'h00000000000000000000000000000000, /* 3667 */
128'h00000000000000000000000000000000, /* 3668 */
128'h00000000000000000000000000000000, /* 3669 */
128'h00000000000000000000000000000000, /* 3670 */
128'h00000000000000000000000000000000, /* 3671 */
128'h00000000000000000000000000000000, /* 3672 */
128'h00000000000000000000000000000000, /* 3673 */
128'h00000000000000000000000000000000, /* 3674 */
128'h00000000000000000000000000000000, /* 3675 */
128'h00000000000000000000000000000000, /* 3676 */
128'h00000000000000000000000000000000, /* 3677 */
128'h00000000000000000000000000000000, /* 3678 */
128'h00000000000000000000000000000000, /* 3679 */
128'h00000000000000000000000000000000, /* 3680 */
128'h00000000000000000000000000000000, /* 3681 */
128'h00000000000000000000000000000000, /* 3682 */
128'h00000000000000000000000000000000, /* 3683 */
128'h00000000000000000000000000000000, /* 3684 */
128'h00000000000000000000000000000000, /* 3685 */
128'h00000000000000000000000000000000, /* 3686 */
128'h00000000000000000000000000000000, /* 3687 */
128'h00000000000000000000000000000000, /* 3688 */
128'h00000000000000000000000000000000, /* 3689 */
128'h00000000000000000000000000000000, /* 3690 */
128'h00000000000000000000000000000000, /* 3691 */
128'h00000000000000000000000000000000, /* 3692 */
128'h00000000000000000000000000000000, /* 3693 */
128'h00000000000000000000000000000000, /* 3694 */
128'h00000000000000000000000000000000, /* 3695 */
128'h00000000000000000000000000000000, /* 3696 */
128'h00000000000000000000000000000000, /* 3697 */
128'h00000000000000000000000000000000, /* 3698 */
128'h00000000000000000000000000000000, /* 3699 */
128'h00000000000000000000000000000000, /* 3700 */
128'h00000000000000000000000000000000, /* 3701 */
128'h00000000000000000000000000000000, /* 3702 */
128'h00000000000000000000000000000000, /* 3703 */
128'h00000000000000000000000000000000, /* 3704 */
128'h00000000000000000000000000000000, /* 3705 */
128'h00000000000000000000000000000000, /* 3706 */
128'h00000000000000000000000000000000, /* 3707 */
128'h00000000000000000000000000000000, /* 3708 */
128'h00000000000000000000000000000000, /* 3709 */
128'h00000000000000000000000000000000, /* 3710 */
128'h00000000000000000000000000000000, /* 3711 */
128'h00000000000000000000000000000000, /* 3712 */
128'h00000000000000000000000000000000, /* 3713 */
128'h00000000000000000000000000000000, /* 3714 */
128'h00000000000000000000000000000000, /* 3715 */
128'h00000000000000000000000000000000, /* 3716 */
128'h00000000000000000000000000000000, /* 3717 */
128'h00000000000000000000000000000000, /* 3718 */
128'h00000000000000000000000000000000, /* 3719 */
128'h00000000000000000000000000000000, /* 3720 */
128'h00000000000000000000000000000000, /* 3721 */
128'h00000000000000000000000000000000, /* 3722 */
128'h00000000000000000000000000000000, /* 3723 */
128'h00000000000000000000000000000000, /* 3724 */
128'h00000000000000000000000000000000, /* 3725 */
128'h00000000000000000000000000000000, /* 3726 */
128'h00000000000000000000000000000000, /* 3727 */
128'h00000000000000000000000000000000, /* 3728 */
128'h00000000000000000000000000000000, /* 3729 */
128'h00000000000000000000000000000000, /* 3730 */
128'h00000000000000000000000000000000, /* 3731 */
128'h00000000000000000000000000000000, /* 3732 */
128'h00000000000000000000000000000000, /* 3733 */
128'h00000000000000000000000000000000, /* 3734 */
128'h00000000000000000000000000000000, /* 3735 */
128'h00000000000000000000000000000000, /* 3736 */
128'h00000000000000000000000000000000, /* 3737 */
128'h00000000000000000000000000000000, /* 3738 */
128'h00000000000000000000000000000000, /* 3739 */
128'h00000000000000000000000000000000, /* 3740 */
128'h00000000000000000000000000000000, /* 3741 */
128'h00000000000000000000000000000000, /* 3742 */
128'h00000000000000000000000000000000, /* 3743 */
128'h00000000000000000000000000000000, /* 3744 */
128'h00000000000000000000000000000000, /* 3745 */
128'h00000000000000000000000000000000, /* 3746 */
128'h00000000000000000000000000000000, /* 3747 */
128'h00000000000000000000000000000000, /* 3748 */
128'h00000000000000000000000000000000, /* 3749 */
128'h00000000000000000000000000000000, /* 3750 */
128'h00000000000000000000000000000000, /* 3751 */
128'h00000000000000000000000000000000, /* 3752 */
128'h00000000000000000000000000000000, /* 3753 */
128'h00000000000000000000000000000000, /* 3754 */
128'h00000000000000000000000000000000, /* 3755 */
128'h00000000000000000000000000000000, /* 3756 */
128'h00000000000000000000000000000000, /* 3757 */
128'h00000000000000000000000000000000, /* 3758 */
128'h00000000000000000000000000000000, /* 3759 */
128'h00000000000000000000000000000000, /* 3760 */
128'h00000000000000000000000000000000, /* 3761 */
128'h00000000000000000000000000000000, /* 3762 */
128'h00000000000000000000000000000000, /* 3763 */
128'h00000000000000000000000000000000, /* 3764 */
128'h00000000000000000000000000000000, /* 3765 */
128'h00000000000000000000000000000000, /* 3766 */
128'h00000000000000000000000000000000, /* 3767 */
128'h00000000000000000000000000000000, /* 3768 */
128'h00000000000000000000000000000000, /* 3769 */
128'h00000000000000000000000000000000, /* 3770 */
128'h00000000000000000000000000000000, /* 3771 */
128'h00000000000000000000000000000000, /* 3772 */
128'h00000000000000000000000000000000, /* 3773 */
128'h00000000000000000000000000000000, /* 3774 */
128'h00000000000000000000000000000000, /* 3775 */
128'h00000000000000000000000000000000, /* 3776 */
128'h00000000000000000000000000000000, /* 3777 */
128'h00000000000000000000000000000000, /* 3778 */
128'h00000000000000000000000000000000, /* 3779 */
128'h00000000000000000000000000000000, /* 3780 */
128'h00000000000000000000000000000000, /* 3781 */
128'h00000000000000000000000000000000, /* 3782 */
128'h00000000000000000000000000000000, /* 3783 */
128'h00000000000000000000000000000000, /* 3784 */
128'h00000000000000000000000000000000, /* 3785 */
128'h00000000000000000000000000000000, /* 3786 */
128'h00000000000000000000000000000000, /* 3787 */
128'h00000000000000000000000000000000, /* 3788 */
128'h00000000000000000000000000000000, /* 3789 */
128'h00000000000000000000000000000000, /* 3790 */
128'h00000000000000000000000000000000, /* 3791 */
128'h00000000000000000000000000000000, /* 3792 */
128'h00000000000000000000000000000000, /* 3793 */
128'h00000000000000000000000000000000, /* 3794 */
128'h00000000000000000000000000000000, /* 3795 */
128'h00000000000000000000000000000000, /* 3796 */
128'h00000000000000000000000000000000, /* 3797 */
128'h00000000000000000000000000000000, /* 3798 */
128'h00000000000000000000000000000000, /* 3799 */
128'h00000000000000000000000000000000, /* 3800 */
128'h00000000000000000000000000000000, /* 3801 */
128'h00000000000000000000000000000000, /* 3802 */
128'h00000000000000000000000000000000, /* 3803 */
128'h00000000000000000000000000000000, /* 3804 */
128'h00000000000000000000000000000000, /* 3805 */
128'h00000000000000000000000000000000, /* 3806 */
128'h00000000000000000000000000000000, /* 3807 */
128'h00000000000000000000000000000000, /* 3808 */
128'h00000000000000000000000000000000, /* 3809 */
128'h00000000000000000000000000000000, /* 3810 */
128'h00000000000000000000000000000000, /* 3811 */
128'h00000000000000000000000000000000, /* 3812 */
128'h00000000000000000000000000000000, /* 3813 */
128'h00000000000000000000000000000000, /* 3814 */
128'h00000000000000000000000000000000, /* 3815 */
128'h00000000000000000000000000000000, /* 3816 */
128'h00000000000000000000000000000000, /* 3817 */
128'h00000000000000000000000000000000, /* 3818 */
128'h00000000000000000000000000000000, /* 3819 */
128'h00000000000000000000000000000000, /* 3820 */
128'h00000000000000000000000000000000, /* 3821 */
128'h00000000000000000000000000000000, /* 3822 */
128'h00000000000000000000000000000000, /* 3823 */
128'h00000000000000000000000000000000, /* 3824 */
128'h00000000000000000000000000000000, /* 3825 */
128'h00000000000000000000000000000000, /* 3826 */
128'h00000000000000000000000000000000, /* 3827 */
128'h00000000000000000000000000000000, /* 3828 */
128'h00000000000000000000000000000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00000000000000000000000000000000, /* 3840 */
128'h00000000000000000000000000000000, /* 3841 */
128'h00000000000000000000000000000000, /* 3842 */
128'h00000000000000000000000000000000, /* 3843 */
128'h00000000000000000000000000000000, /* 3844 */
128'h00000000000000000000000000000000, /* 3845 */
128'h00000000000000000000000000000000, /* 3846 */
128'h00000000000000000000000000000000, /* 3847 */
128'h00000000000000000000000000000000, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule

