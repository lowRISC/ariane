/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module etherboot (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 5906;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h87fe7046_00000000,
        64'h87fe7084_00000000,
        64'h00000000_ffffffff,
        64'h00000006_00000000,
        64'h87feb1d0_cc33aa55,
        64'h00000000_2f7c5c2d,
        64'h00000000_87feb018,
        64'h00000000_ffffffff,
        64'h00006772_615f6473,
        64'h0000646d_635f6473,
        64'h00000000_0c000000,
        64'h00000000_ffffffff,
        64'h00000000_00000000,
        64'h00000000_30000000,
        64'h00000000_004b4d47,
        64'h00004b4d_47545045,
        64'h00000003_0f060301,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'haaaaaaaa_aaaaaaaa,
        64'h55555555_55555555,
        64'h5851f42d_4c957f2d,
        64'h10000000_20000000,
        64'h10325476_98badcfe,
        64'hefcdab89_67452301,
        64'hcccccccc_cccccccd,
        64'h00000a0d_70617274,
        64'h00000000_000a7473,
        64'h65742065_68636143,
        64'h00000000_00000a74,
        64'h6f6f6220_50544654,
        64'h00000000_00000a74,
        64'h73657420_4d415244,
        64'h00000000_00000000,
        64'h0a746f6f_62204453,
        64'h00000000_0000000a,
        64'h5825203d_20646565,
        64'h73206d6f_646e6152,
        64'h000a5825_2c582520,
        64'h3d20676e_69747465,
        64'h73206863_74697753,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00000000,
        64'h0a646c25_2e646c25,
        64'h203d2049_5043202c,
        64'h73656c63_79632064,
        64'h6c25202c_736e6f69,
        64'h74637572_74736e69,
        64'h20646c25_202c424b,
        64'h6425203d_20746573,
        64'h5f676e69_6b726f77,
        64'h00000000_00000000,
        64'h0a2e2979_6c6e6f28,
        64'h2032206e_6f697372,
        64'h65762065_736e6563,
        64'h694c2063_696c6275,
        64'h50206c61_72656e65,
        64'h4720554e_47206568,
        64'h74207265_646e7520,
        64'h6465736e_6563694c,
        64'h00000000_0000000a,
        64'h2e6e6f62_617a6143,
        64'h2073656c_72616843,
        64'h20323130_322d3130,
        64'h30322029_43282074,
        64'h68676972_79706f43,
        64'h00000000_0000000a,
        64'h29746962_2d642528,
        64'h20302e33_2e34206e,
        64'h6f697372_65762072,
        64'h65747365_746d656d,
        64'h00000a74_73657420,
        64'h4d415244_206c6174,
        64'h656d2065_7261420a,
        64'h00000a2e_656e6f44,
        64'h00000000_000a6b6f,
        64'h0000203a_73252020,
        64'h00000073_73657264,
        64'h6441206b_63757453,
        64'h00000000_00000a3a,
        64'h00000000_0075252f,
        64'h00752520_706f6f4c,
        64'h00000000_000a7025,
        64'h7830206f_74207025,
        64'h78302073_69206567,
        64'h6e617220_74736574,
        64'h00000000_00082008,
        64'h00000000_00000008,
        64'h08080808_08080808,
        64'h08082020_20202020,
        64'h20202020_20080808,
        64'h08080808_08080808,
        64'h00000000_0000000a,
        64'h2e2e2e74_73657420,
        64'h7478656e_206f7420,
        64'h676e6970_70696b53,
        64'h00000000_000a2e78,
        64'h25783020_74657366,
        64'h666f2074_6120656e,
        64'h696c2073_73657264,
        64'h64612064_61622065,
        64'h6c626973_736f7020,
        64'h3a455255_4c494146,
        64'h00000000_00007525,
        64'h20676e69_74736574,
        64'h00000000_00007525,
        64'h20676e69_74746573,
        64'h00000000_00080808,
        64'h08080808_08080808,
        64'h00000000_00202020,
        64'h20202020_20202020,
        64'h00000000_0000000a,
        64'h7025203d_20327020,
        64'h2c702520_3d203170,
        64'h00000a2e_78257830,
        64'h20746573_66666f20,
        64'h74612078_25783020,
        64'h3d212078_25783020,
        64'h3a455255_4c494146,
        64'h00000000_000a7325,
        64'h206e6f69_74636e75,
        64'h66202c64_2520656e,
        64'h696c202c_73252065,
        64'h6c696620_2c64656c,
        64'h69616620_7325206e,
        64'h6f697472_65737361,
        64'h00000a72_6564616f,
        64'h6c20746f_6f622065,
        64'h67617473_20747372,
        64'h69662064_65736162,
        64'h20746f6f_622d750a,
        64'h00000000_5c2d2f7c,
        64'h00000000_64252065,
        64'h646f6320_68746977,
        64'h2064656c_69616620,
        64'h64616572_20666c65,
        64'h000a7972_6f6d656d,
        64'h20524444_206f7420,
        64'h666c6520_64616f6c,
        64'h00000000_00000000,
        64'h0a2e7365_74796220,
        64'h64252066_6f206e69,
        64'h622e746f_6f62206d,
        64'h6f726620_78252073,
        64'h73657264_64612079,
        64'h726f6d65_6d206f74,
        64'h20736574_79622064,
        64'h25206465_64616f4c,
        64'h00000000_216b7369,
        64'h6420746e_756f6d75,
        64'h206f7420_6c696166,
        64'h00000000_0021656c,
        64'h69662065_736f6c63,
        64'h206f7420_6c696166,
        64'h0000000a_21746f6f,
        64'h62206e65_706f206f,
        64'h74206465_6c696146,
        64'h00000000_00000000,
        64'h6e69622e_746f6f62,
        64'h00000000_00000a79,
        64'h726f6d65_6d206f74,
        64'h6e69206e_69622e74,
        64'h6f6f6220_64616f4c,
        64'h00000000_0000000a,
        64'h21726576_69726420,
        64'h44532074_6e756f6d,
        64'h206f7420_6c696146,
        64'h00000000_00000000,
        64'h0a2e6e6f_69746172,
        64'h65706f20_50544654,
        64'h206c6167_656c6c49,
        64'h00000000_000a2e64,
        64'h656c6c61_63207172,
        64'h775f656c_646e6168,
        64'h00000000_00000a2e,
        64'h646e6520_656c6966,
        64'h20657669_65636552,
        64'h00000000_00000000,
        64'h0a64253d_657a6973,
        64'h6b636f6c_62202c22,
        64'h73252220_3a717277,
        64'h00000000_0000002f,
        64'h00000000_000a646c,
        64'h25202e67_6e6f6c20,
        64'h6f6f7420_68746170,
        64'h20747365_75716552,
        64'h00000000_00000000,
        64'h0a732520_3d202964,
        64'h252c7025_2835646d,
        64'h00000000_0000000a,
        64'h6425203d_20687467,
        64'h6e656c20_656c6946,
        64'h00000000_00636d6d,
        64'h00000029_73252820,
        64'h00006425_203a7325,
        64'h00000000_00004453,
        64'h00000000_434d4d65,
        64'h00000000_00000000,
        64'h0a646e75_6f662074,
        64'h6f6e2064_25206563,
        64'h69766544_20434d4d,
        64'h0000297a_484d3030,
        64'h32282030_30325348,
        64'h00000000_00297a48,
        64'h4d383032_28203430,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282030,
        64'h35524444_20534855,
        64'h00000000_0000297a,
        64'h484d3030_31282030,
        64'h35524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282035,
        64'h32524453_20534855,
        64'h00000000_00000029,
        64'h7a484d35_32282032,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d32_35282032,
        64'h35524444_20434d4d,
        64'h0000297a_484d3235,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000029_7a484d30,
        64'h35282064_65657053,
        64'h20686769_48204453,
        64'h0000297a_484d3632,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000000_00000079,
        64'h63616765_4c204453,
        64'h00000000_00007963,
        64'h6167656c_20434d4d,
        64'h00000064_252e6425,
        64'h00000000_63256325,
        64'h63256325_63256325,
        64'h00000078_34302578,
        64'h34302520_726e5320,
        64'h78363025_206e614d,
        64'h00000000_00000a21,
        64'h646e756f_66206473,
        64'h635f7478_65206f4e,
        64'h00000000_00000000,
        64'h0a65646f_6d206120,
        64'h7463656c_6573206f,
        64'h7420656c_62616e75,
        64'h00000000_00000000,
        64'h0a217463_656c6573,
        64'h20656761_746c6f76,
        64'h206f7420_646e6f70,
        64'h73657220_746f6e20,
        64'h64696420_64726143,
        64'h0000000a_746e6573,
        64'h65727020_64726163,
        64'h206f6e20_3a434d4d,
        64'h00000000_0000000a,
        64'h64656e6f_69746974,
        64'h72617020_79646165,
        64'h726c6120_64726143,
        64'h00000000_000a7367,
        64'h6e697474_65732079,
        64'h74696c69_6261696c,
        64'h65722065_74697277,
        64'h206e6f69_74697472,
        64'h61702064_656c6c6f,
        64'h72746e6f_63207473,
        64'h6f682074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000a29_7525203e,
        64'h20752528_206d756d,
        64'h6978616d_20736465,
        64'h65637865_20657a69,
        64'h73206465_636e6168,
        64'h6e65206c_61746f54,
        64'h00000000_0000000a,
        64'h65747562_69727474,
        64'h61206465_636e6168,
        64'h6e652074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0a64656e,
        64'h67696c61_20657a69,
        64'h73207075_6f726720,
        64'h50572043_4820746f,
        64'h6e206e6f_69746974,
        64'h72617020_69255047,
        64'h0000000a_64656e67,
        64'h696c6120_657a6973,
        64'h2070756f_72672050,
        64'h57204348_20746f6e,
        64'h20616572_61206465,
        64'h636e6168_6e652061,
        64'h74616420_72657355,
        64'h00000a65_7a697320,
        64'h70756f72_67205057,
        64'h20434820_656e6966,
        64'h65642074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_000a676e,
        64'h696e6f69_74697472,
        64'h61702074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0000000a,
        64'h61657261_20617461,
        64'h64207265_73752064,
        64'h65636e61_686e6520,
        64'h726f6620_64657269,
        64'h75716572_20342e34,
        64'h203d3e20_434d4d65,
        64'h00000000_000a2978,
        64'h6c257830_2878616d,
        64'h20736465_65637865,
        64'h20786c25_78302072,
        64'h65626d75_6e206b63,
        64'h6f6c6220_3a434d4d,
        64'h00000000_00000a64,
        64'h6d632070_6f747320,
        64'h646e6573_206f7420,
        64'h6c696166_20636d6d,
        64'h00000000_000a7964,
        64'h61657220_64726163,
        64'h20676e69_74696177,
        64'h2074756f_656d6954,
        64'h0000000a_58383025,
        64'h7830203a_726f7272,
        64'h45207375_74617453,
        64'h00000000_65646f6d,
        64'h206e776f_6e6b6e55,
        64'h00000000_00006473,
        64'h5f637369_72776f6c,
        64'h00000078_25782520,
        64'h00000020_3a78250a,
        64'h00000000_0a732574,
        64'h69622d64_25203a68,
        64'h74646957_20737542,
        64'h00000000_0000203a,
        64'h79746963_61706143,
        64'h00000000_00000a73,
        64'h25203a79_74696361,
        64'h70614320_68676948,
        64'h00000a64_25203a64,
        64'h65657053_20737542,
        64'h00000000_00000a20,
        64'h63256325_63256325,
        64'h6325203a_656d614e,
        64'h00000000_00000000,
        64'h0a782520_3a4d454f,
        64'h00000000_0a782520,
        64'h3a444920_72657275,
        64'h74636166_756e614d,
        64'h00000000_000a7325,
        64'h203a6563_69766544,
        64'h00202020_3a434d4d,
        64'h00000000_52444420,
        64'h00000000_00006f4e,
        64'h00000000_00736559,
        64'h0000000a_7825203d,
        64'h2074736f_68202c78,
        64'h25207461_20646574,
        64'h61657263_20636d6d,
        64'h00000000_00000a64,
        64'h25206f74_20646567,
        64'h6e616863_206b7361,
        64'h6d202c64_65747265,
        64'h736e6920_64726143,
        64'h00000000_0000000a,
        64'h6425206f_74206465,
        64'h676e6168_63206b73,
        64'h616d202c_6465766f,
        64'h6d657220_64726143,
        64'h000a7475_6f656d69,
        64'h74207325_203a6473,
        64'h5f637369_72776f6c,
        64'h00726464_615f6573,
        64'h61625f64_73203d3d,
        64'h20657361_625f6473,
        64'h00000000_00000063,
        64'h2e636d6d_5f637369,
        64'h72776f6c_2f637273,
        64'h00000000_00000000,
        64'h66656463_62613938,
        64'h37363534_33323130,
        64'h007f7c5d_5b3f3e3d,
        64'h3c3b3a2e_2c2b2a22,
        64'h00007f7c_5d5b3f3e,
        64'h3d3c3b3a_2c2b2a22,
        64'h00000000_0a2e2e2e,
        64'h20726574_6f6f6220,
        64'h2c657962_646f6f47,
        64'h00000000_000a2e2e,
        64'h2e6d6172_676f7270,
        64'h20646564_616f6c20,
        64'h65687420_746f6f42,
        64'h00000000_00000000,
        64'h0a646c25_203d2073,
        64'h75746174_73207470,
        64'h75727265_746e6920,
        64'h74656e72_65687445,
        64'h0000000a_2e783230,
        64'h253a7832_30253a78,
        64'h3230253a_78323025,
        64'h3a783230_253a7832,
        64'h3025203d_20737365,
        64'h72646461_2043414d,
        64'h00000a78_6c253a78,
        64'h6c25203d_2043414d,
        64'h000a7264_64612043,
        64'h414d2070_75746553,
        64'h0000000a_21747075,
        64'h72726574_6e692064,
        64'h656c646e_61686e75,
        64'h00000000_00000a78,
        64'h25783020_3d206570,
        64'h79745f6f_746f7270,
        64'h00000000_0a297825,
        64'h28206465_74726f70,
        64'h7075736e_75203d20,
        64'h6f746f72_70205049,
        64'h000a5741_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a534c50_4d203d20,
        64'h6f746f72_50205049,
        64'h00000000_000a4554,
        64'h494c5044_55203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505443_53203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a504d4f_43203d20,
        64'h6f746f72_50205049,
        64'h00000000_0000004d,
        64'h00000000_0000000a,
        64'h5041434e_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000a48,
        64'h50544545_42203d20,
        64'h6f746f72_50205049,
        64'h000a5054_4d203d20,
        64'h6f746f72_50205049,
        64'h00000a48_41203d20,
        64'h6f746f72_50205049,
        64'h000a5053_45203d20,
        64'h6f746f72_50205049,
        64'h000a4552_47203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505653_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000036,
        64'h00000000_00000000,
        64'h0a504343_44203d20,
        64'h6f746f72_50205049,
        64'h00000a50_54203d20,
        64'h6f746f72_50205049,
        64'h000a5044_49203d20,
        64'h6f746f72_50205049,
        64'h000a3a73_746e6574,
        64'h6e6f6320_74736574,
        64'h0000000a_3a726564,
        64'h61656820_74736574,
        64'h000a5055_50203d20,
        64'h6f746f72_50205049,
        64'h000a5047_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000054,
        64'h00000000_00000000,
        64'h0a504950_49203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000047,
        64'h00006425_2b544553,
        64'h46464f5f_524c5052,
        64'h00000000_3f3f3f3f,
        64'h00000000_00544553,
        64'h46464f5f_524c5052,
        64'h00000000_00544553,
        64'h46464f5f_44414252,
        64'h00000000_00005445,
        64'h5346464f_5f525352,
        64'h00000000_00544553,
        64'h46464f5f_53434652,
        64'h00544553_46464f5f,
        64'h4c525443_4f49444d,
        64'h00000000_00544553,
        64'h46464f5f_53434654,
        64'h00000000_00544553,
        64'h46464f5f_524c5054,
        64'h00000000_54455346,
        64'h464f5f49_4843414d,
        64'h00000000_54455346,
        64'h464f5f4f_4c43414d,
        64'h00000000_000a3b29,
        64'h78257830_2c302c78,
        64'h25287465_736d656d,
        64'h00000a3b_29782578,
        64'h302c7825_78302c78,
        64'h25287970_636d656d,
        64'h000a7825_203d206c,
        64'h61757463_61202c58,
        64'h25203d20_64657269,
        64'h75716572_206e656c,
        64'h00000020_3a5d6425,
        64'h5b6e6f69_74636553,
        64'h000a7325_20202020,
        64'h00786c6c_2a302520,
        64'h00003a78_6c383025,
        64'h00732542_69632520,
        64'h00000000_00732573,
        64'h65747942_20756c25,
        64'h0073257a_48632520,
        64'h00000000_646c252e,
        64'h00000000_00756c25,
        64'h00000000_00000000,
        64'h73257a48_20756c25,
        64'h00000000_00007325,
        64'h00000000_00732520,
        64'h3a646c69_7542202c,
        64'h00000000_73257325,
        64'h00000000_00000a0a,
        64'h00000058_32302520,
        64'h00000000_0000002e,
        64'h00000000_00006325,
        64'h00000000_00000020,
        64'h20202020_20202020,
        64'h000a5245_46464f5f,
        64'h50434844_20726f66,
        64'h20676e69_74696157,
        64'h00000a73_25203a73,
        64'h25206563_69766564,
        64'h206e6f20_59524556,
        64'h4f435349_44205043,
        64'h48442064_6e657320,
        64'h74276e64_6c756f43,
        64'h000a5832_30253a58,
        64'h3230253a_58323025,
        64'h3a583230_253a5832,
        64'h30253a58_32302520,
        64'h3a204341_4d207325,
        64'h00000000_30687465,
        64'h00000000_000a2973,
        64'h2528726f_72726570,
        64'h000a5952_45564f43,
        64'h5349445f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_0000000a,
        64'h64252065_646f6370,
        64'h6f205043_48442064,
        64'h656c646e_61686e55,
        64'h00000000_0a642520,
        64'h6e6f6974_706f2064,
        64'h656c646e_61686e75,
        64'h00000000_0000000a,
        64'h73252072_6f727245,
        64'h00000000_00000a64,
        64'h65737566_65722073,
        64'h73657264_64612064,
        64'h65747365_75716552,
        64'h00000000_0000000a,
        64'h4b414e20_50434844,
        64'h00000000_0a444550,
        64'h50494b53_204b4341,
        64'h00000a22_73252220,
        64'h3d207265_76726573,
        64'h00000a22_73252220,
        64'h3d206e69_616d6f64,
        64'h00000000_00000000,
        64'h0a642520_3d20656d,
        64'h69742065_7361654c,
        64'h000a6425_2e64252e,
        64'h64252e64_2520203a,
        64'h73736572_64646120,
        64'h6b73616d_2074654e,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h61207265_74756f52,
        64'h00000000_00000000,
        64'h0a64252e_64252e64,
        64'h252e6425_20203a73,
        64'h73657264_64412050,
        64'h49207265_76726553,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h41205049_20746e65,
        64'h696c4320_50434844,
        64'h00000000_0000000a,
        64'h4b434120_50434844,
        64'h0000000a_54534555,
        64'h5145525f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_00000000,
        64'h0a702520_2c726f72,
        64'h7265206c_616e7265,
        64'h746e6920_70636864,
        64'h00000a29_73252c73,
        64'h25287075_6b6f6f6c,
        64'h000a6563_69766564,
        64'h206e776f_6e6b6e75,
        64'h00000000_203a6425,
        64'h20656369_7665440a,
        64'h00203a64_25206563,
        64'h69766564_2073250a,
        64'h00000000_00203a64,
        64'h25206563_69766544,
        64'h00000000_00000000,
        64'h73736572_6464612d,
        64'h63616d2d_6c61636f,
        64'h6c006874_6469772d,
        64'h6f692d67_65720074,
        64'h66696873_2d676572,
        64'h00737470_75727265,
        64'h746e6900_746e6572,
        64'h61702d74_70757272,
        64'h65746e69_00646565,
        64'h70732d74_6e657272,
        64'h75630076_65646e2c,
        64'h76637369_72007974,
        64'h69726f69_72702d78,
        64'h616d2c76_63736972,
        64'h0073656d_616e2d67,
        64'h65720064_65646e65,
        64'h7478652d_73747075,
        64'h72726574_6e690073,
        64'h65676e61_7200656c,
        64'h646e6168_702c7875,
        64'h6e696c00_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h00100000_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_00000064,
        64'h6e727768_2d637369,
        64'h72776f6c_1b000000,
        64'h0e000000_03000000,
        64'h00003030_30303030,
        64'h30344064_6e727768,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h00800000_00000000,
        64'h00000030_00000000,
        64'h67000000_10000000,
        64'h03000000_00007fe3,
        64'h023e1800_47010000,
        64'h06000000_03000000,
        64'h03000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_00636d6d,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_02000000,
        64'h25010000_04000000,
        64'h03000000_02000000,
        64'h14010000_04000000,
        64'h03000000_00000100,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40636d6d,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h04000000_3a010000,
        64'h04000000_03000000,
        64'h02000000_30010000,
        64'h04000000_03000000,
        64'h01000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h00c20100_06010000,
        64'h04000000_03000000,
        64'h80f0fa02_4b000000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000010_00000000,
        64'h67000000_10000000,
        64'h03000000_00303537,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000000,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'hffff0000_01000000,
        64'hca000000_08000000,
        64'h03000000_00333130,
        64'h2d677562_65642c76,
        64'h63736972_1b000000,
        64'h10000000_03000000,
        64'h00003040_72656c6c,
        64'h6f72746e_6f632d67,
        64'h75626564_01000000,
        64'h02000000_02000000,
        64'hbb000000_04000000,
        64'h03000000_02000000,
        64'hb5000000_04000000,
        64'h03000000_03000000,
        64'hfb000000_04000000,
        64'h03000000_07000000,
        64'he8000000_04000000,
        64'h03000000_00000004,
        64'h00000000_0000000c,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h09000000_01000000,
        64'h0b000000_01000000,
        64'hca000000_10000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00000c00,
        64'h00000000_00000002,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_01000000,
        64'h03000000_01000000,
        64'hca000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6e696c63,
        64'h01000000_c3000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000008_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h01000000_bb000000,
        64'h04000000_03000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00007663_73697200,
        64'h656e6169_7261202c,
        64'h7a687465_1b000000,
        64'h13000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha8060000_59010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'he0060000_38000000,
        64'h39080000_edfe0dd0,
        64'h00000000_64726143,
        64'h2d445320_726f6620,
        64'h746f6f62_2d752064,
        64'h6573696d_696e696d,
        64'h20435349_52776f4c,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00020000_00010000,
        64'h0000c000_00008000,
        64'h00006000_00004000,
        64'h00002000_00001000,
        64'h00000800_00000400,
        64'h00000200_00000100,
        64'h00000080_00000040,
        64'h00000020_00000000,
        64'h0bebc200_0c65d400,
        64'h02faf080_05f5e100,
        64'h02faf080_017d7840,
        64'h03197500_03197500,
        64'h02faf080_018cba80,
        64'h017d7840_017d7840,
        64'h00989680_000f4240,
        64'h000186a0_00002710,
        64'h50463c37_322d2823,
        64'h1e19140f_0d0c0a00,
        64'h00000000_00000000,
        64'h00000000_10000000,
        64'h00000001_00000000,
        64'h20000000_00000002,
        64'h00000000_40000000,
        64'h00000005_00000001,
        64'h20000000_00000006,
        64'h00000001_40000000,
        64'h70000000_00000000,
        64'h70000000_00000002,
        64'h70000000_00000004,
        64'h60000000_00000005,
        64'h30000000_00000001,
        64'h30000000_00000003,
        64'h00000000_40050100,
        64'h40050000_40040500,
        64'h40040401_40040400,
        64'h40040300_40040200,
        64'h40040100_40040000,
        64'h00000000_87feb180,
        64'h00000000_87feb168,
        64'h00000000_87feb150,
        64'h00000000_87feb138,
        64'h00000000_87feb120,
        64'h00000000_87feb108,
        64'h00000000_87feb0f0,
        64'h00000000_87feb0d8,
        64'h00000000_87feb0c0,
        64'h00000000_87feb0a8,
        64'h00000000_87feb098,
        64'h00000000_87feb088,
        64'hffffbd72_ffffbd72,
        64'hffffbd72_ffffbd72,
        64'hffffbd6e_ffffbd6a,
        64'hffffbd6a_ffffbd44,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_87fe4cf8,
        64'h00000000_87fe4a9a,
        64'h00000000_87fe4e8c,
        64'h00646374_65675f63,
        64'h6d6d5f64_72616f62,
        64'h00000002_0000ffff,
        64'h004c4b40_004c4b40,
        64'h00300000_20000000,
        64'h00000000_87fe9a88,
        64'h00000000_87fead70,
        64'h00717269_5f646e65,
        64'h5f617461_645f6473,
        64'h5f637369_72776f6c,
        64'h00000000_00007172,
        64'h695f646d_635f6473,
        64'h5f637369_72776f6c,
        64'h00007172_695f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0067616c,
        64'h665f7470_75727265,
        64'h746e695f_74696177,
        64'h5f637369_72776f6c,
        64'h00000000_646d635f,
        64'h74726174_735f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0000006e,
        64'h655f7172_695f6473,
        64'h00000000_00007475,
        64'h6f656d69_745f6473,
        64'h00000000_0000657a,
        64'h69736b6c_625f6473,
        64'h00000000_00000074,
        64'h6e636b6c_625f6473,
        64'h00000000_00000000,
        64'h74657365_725f6473,
        64'h00000000_74726174,
        64'h735f646d_635f6473,
        64'h00000000_0000676e,
        64'h69747465_735f6473,
        64'h00000000_00007669,
        64'h645f6b6c_635f6473,
        64'h00000000_00000000,
        64'h6e67696c_615f6473,
        64'h00000000_00006465,
        64'h6c5f7465_735f6473,
        64'h5f637369_72776f6c,
        64'h09020b04_0d060f08,
        64'h010a030c_050e0700,
        64'h020f0c09_0603000d,
        64'h0a070401_0e0b0805,
        64'h0c07020d_08030e09,
        64'h040f0a05_000b0601,
        64'heb86d391_2ad7d2bb,
        64'hbd3af235_f7537e82,
        64'h4e0811a1_a3014314,
        64'hfe2ce6e0_6fa87e4f,
        64'h85845dd1_ffeff47d,
        64'h8f0ccc92_655b59c3,
        64'hfc93a039_ab9423a7,
        64'h432aff97_f4292244,
        64'hc4ac5665_1fa27cf8,
        64'he6db99e5_d9d4d039,
        64'h04881d05_d4ef3085,
        64'heaa127fa_289b7ec6,
        64'hbebfbc70_f6bb4b60,
        64'h4bdecfa9_a4beea44,
        64'hfde5380c_6d9d6122,
        64'h8771f681_fffa3942,
        64'h8d2a4c8a_676f02d9,
        64'hfcefa3f8_a9e3e905,
        64'h455a14ed_f4d50d87,
        64'hc33707d6_21e1cde6,
        64'he7d3fbc8_d8a1e681,
        64'h02441453_d62f105d,
        64'he9b6c7aa_265e5a51,
        64'hc040b340_f61e2562,
        64'h49b40821_a679438e,
        64'hfd987193_6b901122,
        64'h895cd7be_ffff5bb1,
        64'h8b44f7af_698098d8,
        64'hfd469501_a8304613,
        64'h4787c62a_f57c0faf,
        64'hc1bdceee_242070db,
        64'he8c7b756_d76aa478,
        64'h02020202_02020202,
        64'h10020202_02020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02010101_01010101,
        64'h10010101_01010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h08101010_10020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02424242_42424210,
        64'h10101010_10010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h01414141_41414110,
        64'h10101010_10100404,
        64'h04040404_04040404,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h08080808_08080808,
        64'h08080808_08080808,
        64'h08082828_28282808,
        64'h08080808_08080808,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h0000b7e9_ee5ff0ef,
        64'h96cfc0ef_0e450513,
        64'h00002517_bff1f7af,
        64'h80ef97ef_c0ef0e65,
        64'h05130000_2517b7fd,
        64'he0dff0ef_990fc0ef,
        64'h0e850513_00002517,
        64'ha001bfdf_e0ef8522,
        64'h9a4fc0ef_0ec50513,
        64'h00002517_00e78c63,
        64'h470504e7_8163470d,
        64'h02e78b63_47090064,
        64'h57930ff4_7413fd39,
        64'h1de39cef_c0ef8552,
        64'h488c0004_a8239daf,
        64'hc0ef8622_24014480,
        64'h448cc09c_09058556,
        64'h0007c783_016907b3,
        64'h4991122a_0a130000,
        64'h2a17112a_8a930000,
        64'h2a974000_04b72e6b,
        64'h0b130000_2b174901,
        64'hb33fe0ef_11c50513,
        64'h00002517_b0dfe0ef,
        64'hf822e05a_e456e852,
        64'hec4ef04a_f426fc06,
        64'h7139b55f_e06f1be5,
        64'h05130000_25178082,
        64'h4b880007_a8234000,
        64'h07b78082_47884000,
        64'h07b78082_c3884000,
        64'h07b7bff1_f5dff0ef,
        64'h4541f63f_f0ef4521,
        64'hf69ff0ef_4511f6ff,
        64'hf0ef4509_f75ff0ef,
        64'h4505f7bf_f0ef4501,
        64'he4061141_bf51c000,
        64'h28f3c020_26f3fac7,
        64'h10e3a96f_c06f1565,
        64'h05130000_251702a7,
        64'h473302a7_67b302b3,
        64'h45bb02c7_47334000,
        64'h059302a6_87334116,
        64'h86b33e80_0513c000,
        64'h26f38e15_c0202673,
        64'h02b71d63_2705fe08,
        64'h13e397aa_387d0007,
        64'h802397aa_00078023,
        64'h97aa0007_802397aa,
        64'h00078023_40000813,
        64'h87f245a9_01f61e13,
        64'h46814881_470100c5,
        64'h131b4605_80828082,
        64'h614569a2_694264e2,
        64'h740270a2_ff2417e3,
        64'he6dff0ef_24050135,
        64'h85334605_46850084,
        64'h95b34979_01f49993,
        64'h4441b36f_c0ef4485,
        64'he7050513_00002517,
        64'hb44fc0ef_1bc50513,
        64'h00002517_b50fc0ef,
        64'h19850513_00002517,
        64'hb5cfc0ef_17c50513,
        64'h00002517_04000593,
        64'hc8bfe0ef_e44ee84a,
        64'hec26f022_f40617e5,
        64'h05130000_25177179,
        64'hbfa10485_b88fc0ef,
        64'hec050513_00002517,
        64'hb7e94a89_b98fc0ef,
        64'h19050513_00002517,
        64'h97828522_85ce6642,
        64'h008a3783_bb0fc0ef,
        64'h1a050513_00002517,
        64'hc58d000a_358302f7,
        64'h49636762_010a2783,
        64'hbccfc0ef_856eed15,
        64'h920ff0ef_852265a2,
        64'hbdcfc0ef_856a85e6,
        64'hbe4fc0ef_8562beaf,
        64'hc0ef855e_85ca0009,
        64'h0663bf6f_c0ef855a,
        64'h85a68082_61497da2,
        64'h7d427ce2_6c066ba6,
        64'h6b466ae6_7a0679a6,
        64'h794674e6_8556640a,
        64'h60aac1ef_c0ef21e5,
        64'h05130000_25170299,
        64'h7863aeaa_0a130000,
        64'h3a1722ad_8d930000,
        64'h2d9722ad_0d130000,
        64'h2d17222c_8c930000,
        64'h2c97222c_0c130000,
        64'h2c17222b_8b930000,
        64'h2b97222b_0b130000,
        64'h2b174485_4a81e43e,
        64'h99a20034_d793e83e,
        64'h0014d993_0044d793,
        64'hc7cfc0ef_ec36e506,
        64'hf46ef86a_fc66e0e2,
        64'he4dee8da_ecd6f0d2,
        64'hf4ce23a5_05130000,
        64'h251785aa_962a84ae,
        64'h842afca6_e122fff5,
        64'h86138932_f8ca7175,
        64'h80826505_b789547d,
        64'hbf290d85_ee5fe0ef,
        64'h0007c503_97ea8b8d,
        64'h00078b1b_001b079b,
        64'hef9fe0ef_4521ef91,
        64'h034df7b3_00f69323,
        64'h93c117c2_0064d783,
        64'h00f69223_93c117c2,
        64'h0044d783_00f69123,
        64'h93c117c2_0024d783,
        64'h00f69023_93c117c2,
        64'h0004d783_e38866c2,
        64'h67e2bea7_b9230000,
        64'h37978d41_91011402,
        64'h15028c51_8d590106,
        64'h161b0105_151b6702,
        64'h662287ef_e0efe02a,
        64'h884fe0ef_e42a88af,
        64'he0ef842a_890fe0ef,
        64'he836ec3e_b7758c4a,
        64'h8bce4a85_80826149,
        64'h7da27d42_7ce26c06,
        64'h6ba66b46_6ae67a06,
        64'h79a67946_74e6640a,
        64'h60aa8522_d78fc0ef,
        64'h31850513_00002517,
        64'h020a8863_e579842a,
        64'ha82ff0ef_854a85ce,
        64'h866e059d_956397de,
        64'h00fc06b3_003d9793,
        64'h4d818c4e_8bca67ed,
        64'h0d130000_2d179c4a,
        64'h0a13c924_84930000,
        64'h34974a81_fe5fe0ef,
        64'h4b018cb2_f46ee122,
        64'he506f86a_fc66e0e2,
        64'he4dee8da_ecd6fca6,
        64'h6a050200_051389ae,
        64'h892af0d2_f4cef8ca,
        64'h7175bfa1_547dbf0d,
        64'h0d8581af_f0ef0007,
        64'hc50397e6_8b8d0007,
        64'h8a9b001a_879b82ef,
        64'hf0ef4521_ef910ba1,
        64'h033df7b3_ffa795e3,
        64'h00d60023_0ff6f693,
        64'h078500fb_86330006,
        64'hc6830187_86b34781,
        64'he288d0a7_b5230000,
        64'h37978d41_66e29101,
        64'h14021502_8c510106,
        64'h161b8d5d_0105151b,
        64'h664267a2_9a0fe0ef,
        64'he42a9a6f_e0efe82a,
        64'h9acfe0ef_842a9b2f,
        64'he0efec36_b7758ba6,
        64'h8b4a4a05_80826149,
        64'h7da27d42_7ce26c06,
        64'h6ba66b46_6ae67a06,
        64'h79a67946_74e6640a,
        64'h60aa8522_e98fc0ef,
        64'h43850513_00002517,
        64'h020a0863_ed45842a,
        64'hba2ff0ef_852685ca,
        64'h866e04fd_956396da,
        64'h003d9693_67824d21,
        64'h4d818bca_8b2679ec,
        64'h8c930000_2c979c49,
        64'h8993daac_0c130000,
        64'h3c174a01_904ff0ef,
        64'h4a81e032_f46ef86a,
        64'he122e506_fc66e0e2,
        64'he4dee8da_ecd6f0d2,
        64'h69850200_0513892e,
        64'h84aaf4ce_f8cafca6,
        64'h7175b7e9_5b7db749,
        64'h060500b8_3023e30c,
        64'h85d6e111_85e20016,
        64'h75138082_61096de2,
        64'h7d027ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_855a7446,
        64'h70e6f46f_c0ef4be5,
        64'h05130000_2517fafb,
        64'h90e30400_07932b85,
        64'hfbb41be3_8c562405,
        64'he9318b2a_c5eff0ef,
        64'h854a85ce_6622f72f,
        64'hc0ef856a_85daf7af,
        64'hc0efe432_855206f6,
        64'h1063974e_00e90833,
        64'h00361713_67824601,
        64'hfffc4a93_f98fc0ef,
        64'h856685da_00848b3b,
        64'hfa4fc0ef_85524401,
        64'h003b949b_01779c33,
        64'h47854da1_4c4d0d13,
        64'h00002d17_4bcc8c93,
        64'h00002c97_4b4a0a13,
        64'h00002a17_fd0fc0ef,
        64'h4b81e032_89aef862,
        64'he0dae4d6_f4a6f8a2,
        64'hfc86ec6e_f06af466,
        64'hfc5ee8d2_ecce4ce5,
        64'h05130000_2517892a,
        64'hf0ca7119_bf755dfd,
        64'hbfc585ba_fe081be3,
        64'h85c6b761_0605e10c,
        64'he28c85be_00081363,
        64'h859a008b_ea630016,
        64'h78138082_61096de2,
        64'h7d027ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_856e7446,
        64'h70e6847f_c0ef5be5,
        64'h05130000_2517f8f4,
        64'h1be30800_07932405,
        64'hed298daa_d56ff0ef,
        64'h852685ca_662286bf,
        64'hc0ef8566_85a2873f,
        64'hc0efe432_854e0546,
        64'h1c6396ca_00d48533,
        64'h00361693_4601fff7,
        64'hc313fff7_48938fd5,
        64'h008d16b3_00fd17b3,
        64'h0024079b_8f5d00ed,
        64'h173300fd_17b3408b,
        64'h07bb408a_873b8b3f,
        64'hc0ef8562_85a28bbf,
        64'hc0ef854e_5ccc8c93,
        64'h00002c97_03f00b93,
        64'h08100b13_4d0507f0,
        64'h0a935d2c_0c130000,
        64'h2c175ca9_89930000,
        64'h29978e7f_c0ef4401,
        64'h8a32892e_ec6efc86,
        64'hf06af466_f862fc5e,
        64'he0dae4d6_e8d2ecce,
        64'hf0caf8a2_5e450513,
        64'h00002517_84aaf4a6,
        64'h7119b7f1_5dfdbfe5,
        64'he19ce31c_bf610605,
        64'he194e314_008c6663,
        64'h80826109_6de27d02,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e67906,
        64'h74a6856e_744670e6,
        64'h94dfc0ef_6c450513,
        64'h00002517_fb5417e3,
        64'h2405e139_8daae58f,
        64'hf0ef8526_85ca6622,
        64'h96dfc0ef_856a85a2,
        64'h975fc0ef_e4328552,
        64'h05661a63_974a00e4,
        64'h85b30036_17134601,
        64'hfff6c693_fff7c793,
        64'h008996b3_00f997b3,
        64'h408b87bb_9a1fc0ef,
        64'h856685a2_9a9fc0ef,
        64'h85520800_0a936bed,
        64'h0d130000_2d1703f0,
        64'h0c134985_07f00b93,
        64'h6c0c8c93_00002c97,
        64'h6b8a0a13_00002a17,
        64'h9d5fc0ef_44018b32,
        64'h892eec6e_fc86f06a,
        64'hf466f862_fc5ee0da,
        64'he4d6e8d2_eccef0ca,
        64'hf8a26d25_05130000,
        64'h251784aa_f4a67119,
        64'hb7f15dfd_bfe5e298,
        64'he398bf61_0605e28c,
        64'he38c008c_66638082,
        64'h61096de2_7d027ca2,
        64'h7c427be2_6b066aa6,
        64'h6a4669e6_790674a6,
        64'h856e7446_70e6a3bf,
        64'hc0ef7b25_05130000,
        64'h2517fb54_1be32405,
        64'he1398daa_f46ff0ef,
        64'h852685ca_6622a5bf,
        64'hc0ef856a_85a2a63f,
        64'hc0efe432_85520566,
        64'h1a6397ca_00f486b3,
        64'h00361793_46010089,
        64'h95b300e9_9733408b,
        64'h873ba87f_c0ef8566,
        64'h85a2a8ff_c0ef8552,
        64'h08000a93_7a4d0d13,
        64'h00002d17_03f00c13,
        64'h498507f0_0b937a6c,
        64'h8c930000_2c9779ea,
        64'h0a130000_2a17abbf,
        64'hc0ef4401_8b32892e,
        64'hec6efc86_f06af466,
        64'hf862fc5e_e0dae4d6,
        64'he8d2ecce_f0caf8a2,
        64'h7b850513_00002517,
        64'h84aaf4a6_7119bff1,
        64'h59fdb74d_0605e29c,
        64'he31c8082_61256c42,
        64'h6be27b02_7aa27a42,
        64'h79e26906_64a6854e,
        64'h644660e6_b11fc0ef,
        64'h88850513_00003517,
        64'hf94c19e3_0c05e91d,
        64'h89aa81df_f0ef8522,
        64'h85a66622_b31fc0ef,
        64'h855e85ce_b39fc0ef,
        64'he432854a_05561763,
        64'h972600e4_06b30036,
        64'h17134601_8fd9038c,
        64'h17138fd9_030c1713,
        64'h8fd9028c_17138fd9,
        64'h020c1713_8fd9018c,
        64'h17130187_e7b38fd9,
        64'h010c1793_008c1713,
        64'hb7dfc0ef_855a85ce,
        64'h000c099b_b89fc0ef,
        64'h854a1000_0a1389eb,
        64'h8b930000_3b97896b,
        64'h0b130000_3b1788e9,
        64'h09130000_3917babf,
        64'hc0ef4c01_8ab284ae,
        64'hfc4eec86_e862ec5e,
        64'hf05af456_f852e0ca,
        64'he4a68a25_05130000,
        64'h3517842a_e8a2711d,
        64'hb7e15d7d_b7790605,
        64'he198e398_872ac291,
        64'h876a0016_7693bf49,
        64'h000b3d03_80826165,
        64'h6d426ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h694664e6_856a7406,
        64'h70a6c0ff_c0ef9865,
        64'h05130000_3517fb44,
        64'h1ae32405_e5298d2a,
        64'h91bff0ef_852685ca,
        64'h6622c2ff_c0ef8566,
        64'h85a2c37f_c0efe432,
        64'h854e0556_1c6397ca,
        64'h00f485b3_00361793,
        64'hfffd4513_4601c53f,
        64'hc0ef8562_85a2000b,
        64'hbd03cba5_00147793,
        64'hc65fc0ef_854e0400,
        64'h0a1397ac_8c930000,
        64'h3c97972c_0c130000,
        64'h3c17c3ab_8b930000,
        64'h3b97c3ab_0b130000,
        64'h3b1797a9_89930000,
        64'h3997c97f_c0ef4401,
        64'h8ab2892e_e86af486,
        64'hec66f062_f45ef85a,
        64'hfc56e0d2_e4cee8ca,
        64'hf0a29925_05130000,
        64'h351784aa_eca67159,
        64'hbfc154fd_bf590605,
        64'he198e398_8726c291,
        64'h87660016_76938082,
        64'h61656ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h64e66946_85267406,
        64'h70a6cf7f_c0efa6e5,
        64'h05130000_3517fb54,
        64'h1be32405_e12984aa,
        64'ha03ff0ef_854a85ce,
        64'h6622d17f_c0ef8562,
        64'h85a2d1ff_c0efe432,
        64'h85520566_186397ce,
        64'h00f905b3_00361793,
        64'h14fd4601_40900cb3,
        64'hd3dfc0ef_8885855e,
        64'h85a2fff4_4493d4bf,
        64'hc0ef8552_04000a93,
        64'ha60c0c13_00003c17,
        64'ha58b8b93_00003b97,
        64'ha50a0a13_00003a17,
        64'hd6dfc0ef_44018b32,
        64'h89aeec66_eca6f486,
        64'hf062f45e_f85afc56,
        64'he0d2e4ce_f0a2a665,
        64'h05130000_3517892a,
        64'he8ca7159_bfc90705,
        64'h00a83023_e28800f7,
        64'h0533a9df_f06f6121,
        64'h863a69e2_854e7902,
        64'h74a270e2_744200c7,
        64'h1c6396ae_00d98833,
        64'h00371693_47018fc5,
        64'h90811782_65a26602,
        64'h14828fc1_8cc90109,
        64'h179b0105_151b92bf,
        64'he0ef84aa_931fe0ef,
        64'h892a937f_e0ef842a,
        64'h93dfe0ef_89aaec4e,
        64'hf04af426_f822fc06,
        64'he032e42e_7139b7f1,
        64'h00e83023_8f690008,
        64'h3703e314_8ee90785,
        64'h6314b15f_f06f6121,
        64'h863e69e2_854e7902,
        64'h74a270e2_744200c7,
        64'h9c63974e_00e58833,
        64'h00379713_47818d5d,
        64'h91011782_65a26602,
        64'h15028fc1_8d450109,
        64'h179b0105_151b9a3f,
        64'he0ef84aa_9a9fe0ef,
        64'h892a9aff_e0ef842a,
        64'h9b5fe0ef_89aaec4e,
        64'hf04af426_f822fc06,
        64'he032e42e_7139b7f1,
        64'h00e83023_8f490008,
        64'h3703e314_8ec90785,
        64'h6314b8df_f06f6121,
        64'h863e69e2_854e7902,
        64'h74a270e2_744200c7,
        64'h9c63974e_00e58833,
        64'h00379713_47818d5d,
        64'h91011782_65a26602,
        64'h15028fc1_8d450109,
        64'h179b0105_151ba1bf,
        64'he0ef84aa_a21fe0ef,
        64'h892aa27f_e0ef842a,
        64'ha2dfe0ef_89aaec4e,
        64'hf04af426_f822fc06,
        64'he032e42e_7139b7d1,
        64'h00e83023_02a75733,
        64'h00083703_e31402a6,
        64'hd6b30785_63144505,
        64'he111c0df_f06f6121,
        64'h863e69e2_854e7902,
        64'h74a270e2_744200c7,
        64'h9c63974e_00e58833,
        64'h00379713_47818d5d,
        64'h91011782_65a26602,
        64'h15028fc1_8d450109,
        64'h179b0105_151ba9bf,
        64'he0ef84aa_aa1fe0ef,
        64'h892aaa7f_e0ef842a,
        64'haadfe0ef_89aaec4e,
        64'hf04af426_f822fc06,
        64'he032e42e_7139b7e1,
        64'h00e83023_02a70733,
        64'h00083703_e31402a6,
        64'h86b30785_6314c89f,
        64'hf06f6121_863e69e2,
        64'h854e7902_74a270e2,
        64'h744200c7_9c63974e,
        64'h00e58833_00379713,
        64'h47818d5d_91011782,
        64'h65a26602_15028fc1,
        64'h8d450109_179b0105,
        64'h151bb17f_e0ef84aa,
        64'hb1dfe0ef_892ab23f,
        64'he0ef842a_b29fe0ef,
        64'h89aaec4e_f04af426,
        64'hf822fc06_e032e42e,
        64'h7139b7f1_00e83023,
        64'h8f090008_3703e314,
        64'h8e890785_6314d01f,
        64'hf06f6121_863e69e2,
        64'h854e7902_74a270e2,
        64'h744200c7_9c63974e,
        64'h00e58833_00379713,
        64'h47818d5d_91011782,
        64'h65a26602_15028fc1,
        64'h8d450109_179b0105,
        64'h151bb8ff_e0ef84aa,
        64'hb95fe0ef_892ab9bf,
        64'he0ef842a_ba1fe0ef,
        64'h89aaec4e_f04af426,
        64'hf822fc06_e032e42e,
        64'h7139b7f1_00e83023,
        64'h8f290008_3703e314,
        64'h8ea90785_6314d79f,
        64'hf06f6121_863e69e2,
        64'h854e7902_74a270e2,
        64'h744200c7_9c63974e,
        64'h00e58833_00379713,
        64'h47818d5d_91011782,
        64'h65a26602_15028fc1,
        64'h8d450109_179b0105,
        64'h151bc07f_e0ef84aa,
        64'hc0dfe0ef_892ac13f,
        64'he0ef842a_c19fe0ef,
        64'h89aaec4e_f04af426,
        64'hf822fc06_e032e42e,
        64'h7139b7ad_0485b0ff,
        64'hf0ef0007_c50397e2,
        64'h0039f793_0985b1ff,
        64'hf0ef4521_ef8100ad,
        64'hb02300ac_b0238d41,
        64'h91011402_150201a4,
        64'h643300a9_6533010d,
        64'h1d1b0105_151b0344,
        64'hf7b3c6ff_e0ef892a,
        64'hc75fe0ef_8d2ac7bf,
        64'he0ef842a_c81fe0ef,
        64'he33ff06f_61657ae2,
        64'h85567b42_64e685da,
        64'h86266da2_6d426ce2,
        64'h7c027ba2_6a0669a6,
        64'h694670a6_7406962f,
        64'hd0eff025_05130000,
        64'h35170374_9b6300fb,
        64'h0cb300fa_8db30034,
        64'h9793252c_0c130000,
        64'h3c179c4a_0a134981,
        64'hbb1ff0ef_44818bb2,
        64'h8b2ee46e_e86aec66,
        64'he8caf0a2_f486f062,
        64'hf45ef85a_e4ceeca6,
        64'h02000513_8aaa6a05,
        64'hfc56e0d2_7159bfa5,
        64'h07a10585_80826125,
        64'h6ca26c42_6be27b02,
        64'h7aa27a42_79e26906,
        64'h64a66446_60e6557d,
        64'h9dcfd0ef_f3450513,
        64'h00003517_9e8fd0ef,
        64'hf0850513_00003517,
        64'h058e02e6_0d6340e9,
        64'h87330035_9713c689,
        64'h873e8a85_63900085,
        64'h86b3bf5d_07a10485,
        64'h6398e398_40e98733,
        64'h00349713_c689873e,
        64'h8a850084_86b3a889,
        64'h4501a2ef_d0effa65,
        64'h05130000_3517fd54,
        64'h17e30405_02b49b63,
        64'h458187ca_a48fd0ef,
        64'h856285e6_a50fd0ef,
        64'h85520364_98634481,
        64'h87caa5ef_d0ef855e,
        64'h85e60004_0c9ba6af,
        64'hd0ef8552_4ac1f7ec,
        64'h0c130000_3c17fff9,
        64'h4993f7ab_8b930000,
        64'h3b97f72a_0a130000,
        64'h3a17a8ef_d0ef4401,
        64'h8b2ee466_e4a6ec86,
        64'he862ec5e_f05af456,
        64'hf852fc4e_e8a2f865,
        64'h05130000_3517892a,
        64'he0ca711d_bf5d0785,
        64'ha001abef_d0eff865,
        64'h05130000_351785a2,
        64'h8626acef_d0eff6e5,
        64'h05130000_35176090,
        64'h600c02e8_03636098,
        64'h00043803_80826105,
        64'h450164a2_644260e2,
        64'h00c79863_00d50433,
        64'h00d584b3_00379693,
        64'h4781e426_e822ec06,
        64'h1101c2df_f06f8082,
        64'h45018082_45018082,
        64'h80828082_80824509,
        64'h80824509_80824509,
        64'hbff92605_20040413,
        64'h6622edbf_c0efe432,
        64'h852285b2_80826145,
        64'h450164e2_740270a2,
        64'h00961863_00c684bb,
        64'h842ef406_ec26f022,
        64'h71798082_45058082,
        64'h45058082_45058082,
        64'h01418d7d_640260a2,
        64'h95224080_07b3f57f,
        64'hf0efe406_952e842a,
        64'he0221141_a001d2df,
        64'hf0ef4505_b90fd0ef,
        64'he406ffa5_05130000,
        64'h351785aa_862e86b2,
        64'h87361141_808202f5,
        64'h553347a9_b0002573,
        64'h80824501_80824501,
        64'h80820141_450160a2,
        64'hf89fc0ef_20000537,
        64'hbccfd0ef_e40600e5,
        64'h05130000_35171141,
        64'h80828082_61056442,
        64'h60e28522_9e8ff0ef,
        64'h45816622_c509842a,
        64'hfd1ff0ef_e4328532,
        64'hec06e822_110102b5,
        64'h06338082_953e055e,
        64'h10d00513_e3089536,
        64'h00178693_00756513,
        64'h157d631c_89c70713,
        64'h00004717_80824501,
        64'h80822405_0513000f,
        64'h4537a001_ddbff0ef,
        64'he4062501_11419002,
        64'h00000023_e8dff0ef,
        64'hc4cfd0ef_84450513,
        64'h00003517_bdddc5af,
        64'hd0ef0725_05130000,
        64'h3517c981_c62e0005,
        64'h059b962f_90ef0184,
        64'h951385a2_c78fd0ef,
        64'h07850513_00003517,
        64'hc84fd0ef_03c50513,
        64'h00003517_85a20184,
        64'h961386a2_0bf00493,
        64'hbf1d03a5_05130000,
        64'h3517c511_2501dabf,
        64'ha0ef4501_d4458593,
        64'h00003597_4605bf91,
        64'h02850513_00003517,
        64'hbfb904a5_05130000,
        64'h3517c919_2501c96f,
        64'hb0ef5402_0808f3f9,
        64'h9cbd47b2_286010ef,
        64'h854edbff_f0ef0004,
        64'h45039452_dc9ff0ef,
        64'h880d4521_0004099b,
        64'h00c4d41b_e5052501,
        64'hfedfa0ef_080895ca,
        64'h66050074_91810204,
        64'h959314aa_0a130000,
        64'h3a170962_0bf00913,
        64'he12d4481_2501e85f,
        64'ha0ef0808_08c58593,
        64'h00003597_4605d3af,
        64'hd0ef07a5_05130000,
        64'h35178082_27010113,
        64'h24013a03_24813983,
        64'h25013903_25813483,
        64'h26013403_26813083,
        64'hd64fd0ef_08450513,
        64'h00003517_c5152501,
        64'he75fa0ef_25413023,
        64'h25313423_25213823,
        64'h24913c23_26813023,
        64'h26113423_a1450513,
        64'h00004517_e2c58593,
        64'h00003597_4605d901,
        64'h01138302_037eab65,
        64'h85930000_25974305,
        64'hf1402573_0ff0000f,
        64'h0000100f_80826105,
        64'h60e2e9ff_f0ef0091,
        64'h4503ea7f_f0ef0081,
        64'h4503f13f_f0efec06,
        64'h002c1101_80826145,
        64'h694264e2_740270a2,
        64'hfe9410e3_ec9ff0ef,
        64'h00914503_ed1ff0ef,
        64'h34610081_4503f3ff,
        64'hf0ef0ff5_7513002c,
        64'h00895533_54e10380,
        64'h0413892a_f406e84a,
        64'hec26f022_71798082,
        64'h61456942_64e27402,
        64'h70a2fe94_10e3f0bf,
        64'hf0ef0091_4503f13f,
        64'hf0ef3461_00814503,
        64'hf81ff0ef_0ff57513,
        64'h002c0089_553b54e1,
        64'h4461892a_f406e84a,
        64'hec26f022_71798082,
        64'h61056442_60e2f43f,
        64'hf0ef0091_4503f4bf,
        64'hf0ef0081_4503fb7f,
        64'hf0ef0ff4_7513002c,
        64'hf5dff0ef_00914503,
        64'hf65ff0ef_00814503,
        64'hfd1ff0ef_ec068121,
        64'h842a002c_e8221101,
        64'h808200f5_802300e5,
        64'h80a30007_c7830007,
        64'h470397aa_973e8111,
        64'h00f57713_b9478793,
        64'h00002797_b7f50405,
        64'hfa5ff0ef_80820141,
        64'h640260a2_e5090004,
        64'h4503842a_e406e022,
        64'h11418082_00e78823,
        64'h02000713_00e78423,
        64'hfc700713_00e78623,
        64'h470d0007_822300e7,
        64'h8023476d_00e78623,
        64'hf8000713_00078223,
        64'h100007b7_808200a7,
        64'h0023dfe5_0207f793,
        64'h01474783_10000737,
        64'h80820205_75130147,
        64'hc5031000_07b78082,
        64'h00054503_808200b5,
        64'h00238082_61056902,
        64'h64a26442_60e2f47d,
        64'hfa1ff0ef_41240433,
        64'h854a8926_0084f363,
        64'h89226804_8493842a,
        64'he04aec06_e8220098,
        64'h94b7e426_11018082,
        64'h61056902_64a26442,
        64'h60e2fe85_6ee3f45f,
        64'hf0ef0405_944a0285,
        64'h54332404_0413000f,
        64'h443702a4_85333700,
        64'h00ef892a_f63ff0ef,
        64'h84aae04a_e426e822,
        64'hec061101_808202a7,
        64'hd5330141_91011502,
        64'h640260a2_02f407b3,
        64'h24078793_000f47b7,
        64'h3a2000ef_842af95f,
        64'hf0efe022_e4061141,
        64'h80826105_64a28d05,
        64'h02a7d533_644260e2,
        64'h91011502_02f407b3,
        64'h3e800793_3ce000ef,
        64'h842afc1f_f0ef84aa,
        64'he426e822_ec061101,
        64'h80824501_80820141,
        64'h8d5d9101_17821502,
        64'h60a21007_e78310a7,
        64'ha22310e1_a0232705,
        64'h1001a703_00e57763,
        64'h878e1041_e7034920,
        64'h00efe406_11418082,
        64'hcf5ff06f_aac58593,
        64'h00004597_4611cb81,
        64'hcc47d783_00004797,
        64'h80822401_01132201,
        64'h39032281_34832301,
        64'h34032381_3083f63f,
        64'hf0ef8522_002ced4f,
        64'hf0efe802_c44a0828,
        64'h20400613_85a6e92f,
        64'hf0ef2211_3c230028,
        64'h21800613_45818932,
        64'h84ae842a_23213023,
        64'h22913423_22813823,
        64'hdc010113_ebfff06f,
        64'h614505c1_70a24190,
        64'h7402d8df_f06f6145,
        64'h70a265a2_74028522,
        64'h8d5fd0ef_e42e3be5,
        64'h05130000_3517842a,
        64'h8e5fd06f_61453e65,
        64'h05130000_351770a2,
        64'h740202e7_8a63470d,
        64'h00e78e63_01e15783,
        64'h00f10f23_0115c783,
        64'h00f10fa3_47090105,
        64'hc783f022_f4067179,
        64'h80826105_690264a2,
        64'h644260e2_d61ff06f,
        64'h61056902_64a260e2,
        64'h6442937f_d0ef4065,
        64'h05130000_35170087,
        64'hcf63278d_439cdae7,
        64'h87930000_4797daf7,
        64'h1d230000_47172785,
        64'h0007d783_dc878793,
        64'h00004797_240000ef,
        64'h02000513_d35ff0ef,
        64'h4515dde5_d5830000,
        64'h45972560_00ef4535,
        64'he2dff0ef_854abe65,
        64'h85930000_4597bea7,
        64'h98230000_47974611,
        64'hd23ff0ef_e0855503,
        64'h00004517_c0a79223,
        64'h00004797_d37ff0ef,
        64'h4511dc3f_f0ef0044,
        64'h8513ffc4_059b06a7,
        64'h9a632501_0024d783,
        64'hd53ff0ef_e3855503,
        64'h00004517_08a79563,
        64'h25010004_d783d69f,
        64'hf0ef84ae_450d892a,
        64'h08c7df63_8432478d,
        64'he04ae426_ec06e822,
        64'h1101b799_e6879423,
        64'h00004797_eb1ff0ef,
        64'h854ec6a5_85930000,
        64'h45974611_c6a79b23,
        64'h00004797_da7ff0ef,
        64'h4501c8a7_91230000,
        64'h4797db5f_f0efeaf7,
        64'h33230000_4717eaf7,
        64'h33230000_47174511,
        64'h01f41793_4405a4bf,
        64'hd0ef4fa5_05130000,
        64'h3517858a_4390ebe7,
        64'h87930000_4797e22f,
        64'hf0ef850a_85a2e2af,
        64'hf0ef850a_51458593,
        64'h00003597_00f70963,
        64'h02f00793_01294703,
        64'he1aff0ef_850a31e5,
        64'h85930000_3597893f,
        64'hf0ef850a_45811000,
        64'h0613b755_f0f72223,
        64'h00004717_20000793,
        64'h80826155_69b26952,
        64'h64f27412_70b2abbf,
        64'hd0ef5425_05130000,
        64'h351700a4_05b3f54f,
        64'hf0ef3625_05130000,
        64'h3517842a_f62ff0ef,
        64'h852204a7_f2630ff0,
        64'h07939526_f72ff0ef,
        64'h38050513_00003517,
        64'h84aaf80f_f0ef8522,
        64'hf6a7a023_00004797,
        64'h04e7ee63_1ff00793,
        64'hfff5071b_eabff0ef,
        64'h95260505_fa2ff0ef,
        64'h852600a4_04b30505,
        64'hfaeff0ef_892eea4a,
        64'hee26f606_852289aa,
        64'he64e0125_8413f222,
        64'h71698082_45018082,
        64'h01416402_60a2557d,
        64'h00850363_8c0fa0ef,
        64'h8432e406_e0221141,
        64'h83026105_250106e5,
        64'h85930000_25976902,
        64'h834a64a2_60e26442,
        64'hf1402573_0ff0000f,
        64'h0000100f_b81fd0ef,
        64'h5f050513_00003517,
        64'h862286aa_608ce77f,
        64'hc0ef85a2_6088b9bf,
        64'hd0ef85a2_4124043b,
        64'hec065fa5_05130000,
        64'h35170004_b9036380,
        64'he04ae822_02448493,
        64'h00004497_03478793,
        64'h00004797_e4261101,
        64'h80826105_64a26442,
        64'he00c95a6_60e2600c,
        64'ha2fff0ef_ec066008,
        64'h85aa84ae_862ee426,
        64'h06040413_00004417,
        64'he8221101_808206f7,
        64'h37230000_471706f7,
        64'h37230000_471707fe,
        64'h47854e60_006f0305,
        64'h05130141_60a26402,
        64'h02a4753b_4529fe7f,
        64'hf0ef357d_02b455bb,
        64'h45a900b7_f86347a5,
        64'h00a04563_842ee406,
        64'he0221141_bff90505,
        64'hfd07879b_9fb902f5,
        64'h87bb00d6_67630ff6,
        64'hf693fd07_069b8082,
        64'h853ee319_00054703,
        64'h45a94625_47818082,
        64'h014100e1_550300a1,
        64'h07238121_00a107a3,
        64'h1141fa5f_f06f4581,
        64'hd7dff06f_01410505,
        64'h45814629_60a26402,
        64'hf77d8b11_00074703,
        64'h973e0005_4703fea4,
        64'h7ae3157d_80820141,
        64'h557d6402_60a2e719,
        64'h8b110007_4703973e,
        64'hfff58513_c3c78793,
        64'h00002797_fff5c703,
        64'h00a405b3_95bff0ef,
        64'he589842a_e406e022,
        64'h1141bfd5_0789bff1,
        64'h052a052a_b7e9e01c,
        64'h078d00e6_98630420,
        64'h07130027_c683fce6,
        64'h9fe3052a_06900713,
        64'h0017c683_fed716e3,
        64'h06b00693_02d70763,
        64'h04d00693_80820141,
        64'h640260a2_02d70e63,
        64'h04700693_00e6ea63,
        64'h02d70463_0007c703,
        64'h04b00693_601cf87f,
        64'hf0ef842e_e406e022,
        64'h1141b7e1_e008b7cd,
        64'hfc97879b_0ff7f793,
        64'hfe07079b_c6098a09,
        64'hb7d196be_050502d5,
        64'h86b3feb7_f4e3fd07,
        64'h879b0008_8b630046,
        64'h78938082_61058536,
        64'h644260e2_ec050008,
        64'h98630446_78930006,
        64'h460300f8_06330007,
        64'h079b0005_4703d168,
        64'h08130000_28174681,
        64'h00c16583_e0fff0ef,
        64'hc632ec06_006c842e,
        64'he8221101_bfd50789,
        64'hbff1052a_052ab7e9,
        64'he01c078d_00e69863,
        64'h04200713_0027c683,
        64'hfce69fe3_052a0690,
        64'h07130017_c683fed7,
        64'h16e306b0_069302d7,
        64'h076304d0_06938082,
        64'h01416402_60a202d7,
        64'h0e630470_069300e6,
        64'hea6302d7_04630007,
        64'hc70304b0_0693601c,
        64'hf0dff0ef_842ee406,
        64'he0221141_80820141,
        64'h40a00533_60a2f23f,
        64'hf0efe406_05051141,
        64'hf2dff06f_00e68463,
        64'h02d00713_00054683,
        64'hb7e94501_e088fcf7,
        64'h18e347a9_fd279be3,
        64'h07858f81_cb010007,
        64'hc703fe87_82e367e2,
        64'hf5dff0ef_8522082c,
        64'h892a862e_80826121,
        64'h790274a2_744270e2,
        64'h5529e901_65a2b0df,
        64'hf0ef84b2_842ae42e,
        64'h00063023_f04afc06,
        64'hf426f822_7139b7e1,
        64'he008b7cd_fc97879b,
        64'h0ff7f793_fe07079b,
        64'hc6098a09_b7d196be,
        64'h050502d5_86b3feb7,
        64'hf4e3fd07_879b0008,
        64'h8b630046_78938082,
        64'h61058536_644260e2,
        64'hec050008_98630446,
        64'h78930006_460300f8,
        64'h06330007_079b0005,
        64'h4703e6a8_08130000,
        64'h28174681_00c16583,
        64'hf63ff0ef_c632ec06,
        64'h006c842e_e8221101,
        64'hbf6d47a9_bf7d47a1,
        64'h80820509_00e79363,
        64'h07800713_0ff7f793,
        64'h0207879b_c7098b05,
        64'h00074703_973eeae7,
        64'h07130000_27170015,
        64'h478302f7_16630300,
        64'h07930005_470302f7,
        64'h1c6347c1_4198c19c,
        64'h47c1c3b1_0447f793,
        64'h0007c783_97ba0025,
        64'h470304d7_1b630780,
        64'h06930ff7_77130207,
        64'h071bc689_8a850006,
        64'hc68300e7_86b3efe7,
        64'h87930000_27970015,
        64'h470308f7_11630300,
        64'h07930005_4703e7a9,
        64'h419cb7f1_377d87aa,
        64'hbfa5fef5_1be30785,
        64'hf8b712e3_0007c703,
        64'h00d80a63_00878513,
        64'h0007b803_bfcd367d,
        64'h0785f8b7_1fe30007,
        64'hc703d24d_8a1deb11,
        64'h87aa2701_8edd0036,
        64'h57130207_96938fd9,
        64'h01071793_00b7e733,
        64'h00859793_8e1d953e,
        64'h93810207_1793faf5,
        64'h078536fd_fcb81ce3,
        64'h0007c803_87aa0007,
        64'h069b40e7_873b47a1,
        64'hc31d0075_7713b7f5,
        64'h367d0785_feb71ce3,
        64'h0007c703_8082853e,
        64'h4781e601_87aa2601,
        64'h00c7ef63_0ff5f593,
        64'h47c1b7ed_853efeb7,
        64'h0be30015_07930005,
        64'h47038082_450100c5,
        64'h14630ff5_f593962a,
        64'hbfe90405_d175f8bf,
        64'hf0ef397d_852285ce,
        64'h86268082_614569a2,
        64'h694264e2_740270a2,
        64'h85224401_00995b63,
        64'h0005091b_d13ff0ef,
        64'h8522c889_0005049b,
        64'hd1fff0ef_89aee84a,
        64'hf406e44e_ec26852e,
        64'h842af022_7179bfc5,
        64'h0505feb7_8de30005,
        64'h47838082_00c51363,
        64'h962ab7dd_05850505,
        64'hfbed9f99_0005c703,
        64'h00054783_8082853e,
        64'h478100c5_1563962a,
        64'hb7fd00f6_802316fd,
        64'h0005c783_15fdd7e5,
        64'h00e587b3_40b60733,
        64'h00c506b3_95b28082,
        64'h01416402_60a28522,
        64'hf57ff0ef_00a5e963,
        64'h842ae406_e0221141,
        64'h80826145_64e26942,
        64'h85267402_70a20004,
        64'h0023f79f_f0ef944a,
        64'h864a8522_fff60913,
        64'h00c56463_6582892a,
        64'hce1184aa_6622dcdf,
        64'hf0efe02e_e84af406,
        64'he432ec26_852e842a,
        64'hf0227179_bf65fee7,
        64'h8fa30785_fff5c703,
        64'h0585bfe1_469d00c5,
        64'h08b387aa_872ebfc1,
        64'h00e507b3_963e95ba,
        64'h070e02f7_07b357e1,
        64'h00365713_ff06e8e3,
        64'h40f88833_ff07bc23,
        64'h07a1ff87_38030721,
        64'h808202c7_9e63963e,
        64'h87aacb9d_8b9d00a5,
        64'he7b300b5_0a63bf6d,
        64'hfeb78fa3_0785bfe1,
        64'hfef73c23_0721bfd1,
        64'h0ff5f693_4725bfc1,
        64'h963a97aa_078e02e7,
        64'h87335761_00365793,
        64'h0106ef63_40e88833,
        64'h469d00c5_08b3872a,
        64'hff6d377d_8fd507a2,
        64'h808204c7_9063963e,
        64'h87aacb9d_00757793,
        64'h80824501_b7e50789,
        64'h00d780a3_00e78023,
        64'h8082e311_0017c703,
        64'hce810007_c68387aa,
        64'hcf990005_4783c11d,
        64'h80826105_64a28526,
        64'h644260e2_e0080505,
        64'h00050023_c501f73f,
        64'hf0ef8526_842ac891,
        64'he822ec06_6104e426,
        64'h1101bfd9_4aa7b623,
        64'h00004797_05050005,
        64'h0023c781_00054783,
        64'hc519f9ff_f0ef8522,
        64'h85a68082_610564a2,
        64'h644260e2_85224401,
        64'h4c07bc23_00004797,
        64'hef810004_4783942a,
        64'hf9dff0ef_85a68522,
        64'hcc116380_4f478793,
        64'h00004797_e519842a,
        64'h84aeec06_e426e822,
        64'h1101bfd5_87aeb7e5,
        64'h0505fafd_0007c683,
        64'h0785fee6_8fe38082,
        64'h4501eb19_00054703,
        64'hbff90785_bfd5872e,
        64'h8082fe08_1be30007,
        64'h48030705_00c80a63,
        64'h8082ea11_40d78533,
        64'h0007c603_87aa86aa,
        64'hbfcd872e_b7d50785,
        64'hfe081be3_00074803,
        64'h0705fed8_0fe38082,
        64'hea9940c7_85330007,
        64'hc68387aa_862ab7fd,
        64'h07858082_40a78533,
        64'he7010007_c70300b7,
        64'h856387aa_95aa8082,
        64'h61056442_60e24501,
        64'hfe857be3_157d00b7,
        64'h86630005_47830ff5,
        64'hf5939522_65a2fe5f,
        64'hf0efec06_842ae42e,
        64'he8221101_bfcd0785,
        64'h808240a7_8533e701,
        64'h0007c703_87aabfcd,
        64'h0505dffd_808200b7,
        64'h93630005_47830ff5,
        64'hf5938082_4501bfcd,
        64'h0505c399_808200b7,
        64'h93630005_47830ff5,
        64'hf5938082_853eff79,
        64'h0505e399_4187d79b,
        64'h0187979b_40f707bb,
        64'hfff5c783_00054703,
        64'h0585a839_478100c5,
        64'h9463962e_8082853e,
        64'hf37d0505_e3994187,
        64'hd79b0187_979b40f7,
        64'h07bbfff5_c7830005,
        64'h47030585_b7cd87ba,
        64'h80820007_80a300c7,
        64'h15638082_e291fed7,
        64'h0fa30017_8713fff5,
        64'hc6830585_963efb7d,
        64'h00178693_0007c703,
        64'h87b68082_e21987aa,
        64'hb7d587b6_8082fb75,
        64'hfee78fa3_0785fff5,
        64'hc7030585_eb090017,
        64'h86930007_c70387aa,
        64'h8082fb65_fee78fa3,
        64'h0785fff5_c7030585,
        64'h00c78963_87aa962a,
        64'h8082fb75_fee78fa3,
        64'h0785fff5_c7030585,
        64'h87aa8082_01416402,
        64'h60a28d41_15029001,
        64'hfd1ff0ef_14020005,
        64'h041bfdbf_f0efe022,
        64'he4061141_80820141,
        64'h25016402_60a28d41,
        64'h0105151b_fe9ff0ef,
        64'h842afeff_f0efe022,
        64'he4061141_fc3ff06f,
        64'h6f850513_00004517,
        64'h80822501_8d5d00f7,
        64'h17bb40f0_07b300f7,
        64'h553b93ed_836d8f3d,
        64'h0127d713_e1189736,
        64'h00176713_02d786b3,
        64'h65186294_611c4966,
        64'h86930000_46971180,
        64'h106f8082_61056902,
        64'h64a26442_60e28522,
        64'he99ff0ef_10f40023,
        64'h0247c783_85220ea4,
        64'h2e23681c_18f43423,
        64'h20a78793_00001797,
        64'h18f43023_21a78793,
        64'h00001797_16f43c23,
        64'h91c78793_fffff797,
        64'he65ff0ef_04052823,
        64'h03253023_e90410f5,
        64'h02a34785_0ef52c23,
        64'h4799c57c_57fdcd21,
        64'h842a15c0_10ef4505,
        64'h1c000593_84aa892e,
        64'hc7ad639c_c7bd651c,
        64'hcbad511c_cbbd4d5c,
        64'hcfad4401_4d1cc141,
        64'h4401e04a_e426ec06,
        64'he8221101_b7716000,
        64'h286010ef_57450513,
        64'h00003517_01a98863,
        64'hda4fe0ef_856685e2,
        64'h00978e63_601cdb2f,
        64'he0ef855e_85ca0009,
        64'h0663dbef_e0ef638c,
        64'h855a0fc4_2603681c,
        64'h89560007_c3638952,
        64'h4c1cc791_4901541c,
        64'hddcfe06f_61251165,
        64'h05130000_45176d02,
        64'h6ca26c42_6be27b02,
        64'h7aa27a42_79e26906,
        64'h64a660e6_64460294,
        64'h15634d29_5ecc8c93,
        64'h00003c97_00050c1b,
        64'h058b8b93_00004b97,
        64'h058b0b13_00004b17,
        64'h050a8a93_00004a97,
        64'h060a0a13_00004a17,
        64'h89aae0ca_ec86e06a,
        64'he466e862_ec5ef05a,
        64'hf456f852_fc4e6080,
        64'he8a28824_84930000,
        64'h5497e4a6_711d8082,
        64'he308e518_e11ce788,
        64'h679889a7_87930000,
        64'h5797e508_80827207,
        64'hab230000_4797e79c,
        64'he39c8b27_87930000,
        64'h5797b7d5_6000a9cf,
        64'hf0ef8522_c78119a4,
        64'h47838082_610564a2,
        64'h644260e2_00941763,
        64'h84beec06_e4266380,
        64'he8228e27_87930000,
        64'h57971101_80824388,
        64'h78078793_00004797,
        64'h80820f85_05138082,
        64'hc3980015_071b4388,
        64'h79878793_00004797,
        64'hbfd55535_80826105,
        64'h64a26442_60e2e080,
        64'h0f840413_e501cf0f,
        64'hf0ef842a_cd09f7df,
        64'hf0ef84ae_e822ec06,
        64'he4261101_bfcdf840,
        64'h0513bfe5_45018082,
        64'h610560e2_5535eb3f,
        64'he06f6105_60e200f7,
        64'h0c630ff0_07930815,
        64'h470302b7_006365a2,
        64'h10354703_c105fbdf,
        64'hf0efe42e_ec061101,
        64'h41488082_853ebfd1,
        64'h87b600a6_04630fc7,
        64'ha6038082_0141853e,
        64'h478160a2_f60fe0ef,
        64'he4061725_05130000,
        64'h451785aa_114102e7,
        64'h90636394_631c9ae7,
        64'h07130000_57178082,
        64'h45018082_01414501,
        64'h640260a2_0dc000ef,
        64'h13e000ef_02c00513,
        64'hfc5ff0ef_85220005,
        64'h5563aeef_e0ef8522,
        64'h12a000ef_9ef72023,
        64'h00005717_842ae406,
        64'he0224785_1141ef9d,
        64'h439c9f67_87930000,
        64'h57978082_18b50d23,
        64'h8082557d_8082557d,
        64'h80824501_c56ce54f,
        64'hf06ffa10_0413f0ef,
        64'hf06f2006_061b4001,
        64'h0637f0a6_09634505,
        64'hf0c54363_8ca602e3,
        64'h45098a3d_01a6d61b,
        64'hf2c51a63_40000637,
        64'h06bba423_06eba223,
        64'h06fba023_04dbae23,
        64'h018ba503_45e64756,
        64'h47c646b6_ea051163,
        64'h842a93bf_e0efc4be,
        64'h855e0107_979b008c,
        64'h460107cb_d783c2be,
        64'h479d04f1_102347a5,
        64'h06fb9e23_04e15783,
        64'h0007d663_018ba783,
        64'hec051b63_842a96ff,
        64'he0efc2be_47d5855e,
        64'hc4be0107_979b008c,
        64'h460107cb_d78304f1,
        64'h1023478d_6da000ef,
        64'h06cb8513_00ec4641,
        64'hbf6d1187_2583974e,
        64'h83790207_9713fcfc,
        64'h65e34581_b7c9f521,
        64'hd31fe0ef_855e4585,
        64'h0b700613_0ff6f693,
        64'hbb91fd31_9fdfe0ef,
        64'h855ecb0f_f0ef855e,
        64'h460118fb_ae2308bb,
        64'ha2230017_b79317ed,
        64'h088ba583_ef8d1afb,
        64'ha823409c_e79d0046,
        64'hf7930089_2683f941,
        64'h808ff0ef_855e408c,
        64'h933fe0ef_855e02eb,
        64'haa230017_b71341b7,
        64'h87b301a7_86634711,
        64'h00d78963_47214000,
        64'h06b70009_2783bb6d,
        64'h925fe0ef_1c450513,
        64'h00004517_f7649fe3,
        64'h04a1fb99_11e30931,
        64'h973fe0ef_855e035b,
        64'haa2308fb_a223180b,
        64'hae231a0b_a823088b,
        64'ha783ddbf_e0ef855e,
        64'h45850b70_06134681,
        64'hc131debf_e0ef855e,
        64'h0fb6f693_45850b70,
        64'h06130089_4683c3a1,
        64'h8ff900fa_77b30009,
        64'h270340dc_04f71863,
        64'h0017b793_17ed0049,
        64'h4703409c_10000db7,
        64'h20000d37_da490913,
        64'h00003917_cbb52781,
        64'h00fa77b3_00fa97bb,
        64'h409cdf6c_8c930000,
        64'h3c974c2d_dc4b0b13,
        64'h00003b17_4a85db4f,
        64'hf0efdb24_84930000,
        64'h349700fa_7a33855e,
        64'h4601088b_a583044b,
        64'ha783040b_aa0304fb,
        64'ha02300c7_e793040b,
        64'ha783c799_8b8504eb,
        64'ha0230107_6713040b,
        64'ha70304eb_a0230217,
        64'h071bc689_00c7f693,
        64'hce910027_f6931adb,
        64'ha42303f7_f6930c46,
        64'hc78304fb_a0230017,
        64'h079b7000_0737bb95,
        64'h2f050513_00004517,
        64'he691ecf7_6ce31a0b,
        64'hb6834004_07b704fb,
        64'ha0232785_100007b7,
        64'hb8d102fb_a4234785,
        64'h740010ef_8526a3ff,
        64'he0ef8a3d_8abd0146,
        64'h561b0106_569b0624,
        64'h85133725_85930000,
        64'h4597074b_a603a5ff,
        64'he0ef04d4_85133765,
        64'h85930000_45972681,
        64'h0ff77713_0ff87813,
        64'h0ff7f793_0188569b,
        64'h0108571b_0088579b,
        64'h06cbc603_077bc883,
        64'h070ba803_a95fe0ef,
        64'hfef53623_02450513,
        64'h39858593_00004597,
        64'h84aa06fb_c603074b,
        64'hd68307ab_d70302c7,
        64'hd7b3ed10_92010a8b,
        64'hb783d11c_9fb90712,
        64'h00e03733_8f750207,
        64'h161376c1_9fb5068e,
        64'h00d036b3_8ef9f006,
        64'h8693ff01_06b79fb5,
        64'h068a00d0_36b38ef9,
        64'h0f068693_f0f0f6b7,
        64'h9fb500f0_37b30686,
        64'h00d036b3_27818ef9,
        64'h8ff9ccc6_8693aaa7,
        64'h8793cccc_d6b7aaaa,
        64'hb7b708cb_a7030005,
        64'h06230005_15234840,
        64'h00ef855e_08fba823,
        64'h08fba623_20000793,
        64'hc79919cb_a7831afb,
        64'haa231b0b_a7830adb,
        64'ha2230afb_a02302d6,
        64'h06bb02f7_57bb8a8d,
        64'h0106d69b_02e6073b,
        64'h3e800613_c305c38d,
        64'h03f77713_27810126,
        64'hd71b8fd1_0186d61b,
        64'h8ff917fd_67c100cc,
        64'ha68308fb_ae230087,
        64'h171b1487_a78397b6,
        64'h078af026_86930000,
        64'h369704d6_1c638003,
        64'h06b7018b_a60300f6,
        64'hf8638bbd_00c7579b,
        64'h46a5008c_a703fdb5,
        64'h9ee3fefd_ae238fd9,
        64'h8ff58f51_0087d79b,
        64'h8e690087_961b8f51,
        64'h0187971b_0187d61b,
        64'h0d91000d_a783f006,
        64'h869300ff_0537040d,
        64'h859366c1_b5451187,
        64'h2583974e_83790207,
        64'h9713eaf7_68e34581,
        64'h472db35d_04fba023,
        64'h00876793_da06d9e3,
        64'h040ba703_02e79693,
        64'h8fd18ff5_0087d79b,
        64'h0087961b_f0068693,
        64'h66c144dc_fbe18b85,
        64'h83a54cdc_d0051ce3,
        64'hd61fe0ef_dc3ef84a,
        64'hf426c556_855e010c,
        64'h04000793_1030c33e,
        64'h47d508f1_10234799,
        64'h020a0863_3a7d0905,
        64'h3ac54a15_98811902,
        64'h01000ab7_0ff10493,
        64'h4905bbc5_80030737,
        64'hde075ee3_03079713,
        64'h00ebac23_80020737,
        64'hb519a007_071b8001,
        64'h1737b61d_df400413,
        64'hcbdfe0ef_55c50513,
        64'h00004517_e6f49fe3,
        64'h0b078793_00003797,
        64'h04a1eafa_94e347a1,
        64'h0a918c9f_f0ef855e,
        64'h84058593_4601180b,
        64'hae23096b_a2231afb,
        64'ha823017d_85b74785,
        64'hf3ed37fd_670267a2,
        64'h0e050c63_e0dfe0ef,
        64'he03ac93a_e552e16e,
        64'he43e855e_110c0110,
        64'h04000713_4791d502,
        64'hd33a0af1_102347b5,
        64'h6702e915_e35fe0ef,
        64'hd53ee03a_d33a8cee,
        64'h855e110c_0107979b,
        64'h46014755_07cbd783,
        64'h0af11023_03700793,
        64'hfe07fd93_0ff10793,
        64'h947ff0ef_855e4601,
        64'h18fbae23_08bba223,
        64'h0017b793_17ed088b,
        64'ha5831407_9a631afb,
        64'ha823409c_09b79463,
        64'h8bbd010c_4783e941,
        64'he91fe0ef_c93ee552,
        64'he162855e_110c0400,
        64'h07930110_d53e00fd,
        64'he7b317c1_2d818100,
        64'h07b7d33e_47d50af1,
        64'h10234799_4d850ce7,
        64'h9163470d_01a78663,
        64'h409cdfdf_e0ef855e,
        64'h02fbaa23_001cb793,
        64'h40fc8cb3_100007b7,
        64'h00ec8863_47912000,
        64'h073700ec_8d6347a1,
        64'h40000737_0e051c63,
        64'h8daa971f_f0ef855e,
        64'h0015b593_40bc85b3,
        64'h100005b7_00fc8863,
        64'h45912000_07b700fc,
        64'h8d6345a1_400007b7,
        64'h14078163_0197f7b3,
        64'h00f977b3_40dc0007,
        64'hac8397d6_109c840b,
        64'h0b1b4a81_017d8b37,
        64'h16078563_278100f9,
        64'h77b300e7_97bb4785,
        64'h40980a05_fe07fc13,
        64'h83f97913_0ff10793,
        64'h00f97933_23448493,
        64'h00003497_020d1a13,
        64'h044ba783_f0be4d05,
        64'h040ba903_639ce1e7,
        64'h87930000_57971ef7,
        64'h18638001_07b7018b,
        64'ha70304fb_a0238fd9,
        64'h20000737_040ba783,
        64'h00075963_02d79713,
        64'h00ebac23_80010737,
        64'h20d70263_46892127,
        64'h00638b3d_0187d71b,
        64'h04ebac23_8f558f71,
        64'h8ecd0087_571b8de9,
        64'h0087159b_8ecd0187,
        64'h169b0187_559b40d8,
        64'h04fbaa23_27818fd5,
        64'h8ef1f007_06138fd1,
        64'h67410087_569b8e69,
        64'h8fd50087_161b0187,
        64'h179b0187_569b00ff,
        64'h05374098_b5558b1d,
        64'h938100f7_571b1782,
        64'h8fd501e7_569b8ff5,
        64'h0027979b_16f16685,
        64'hb54d08bb_a82300b5,
        64'h15bb89bd_0165d59b,
        64'hbd994003_0637a7a9,
        64'h40020637_bb45842a,
        64'hfe0a16e3_3a7dc131,
        64'h850ff0ef_d05aec56,
        64'he826855e_108c0810,
        64'h4b210a85_4a11d482,
        64'h06f11023_98810209,
        64'h1a930330_07930bf1,
        64'h04934905_d2caed05,
        64'h880ff0ef_d4bed2ca,
        64'h855e0107_979b108c,
        64'h460107cb_d78306f1,
        64'h10230370_079304fb,
        64'ha0232789_100007b7,
        64'h54075a63_018ba703,
        64'he0051fe3_842affbf,
        64'he0ef855e_00b54583,
        64'h0f7000ef_855ee205,
        64'h1ae3842a_c9aff0ef,
        64'h855e08fb_80a357fd,
        64'h08fbaa23_4785e405,
        64'h16e3842a_8e4ff0ef,
        64'hc4bec2ca_855e008c,
        64'h0107979b_46014955,
        64'h07cbd783_04f11023,
        64'h479d902f_f0efc282,
        64'hc4be04e1_1023855e,
        64'h008c4601_0107979b,
        64'h471100e7_8e63577d,
        64'h04cba783_c21508fb,
        64'ha82300e7_f4632000,
        64'h0793090b_a70308fb,
        64'ha6230107_d4632000,
        64'h07930afb_b8230e0b,
        64'hb0230c0b_bc230c0b,
        64'hb8230c0b_b4230c0b,
        64'hb0230a0b_bc230307,
        64'h87b300e7_97b30709,
        64'h07854721_93811782,
        64'h8fd98ff5_0107571b,
        64'h003f06b7_0107979b,
        64'h14068e63_02cba683,
        64'h090ba823_1408dc63,
        64'h090ba623_00d5183b,
        64'h8abd0107_d69b08db,
        64'ha22308db_a42304cb,
        64'ha823180b_ae231a0b,
        64'ha8238a05_00c7d61b,
        64'h02d606bb_018ba883,
        64'h45051086_a6830f86,
        64'h460396ce_964e068a,
        64'h8a3d41a9_89930000,
        64'h39978a9d_0036d61b,
        64'h00cbac23_4006061b,
        64'h40010637_a0294004,
        64'h06370ea6_1ee34511,
        64'h1aa60f63_450dbf05,
        64'h06fb9e23_478502fb,
        64'ha6238b85_41e7d79b,
        64'h048ba783_00fbac23,
        64'h400007b7_bfe91a50,
        64'h10ef0640_051312a9,
        64'h6ee31170_10ef8526,
        64'h0007cc63_048ba783,
        64'hf155842a_b36ff0ef,
        64'h855e4585_3e800913,
        64'h90810205_149313b0,
        64'h10ef4501_b16ff0ef,
        64'h855e0407_c163180b,
        64'h8c23048b_a7838082,
        64'h615d6db6_6d566cf6,
        64'h7c167bb6_7b567af6,
        64'h6a1a69ba_695a64fa,
        64'h741a70ba_8522d55d,
        64'h842ad99f_f0ef855e,
        64'ha031020b_a423f4fd,
        64'h34fd1005_03e3842a,
        64'haa0ff0ef_855e008c,
        64'h46014495_cf818b85,
        64'h1b8ba783_120500e3,
        64'h842aabaf_f0efc482,
        64'hc2be855e_008c479d,
        64'h460104f1_10234789,
        64'he7b5180b_8ca3198b,
        64'hc783c7b1_199bc783,
        64'h1cd010ef_45018baa,
        64'he3b54401_e6eeeaea,
        64'heee6f2e2_f6defada,
        64'hfed6e352_e74eeb4a,
        64'hef26f706_f3227161,
        64'h551cb585_84aab595,
        64'hfa100493_a10ff0ef,
        64'ha8050513_00005517,
        64'hd965c1cf_f0ef8522,
        64'h4585bfd1_18f40c23,
        64'h47850007_d663443c,
        64'hed09c34f_f0ef8522,
        64'h4581c04f_f0ef8522,
        64'h02f51f63_f9200793,
        64'hb55d18f4_0ca34785,
        64'h06041e23_d45c8b85,
        64'h41e7d79b_c43ccc18,
        64'h80010737_00e68563,
        64'h80020737_4c14bf45,
        64'h2ff010ef_3e800513,
        64'h06090863_397d0007,
        64'hca6347b2_ed1db8ef,
        64'hf0ef8522_858a4601,
        64'hc43e0197_e7b30187,
        64'h1563c43e_0177f7b3,
        64'hc25a4bdc_01511023,
        64'h4c18681c_e13dbb6f,
        64'hf0efc402_c2520131,
        64'h10238522_858a4601,
        64'h40000cb7_80020c37,
        64'h00ff8bb7_4b050290,
        64'h0a934a55_03700993,
        64'h3e900913_cc1c8002,
        64'h07b700f7_15630aa0,
        64'h079300c1_4703e911,
        64'hbf8ff0ef_c23ec43a,
        64'h8522858a_460147d5,
        64'h0aa00713_e3991aa0,
        64'h07138ff9_4bdc00ff,
        64'h8737681c_00f11023,
        64'h47a10005_05a345d0,
        64'h00ef8522_f14984aa,
        64'hcf2ff0ef_8522f1df,
        64'hf0ef8522_45814601,
        64'hb72ff0ef_8522d85c,
        64'h478508f4_22231a04,
        64'h28231804_2e230884,
        64'h2783f945_84aa9782,
        64'h6b9c679c_8522681c,
        64'h3ef010ef_7d000513,
        64'hba2ff0ef_85220204,
        64'h2c2302f4_08234785,
        64'h1af42c23_478df93f,
        64'hf0eff3e5_4481541c,
        64'h80826109_7ca27c42,
        64'h7be26b06_6aa66a46,
        64'h69e674a6_79068526,
        64'h744670e6_f8500493,
        64'hbacff0ef_c0450513,
        64'h00005517_02042423,
        64'heb8d6b9c_679c681c,
        64'hc509f11f_f0ef842a,
        64'hc17c8fd9_f466f862,
        64'hfc5ee0da_e4d6e8d2,
        64'heccef0ca_f4a6fc86,
        64'hf8a2070d_4b9c7119,
        64'h10000737_691c8082,
        64'h8082c2cf_f06f02c5,
        64'h0823dd0c_0007059b,
        64'h00e7f463_85be2781,
        64'h4f1887ae_00f5f363,
        64'h4f5c6918_ee09b7cd,
        64'hc402fef4_14e34785,
        64'h80826121_790274a2,
        64'h744270e2_d34ff0ef,
        64'h8526858a_4601c43e,
        64'h478900f4_1f634791,
        64'hc24a00f1_10234799,
        64'hed19d52f_f0efc43e,
        64'hc24a8526_858a4601,
        64'h0107979b_4955842e,
        64'h07c4d783_00f11023,
        64'h03700793_04f59263,
        64'h55294785_00f58663,
        64'h84aa4791_f04af822,
        64'hfc06f426_71398082,
        64'h01416402_60a24505,
        64'h83020141_60a26402,
        64'h85220003_07630187,
        64'hb303679c_681c0005,
        64'h5e63810f_f0ef842a,
        64'he406e022_1141b32d,
        64'hdd79842a_945ff0ef,
        64'h854a4585_0a700613,
        64'h86cebb3d_842a957f,
        64'hf0ef854a_458509b0,
        64'h06134685_01379b63,
        64'h0a7a4783_d4fb0de3,
        64'h4785ed19_975ff0ef,
        64'h854a4585_09c00613,
        64'h86defdb4_98e30c11,
        64'h0ff4f493_248dffac,
        64'h90e30ffa_fa932ca1,
        64'h2a85e139_99dff0ef,
        64'h854a0ff6_f6930196,
        64'hd6bb4585_8656000c,
        64'h26834c81_8aa609b0,
        64'h0d934d61_ffa492e3,
        64'h2ca10ff4_f4932485,
        64'he9359cbf_f0ef854a,
        64'h45858626_0ff6f693,
        64'h019ad6bb_08f00d13,
        64'h4c81ffb4_92e32d21,
        64'h0ff4f493_2485ed49,
        64'h9f1ff0ef_854a4585,
        64'h86260ff6_f69301ac,
        64'hd6bb08c0_0d934d01,
        64'h08800493_08f92a23,
        64'h00a7979b_0e0a4783,
        64'h0afa07a3_4785e569,
        64'ha21ff0ef_854a4585,
        64'h0af00613_4685e395,
        64'h8b850afa_4783e20b,
        64'h02e3b51d_547ddbaf,
        64'hf0efdf25_05130000,
        64'h5517cb89_8b8509ba,
        64'h4783bfd1_00f9f9b3,
        64'hfff7c793_b5912cc0,
        64'h20efdc25_05130000,
        64'h5517ef89_8b850a6a,
        64'h478302d9_8263fcc5,
        64'h92e3872e_0ff9f993,
        64'h00f9e9b3_c70d4189,
        64'hd99b4187_d79b8b05,
        64'h0189999b_0187979b,
        64'h0027571b_00b517bb,
        64'h02080463_00187813,
        64'h0017581b_4b189726,
        64'h070e0017_059b4611,
        64'h45054701_0016e993,
        64'hc3990fe6_f9938b89,
        64'hc71989b6_0017f713,
        64'h0a7a4683_0084c783,
        64'hb5c1e56f_f0efe0e5,
        64'h05130000_551785ce,
        64'h01367a63_963e09da,
        64'h47839e3d_0087979b,
        64'h0106161b_09ea4783,
        64'h09fa4603_ee0519e3,
        64'h842af94f_f0ef854a,
        64'h85d2fe0a_7a1302f1,
        64'h0a13f006_00e3e1e5,
        64'h05130000_55178a09,
        64'h000b8963_fbc596e3,
        64'h87ae0511_08210133,
        64'h09bb0ffb_fb9300db,
        64'hebb300be_96bbcb89,
        64'h8b850107_c78397a6,
        64'h078e0208_80630065,
        64'h202302e8_d33bb7f1,
        64'h4b814a81_4c81b7c1,
        64'hee4ff0ef_e3c50513,
        64'h00005517_00030d63,
        64'h02e8f33b_0017859b,
        64'h00082883_4e114e85,
        64'h478189d6_856200c4,
        64'h88138c0a_009c9c9b,
        64'he3994b85_02eadabb,
        64'h02c92783_bf415429,
        64'hf24ff0ef_e4450513,
        64'h00005517_cb8902ec,
        64'hf7bb0005_ac83e791,
        64'h02eaf7bb_060a8163,
        64'h0045aa83_db45e3e5,
        64'h05130000_55170989,
        64'h27038082_2a010113,
        64'h23813d83_24013d03,
        64'h24813c83_25013c03,
        64'h25813b83_26013b03,
        64'h26813a83_27013a03,
        64'h27813983_28013903,
        64'h28813483_29013403,
        64'h29813083_8522f840,
        64'h0413f96f_f0efe665,
        64'h05130000_5517e7b9,
        64'h00167793_07e94603,
        64'h00e7eb63_e4450513,
        64'h00005517_84ae8b32,
        64'h892abfe7_87933ffc,
        64'h07b79f3d_bff7879b,
        64'hbffc07b7_4d180ac7,
        64'he9634789_23b13c23,
        64'h25a13023_25913423,
        64'h25813823_25713c23,
        64'h27613023_27513423,
        64'h27413823_27313c23,
        64'h29213023_28913423,
        64'h28813823_28113c23,
        64'hd6010113_80826145,
        64'h69a26942_64e27402,
        64'h70a28522_013505a3,
        64'h15e010ef_8526842a,
        64'h875ff0ef_852685ca,
        64'h00091c63_00f51e63,
        64'h842a57b5_c519cc7f,
        64'hf0ef84aa_45850b30,
        64'h06138edd_892e9be1,
        64'h0079f693_0ff5f993,
        64'h08154783_f022f406,
        64'he44ee84a_ec267179,
        64'hb74d84aa_b75ddf40,
        64'h0493f7d5_0b944783,
        64'he51998df_f0ef854a,
        64'h85a29801_01f10413,
        64'hf1e92581_99f5ffe4,
        64'h059bf571_84aad1ff,
        64'hf0ef892a_45850b90,
        64'h0613842e_4685fef7,
        64'h60e34705_ffc5879b,
        64'h80822401_01132281,
        64'h34832201_39038526,
        64'h23013403_23813083,
        64'h54a9c585_468102b7,
        64'he16302f5_88634789,
        64'h23213023_22913423,
        64'h22813823_22113c23,
        64'hdc010113_bf455929,
        64'hbf555951_bf651a04,
        64'hb0235240_20efd169,
        64'h1a04b503_892abf4d,
        64'h08f4aa23_02f707bb,
        64'h27852705_8bfd8b7d,
        64'h0057d79b_00a7d71b,
        64'h50fc8082_25010113,
        64'h22813983_23013903,
        64'h23813483_854a2401,
        64'h34032481_308308f4,
        64'h80230a74_478308d4,
        64'hac2302f6_86bb00a6,
        64'h969b0dd4_4783f8dc,
        64'h07a60d44_27830009,
        64'h8663c799_54dc08f4,
        64'haa2300a6_979bc7b9,
        64'h8b850e04_46830af4,
        64'h47830af4_07a34785,
        64'hed35e0bf_f0ef8526,
        64'h45850af0_06134685,
        64'hce81e391_8bfd09c4,
        64'h4783c789_8b850a04,
        64'h4783f4fc_07a6c319,
        64'hf4fc54d8_9fb90884,
        64'h47039fb9_0087171b,
        64'h08944703_9fb90107,
        64'h171b0187_979b08a4,
        64'h470308b4_4783f8fc,
        64'h07ce02e7_87b30dd4,
        64'h478302f7_07330e04,
        64'h470397ba_08c44703,
        64'h9fb90087_171b0107,
        64'h979b4685_08d44703,
        64'h08e44783_04098f63,
        64'hfca714e3_0621070d,
        64'he21c07ce_02b787b3,
        64'h0dd44783_02f585b3,
        64'h0e044583_00098c63,
        64'h4685c391_97aeffe7,
        64'h45839fad_0105959b,
        64'h0087979b_00074583,
        64'hfff74783_e0fc07c6,
        64'h468109d4_05130a84,
        64'h4783fcdc_07c60c84,
        64'h86130914_07130e24,
        64'h478306f4_8fa309c4,
        64'h4783c789_8b890a04,
        64'h47830009_8a6308f4,
        64'h80a30b34_4783c789,
        64'h0e244783_e7810019,
        64'hf9938b85_06f48f23,
        64'h09b44983_0a044783,
        64'hf8dc00d7_73630147,
        64'hd69307a6_80070713,
        64'h67050d44_278300e7,
        64'hfd63cc98_1ff78793,
        64'h400407b7_53b897ba,
        64'h078ae0a7_07130000,
        64'h47171cf7_6b634721,
        64'h0c044783_123010ef,
        64'h85a22000_06131e05,
        64'h03631a04_b5031aa4,
        64'hb0236c20_20ef2000,
        64'h0513e799_1a04b783,
        64'h1e051863_892ac09f,
        64'hf0ef84aa_85a29801,
        64'h01f10413_1ce7f563,
        64'h49013ffc_07372331,
        64'h34232291_3c232481,
        64'h30232411_34239fb9,
        64'h23213823_bffc07b7,
        64'hdb010113_4d18bfcd,
        64'hfc79347d_80826121,
        64'h74a27442_70e2d91f,
        64'hf0ef8526_3e800593,
        64'he919c53f_f0ef8526,
        64'h858a4601_440dc436,
        64'h84aafc06_f426f822,
        64'h8ed10106_161b8edd,
        64'h030007b7_0086969b,
        64'hc23e47f5_00f11023,
        64'h47997139_80826121,
        64'h6aa26a42_69e274a2,
        64'h79028526_744270e2,
        64'hfc0999e3_9aa20287,
        64'h84339a22_408989b3,
        64'h08c96783_fc851ae3,
        64'hf01ff0ef_854a85d6,
        64'h865286a2_844e0089,
        64'hf3630207_e4030109,
        64'h378389a6_f96decdf,
        64'hf0ef854a_08c92583,
        64'ha0894481_bd9ff0ef,
        64'h24050513_00005517,
        64'h00b67a63_014485b3,
        64'h68100005_4d638dff,
        64'ha0ef8522_00b44583,
        64'hc11d892a_482010ef,
        64'h8ab684b2_8a2e4148,
        64'h842ace05_e456e852,
        64'hec4ef04a_f426f822,
        64'hfc067139_b7c54401,
        64'hb7d50004_841bb74d,
        64'h02f6063b_bf6147c5,
        64'h80826125_690664a6,
        64'h644660e6_8522c43f,
        64'hf0ef28a5_05130000,
        64'h5517c11d_d55ff0ef,
        64'hd23ed402_854a100c,
        64'h47f54601_02f11023,
        64'h47b10497_f0634785,
        64'he529842a_d75ff0ef,
        64'hc83eca26_d23a854a,
        64'h100c4785_0030cc3e,
        64'he42e4755_d432cf31,
        64'h08c92783_260102f1,
        64'h102302c9_270347c9,
        64'h06d7f663_84b6892a,
        64'h4785e8a2_ec86e0ca,
        64'he4a6711d_80824501,
        64'hbfd54501_80826121,
        64'h74a27442_70e2f8ed,
        64'h34fdc901_dcdff0ef,
        64'h8522858a_46014495,
        64'hcb918b89_1b842783,
        64'hc11dde3f_f0efc23e,
        64'h842af426_fc06f822,
        64'h858a4601_47d5c42e,
        64'h00f11023_47c17139,
        64'he7a919c5_2783bf7d,
        64'hf9200513_d09ff0ef,
        64'h33050513_00005517,
        64'hfc8049e3_4501b755,
        64'h5a6020ef_3e800513,
        64'h00f05763_0014079b,
        64'h347dfe04_c6e334fd,
        64'h80826125_7aa27a42,
        64'h79e26906_64a66446,
        64'h60e6fba0_0513d4bf,
        64'hf0ef35a5_05130000,
        64'h5517c78d_0125f7b3,
        64'h05479363_0135f7b3,
        64'hc7891005_f79345b2,
        64'hed0de73f_f0ef8556,
        64'h858a4601_e00a0a13,
        64'he0098993_08090913,
        64'h4495c43e_842e8aaa,
        64'hec86f456_e4a6e8a2,
        64'h6a056989_fdf94937,
        64'h0107979b_f852fc4e,
        64'he0ca07c5_5783c23e,
        64'h47d500f1_102347b5,
        64'h711d8082_61457402,
        64'h70a2c43c_47b2e119,
        64'hec9ff0ef_8522858a,
        64'h4601c43e_8fd98f55,
        64'h400006b7_8f756000,
        64'h06b78ff5_8ff9f807,
        64'h87934ad4_008007b7,
        64'h45386914_c195842a,
        64'hc402c23e_f406f022,
        64'h478500f1_10234785,
        64'h71798082_61457402,
        64'h70a28522_69a020ef,
        64'h7d000513_e509842a,
        64'hf21ff0ef_c202c402,
        64'h00011023_858a4601,
        64'h85226b80_20eff406,
        64'h3e800513_842af022,
        64'h7179b761_fb600513,
        64'hd55156f0_10ef0d44,
        64'h85130d44_05934611,
        64'h00f71a63_0e044783,
        64'h0e04c703_02f71063,
        64'h0c044783_0c04c703,
        64'h02f71663_0dd44783,
        64'h0dd4c703_02f71c63,
        64'h0a044783_0a04c703,
        64'hf579f95f_f0ef1a05,
        64'h34832211_3c232291,
        64'h342385a2_980101f1,
        64'h04132281_3823dc01,
        64'h01138082_24010113,
        64'h22813483_23013403,
        64'h23813083_45018082,
        64'h450100e6_fe634004,
        64'h07374d14_80826161,
        64'h60a6fd3f_f0efcc3e,
        64'hd402e486_100c2000,
        64'h07930030_e83ee42e,
        64'h07851782_4785d23e,
        64'h47d502f1_102347a1,
        64'h715d8302_0007b303,
        64'h679c691c_80824fe5,
        64'h05130000_55178082,
        64'h6108953e_817525e7,
        64'h87930000_47971502,
        64'h00a7eb63_47ad8082,
        64'h557d8082_01416402,
        64'h60a24501_83020141,
        64'h60a26402_85220003,
        64'h07630207_b303679c,
        64'h681c0005_5e63ff5f,
        64'hf0ef842a_e406e022,
        64'h11418082_557d8082,
        64'h557db7e9_659c95aa,
        64'h058e05e1_35f1bfd9,
        64'h617cbfe9_7d5c8082,
        64'h61054501_e91c64a2,
        64'h644260e2_02f457b3,
        64'h93810204_97930c50,
        64'h10ef7540_f55c08c5,
        64'h2483795c_878297ba,
        64'he426e822_ec061101,
        64'h439c97ba_83f92d67,
        64'h07130000_47170205,
        64'h979304b7_ee63479d,
        64'h80824501_83020003,
        64'h03630087_b303679c,
        64'h691c8082_61356452,
        64'h60f28522_0f7020ef,
        64'h0808842a_e3fff0ef,
        64'he436eec6_eac2e6be,
        64'he2baea22_ee060808,
        64'h10000593_1234862a,
        64'hfe36fa32_f62e710d,
        64'h80826161_60e2e69f,
        64'hf0efe436_e4c6e0c2,
        64'hfc3ef83a_ec061000,
        64'h05931014_862ef436,
        64'hf032715d_80826161,
        64'h60e2e8df_f0efe436,
        64'he4c6e0c2_fc3ef83a,
        64'hec061034_f436715d,
        64'hb7f18522_02010393,
        64'h0005059b_4db010ef,
        64'h85220124_74336000,
        64'h00840b13_b5fd845a,
        64'hd93ff0ef_00840b13,
        64'h02010393_00044503,
        64'ha809ddbf_f0ef0028,
        64'h02010393_0005059b,
        64'he37ff0ef_400845a9,
        64'h46010016_b6930038,
        64'h00840b13_f8b50693,
        64'ha81145c1_00163613,
        64'h46850038_00840b13,
        64'hfa850613_f6e510e3,
        64'h07800713_02e50063,
        64'h07500713_a00d4601,
        64'h46850038_00840b13,
        64'hf6e51ee3_07000713,
        64'h00a76c63_06e50e63,
        64'h07300713_b74d048d,
        64'h0024c503_80826109,
        64'h0007051b_6b066aa6,
        64'h6a4669e6_790674a6,
        64'h744670e6_f55d08f5,
        64'h09630630_079304d5,
        64'h0f630580_069302a6,
        64'heb6306d5_0f630640,
        64'h06930489_0014c503,
        64'h478100f6_f36346a5,
        64'h0ff7f793_fd07879b,
        64'hcb9d0004_c7830355,
        64'h10634781_04890545,
        64'h0f630014_c503bfe1,
        64'he7bff0ef_02010393,
        64'h04850135_086304d7,
        64'hff639381_17827682,
        64'h0017079b_c52d8f1d,
        64'h0004c503_77a27742,
        64'h02095913_03000a93,
        64'h06c00a13_02500993,
        64'hf82af02e_f42afc3e,
        64'h843684b2_e0dafc86,
        64'he4d6e8d2_eccef4a6,
        64'hf8a2597d_011cf0ca,
        64'h7119b7f1_06850117,
        64'h80230066_80232605,
        64'h0006c883_0007c303,
        64'h97ba9381_178240c8,
        64'h07bbb7d9_2585fea6,
        64'h8fa30685_bf5d00a8,
        64'h053b8082_00b61b63,
        64'hfff5081b_86ba2581,
        64'h00068023_0015559b,
        64'h40e6853b_068500f6,
        64'h802302d0_07930008,
        64'h876302f5_e9630300,
        64'h051340e6_85bbfe71,
        64'h8532fea6_8fa30685,
        64'h0ff57513_02b6563b,
        64'h0305051b_046e6763,
        64'h0ff37513_02b6733b,
        64'h0005061b_385986ba,
        64'h4e250ff6_f8130410,
        64'h0693c219_06100693,
        64'h488540a0_053be681,
        64'h00055663_4881bfe9,
        64'h00d70023_07850007,
        64'hc68300d3_b8230017,
        64'h06938082_852e0007,
        64'h002300b6_e6630103,
        64'hb70340a7_86bb87aa,
        64'h9d9dfff7_059b00c6,
        64'hf5638e9d_fff70693,
        64'h0003b703_8f999201,
        64'h02059613_0103b783,
        64'h0083b703_80824501,
        64'h80820007_80234505,
        64'h0103b783_00a70023,
        64'h00f3b823_00170793,
        64'h00d7fe63_93811782,
        64'h278540f7_07b30003,
        64'hb6830083_b7830103,
        64'hb7038082_61454501,
        64'h6a0269a2_694264e2,
        64'h740270a2_2e8000ef,
        64'he2050513_00006517,
        64'hfd249fe3_04052fa0,
        64'h00ef8191_00f5f613,
        64'h2485854e_00044583,
        64'h30c000ef_855285a6,
        64'he78901f4_f7932000,
        64'h09139029_89930000,
        64'h6997902a_0a130000,
        64'h6a174481_ed5ff0ef,
        64'h84264581_852633a0,
        64'h00ef9025_05130000,
        64'h6517bda6_06130000,
        64'h6617e789_87c60613,
        64'h00006617_584c19c4,
        64'h2783db5f_b0efe965,
        64'h85930000_65977448,
        64'h05e030ef_92450513,
        64'h00006517_378000ef,
        64'h91850513_00006517,
        64'h8a058593_00006597,
        64'hc7898b25_85930000,
        64'h6597545c_398000ef,
        64'h92850513_00006517,
        64'h5c0c3a60_00ef2601,
        64'h0ff6f693_0ff7f793,
        64'h0ff77713_0187d61b,
        64'h0107d69b_0087d71b,
        64'h93850513_00006517,
        64'h06c44583_583c3d20,
        64'h00ef91c1_15c20085,
        64'hd59b9425_05130000,
        64'h6517546c_3e8000ef,
        64'h93850513_00006517,
        64'h06f44583_3f8000ef,
        64'h638c93a5_05130000,
        64'h6517681c_206010ef,
        64'h842a4910_10ef4501,
        64'h44b010ef_0001b503,
        64'h10e030ef_95450513,
        64'h00006517_84aa0060,
        64'h30efe052_e44ee84a,
        64'hec26f022_f4062000,
        64'h05137179_7940006f,
        64'h61054685_60e26622,
        64'h644285a2_4d3010ef,
        64'he42eec06_4501842a,
        64'he8221101_80820141,
        64'h640260a2_557de391,
        64'h4505703c_0cc030ef,
        64'h8f050513_00006517,
        64'h8e058593_00006597,
        64'h34c00613_77c68693,
        64'h00004697_02f40263,
        64'h200007b7_e4066380,
        64'he0221141_711c8082,
        64'h25016108_953e050e,
        64'h200007b7_f73ff06f,
        64'h20000537_45814609,
        64'h8082bff9_557d0e80,
        64'h30ef8522_b7e5c45c,
        64'h4785d4fd_45018885,
        64'h80826145_69a26942,
        64'h64e27402_70a24501,
        64'hc45c4789_cb990024,
        64'hf793f404_01242423,
        64'he01c2000_07b70209,
        64'h8b634fe0_00ef9fe5,
        64'h05130000_65178622,
        64'h85aa89aa_785010ef,
        64'h7e050513_00004517,
        64'h85a2cc1d_5551842a,
        64'h100030ef_892e84b2,
        64'he44ef406_e84aec26,
        64'hf0220480_05137179,
        64'h08b04163_5535b7dd,
        64'h87ca0ca1_39a020ef,
        64'he43e002c_46218566,
        64'h639c0087_8913fa97,
        64'h8de394be_00093c83,
        64'h01096483_97a667a1,
        64'hbf41b1df_f0ef8522,
        64'hb77100f9_2623000c,
        64'hb783dbd9_8b85bd95,
        64'h60f020ef_4505d80c,
        64'h8ee3c47f_f0ef8522,
        64'h484cc85c_9bf54c85,
        64'h485cb4df_f0ef8522,
        64'hef8d8b85_00892783,
        64'h00090963_04043023,
        64'h210030ef_855685d2,
        64'h0ca00613_87468693,
        64'h00005697_01748c63,
        64'h04043903_6004cc9d,
        64'h4c858889_c85c9bf9,
        64'h485cc85c_0027e793,
        64'h485ccbb5_603cfeb6,
        64'h90e30791_872a2685,
        64'hc3988f51_8361ff87,
        64'h37030106_8763c390,
        64'h0086161b_ff870513,
        64'h63104591_480d4681,
        64'h00c90793_018c8713,
        64'h08e69f63_0037f693,
        64'h470d0204_3c230049,
        64'h2783cba9_7c1c28e0,
        64'h30ef8556_85d209c0,
        64'h06138da6_86930000,
        64'h5697017c_8c630384,
        64'h39030004_3c83cfb5,
        64'h0014f793_658000ef,
        64'hb3050513_00006517,
        64'h85cad1ff_f0ef85ca,
        64'h00496913_ff397913,
        64'h85220144_2903c395,
        64'h0084f793_680000ef,
        64'hb3050513_00006517,
        64'h85cad47f_f0ef85ca,
        64'h00896913_ff397913,
        64'h85220144_2903c395,
        64'h0044f793_b27ff0ef,
        64'h85224581_b6fff0ef,
        64'h85224581_cc5cf920,
        64'h0793c781_7c1c00f7,
        64'h6f630c89_37830209,
        64'h37031204_8e632481,
        64'h8cfd4c81_485c0709,
        64'h348333a0_30ef8556,
        64'h85d20f20_061386e2,
        64'h01790963_00043903,
        64'hb7116f60_00efb8e5,
        64'h05130000_651796e5,
        64'h85930000_5597000b,
        64'h1d633b7d_20000bb7,
        64'h8b4ebd61_00c4e493,
        64'hbd8537a0_30efb9e5,
        64'h05130000_6517b8e5,
        64'h85930000_65971490,
        64'h061398a6_86930000,
        64'h5697b765_47014781,
        64'h2585e31c_97469381,
        64'h83751782_170200be,
        64'h873b8fd9_8fe90107,
        64'h67330087_d79b01c8,
        64'h78330087_981b0107,
        64'h67330187_971b0187,
        64'hd81bf2e5_00670363,
        64'h16fd0605_27810107,
        64'he7b301e8_183b0705,
        64'h00371f1b_00064803,
        64'hec0689e3_6e89f005,
        64'h051300ff_0e374311,
        64'h47014781_45816390,
        64'h0107e683_65410004,
        64'h3883603c_ee079be3,
        64'h8b85449c_df3ff0ef,
        64'h8522488c_db7ff0ef,
        64'he0248522_44cc8082,
        64'h61654501_6ce27c02,
        64'h7ba27b42_7ae26a06,
        64'h69a66946_64e67406,
        64'h70a6efe9_485cc6ea,
        64'h8a930000_6a976819,
        64'h8993eb7f_f0ef2581,
        64'h0015e593_009899b7,
        64'h85220d89_b583cd1f,
        64'hf0ef8522_4585e93f,
        64'hf0ef8522_24058593,
        64'h000f45b7_d27ff0ef,
        64'h85224581_46054685,
        64'h4705cf5f_f0ef8522,
        64'h4581cbdf_f0ef8522,
        64'h85a6c81f_f0efcaea,
        64'h0a130000_6a178522,
        64'h00095583_c4fff0ef,
        64'hae8c0c13_00005c17,
        64'h85220089_2583be1f,
        64'hf0ef8522_4581d71f,
        64'hf0ef8522_45814605,
        64'h46814705_0144e493,
        64'h16078663_8b85008a,
        64'h2783000a_09638cdd,
        64'h03243c23_4c1c4485,
        64'he391448d_8b89c709,
        64'h0017f713_44810049,
        64'h278316f9_9a630404,
        64'h3a032000_07b70004,
        64'h3983bf5f_f0ef4585,
        64'h60080e04_9c636ca0,
        64'h20ef00c9_05134581,
        64'h4611d01c_e03084b2,
        64'h892e0005_d7830204,
        64'h08a3ec66_f062f45e,
        64'hf85afc56_e0d2e4ce,
        64'hf486e8ca_eca67100,
        64'hf0a27159_80826105,
        64'h690264a2_644260e2,
        64'hc8440499_3c2356e0,
        64'h30efd925_05130000,
        64'h6517d825_85930000,
        64'h65970760_0613b6e6,
        64'h86930000_569702f9,
        64'h026384ae_842a2000,
        64'h07b7ec06_e426e822,
        64'h00053903_e04a1101,
        64'h80826105_64a26442,
        64'h60e2e424_5b4030ef,
        64'hdd850513_00006517,
        64'hdc858593_00006597,
        64'h06f00613_ba468693,
        64'h00005697_02f40263,
        64'h84ae2000_07b7ec06,
        64'he4266100_e8221101,
        64'h80826105_64a26442,
        64'h60e2e0a0_8c7d17fd,
        64'h67855fa0_30efe1e5,
        64'h05130000_6517e0e5,
        64'h85930000_65970680,
        64'h0613bda6_86930000,
        64'h569702f4_8263842e,
        64'h200007b7_ec06e822,
        64'h6104e426_11018082,
        64'h610564a2_644260e2,
        64'hfc809041_144263e0,
        64'h30efe625_05130000,
        64'h6517e525_85930000,
        64'h65970610_0613c0e6,
        64'h86930000_569702f4,
        64'h8263842e_200007b7,
        64'hec06e822_6104e426,
        64'h1101d4df_f06f0141,
        64'h458160a2_64026008,
        64'hf23ff0ef_46054685,
        64'h47054581_8522ef1f,
        64'hf0ef4581_8522f39f,
        64'hf0ef842a_45810405,
        64'h30230205_3c234605,
        64'h46814705_e022e406,
        64'h11418082_01414501,
        64'h640260a2_d97ff0ef,
        64'h45816008_f67ff0ef,
        64'h45814605_46854705,
        64'h8522f35f_f0ef4581,
        64'h8522f7df_f0efe406,
        64'h45818522_46054681,
        64'h47057100_e0221141,
        64'h80826121_69e27902,
        64'h74a202b9_b8238dc5,
        64'h744270e2_88a10125,
        64'he5b30034_949b8dd9,
        64'h00497913_0029191b,
        64'h8b058989_0014159b,
        64'h67227220_30efe43a,
        64'hf4850513_00006517,
        64'hf3858593_00006597,
        64'h05a00613_ce468693,
        64'h00005697_02f98463,
        64'h84368932_84ae2000,
        64'h07b7fc06_f04af426,
        64'hf8220005_3983ec4e,
        64'h71398082_610564a2,
        64'h644260e2_f40476e0,
        64'h30eff925_05130000,
        64'h6517f825_85930000,
        64'h65970530_0613d1e6,
        64'h86930000_569702f4,
        64'h026384ae_200007b7,
        64'hec06e426_6100e822,
        64'h11018082_610564a2,
        64'h644260e2_f0047ae0,
        64'h30effd25_05130000,
        64'h6517fc25_85930000,
        64'h659704c0_0613d4e6,
        64'h86930000_569702f4,
        64'h026384ae_200007b7,
        64'hec06e426_6100e822,
        64'h11018082_610564a2,
        64'h644260e2_ec809001,
        64'h14027f20_30ef0165,
        64'h05130000_65170065,
        64'h85930000_65970450,
        64'h0613c626_86930000,
        64'h769702f4_8263842e,
        64'h200007b7_ec06e822,
        64'h6104e426_11018082,
        64'h610564a2_644260e2,
        64'he8809001_14020370,
        64'h30ef05a5_05130000,
        64'h651704a5_85930000,
        64'h659703e0_0613cae6,
        64'h86930000_769702f4,
        64'h8263842e_200007b7,
        64'hec06e822_6104e426,
        64'h11018082_610564a2,
        64'h644260e2_e4040770,
        64'h30ef09a5_05130000,
        64'h651708a5_85930000,
        64'h65970360_0613e066,
        64'h86930000_569702f4,
        64'h026384ae_200007b7,
        64'hec06e426_6100e822,
        64'h11018082_610564a2,
        64'h644260e2_e0040b70,
        64'h30ef0da5_05130000,
        64'h65170ca5_85930000,
        64'h659702f0_0613e366,
        64'h86930000_569702f4,
        64'h026384ae_200007b7,
        64'hec06e426_6100e822,
        64'h11018082_610564a2,
        64'h644260e2_fc240f70,
        64'h30ef11a5_05130000,
        64'h651710a5_85930000,
        64'h65970880_0613e5e6,
        64'h86930000_569702f5,
        64'h026384ae_842a2000,
        64'h07b7ec06_e426e822,
        64'h11018082_556dbfe5,
        64'h0007ac23_80824501,
        64'hcf980200_071300d7,
        64'h17634691_00d70d63,
        64'h711c46a1_59588082,
        64'h6149640a_60aaf83f,
        64'hf0ef0808_f01ff0ef,
        64'h0808e85f_f0ef0808,
        64'h85a26622_f71ff0ef,
        64'he42ee506_0808842a,
        64'he1227175_80826105,
        64'hf3050513_00007517,
        64'h60e2fca7_1de3fef6,
        64'h8fa3fec6_8f230007,
        64'hc78397ae_00064603,
        64'h8bbd962e_0047d613,
        64'h07050689_0007c783,
        64'h00e107b3_45411a65,
        64'h85930000_6597f6e6,
        64'h86930000_76974701,
        64'h3bf020ef_ec06850a,
        64'h46410505_05931101,
        64'h8082e13c_b6c78793,
        64'h00000797_ed3c639c,
        64'hd2878793_00007797,
        64'he93c0405_3423639c,
        64'hd3078793_00007797,
        64'h80826145_69a26942,
        64'h64e27402_70a2fd24,
        64'hfde34501_97828522,
        64'h603cfc1c_078e643c,
        64'h0124f563_3c9020ef,
        64'h95224581_92011602,
        64'h0006091b_40a9863b,
        64'h449d0400_099300e7,
        64'h802397a2_f8000713,
        64'h00178513_e84af406,
        64'he44eec26_842a03f7,
        64'hf793f022_7179653c,
        64'h80826161_6ba26b42,
        64'h6ae27a02_79a27942,
        64'h74e26406_60a6b7c9,
        64'h97824401_852660bc,
        64'h01741763_99d64159,
        64'h09334810_20ef0144,
        64'h043b8656_00848533,
        64'h85ce020a_da93020a,
        64'h1a930009_0a1b00f9,
        64'h74639381_17820007,
        64'h8a1b408b_07bb0400,
        64'h0b930400_0b13e53c,
        64'h893289ae_84aa97b2,
        64'h03f7f413_ec56f052,
        64'he486e45e_e85af44e,
        64'hf84afc26_e0a2715d,
        64'h653c8082_61056922,
        64'h64c2cd70_cd34c97c,
        64'h05052823_00c8863b,
        64'h00d306bb_00fe07bb,
        64'h010e883b_6462f3ef,
        64'h9de300e5_87bb0005,
        64'h869b0003_861b0f11,
        64'h8f5d0157_171b00b7,
        64'h579b9f3d_00774733,
        64'h9fa18f4d_fff74713,
        64'h0007081b_00b385bb,
        64'h40809fa1_8dd50115,
        64'hd59b94aa_00f5969b,
        64'h048a9db5_ffc2a403,
        64'h8db902c1_0075e5b3,
        64'hfff7c593_023f4483,
        64'h9ead00c7_03bb00c3,
        64'he633400c_9ead0166,
        64'h561b00a6_139b0082,
        64'ha5839e2d_8e3d8e59,
        64'hfff6c613_9db100f8,
        64'h073b0107_683301a8,
        64'h581b0003_a5839e2d,
        64'h0068171b_0107083b,
        64'h0042a583_9f2d942a,
        64'h040a418c_95aa058a,
        64'h93aa038a_020f4583,
        64'h9f2d022f_4403021f,
        64'h43830002_a70300d7,
        64'h45b38f5d_fff64713,
        64'h0b028293_00005297,
        64'hf5f592e3_00e407bb,
        64'h0004069b_0002861b,
        64'h0f918f5d_0177171b,
        64'h0097579b_9f3d8f21,
        64'h9fa50057_47330007,
        64'h081b00d2_843b8ec1,
        64'h00092483_0106d69b,
        64'h9fa50106_941b992a,
        64'h9ea1090a_0056c6b3,
        64'h00e7c6b3_ffc3a483,
        64'h9c3500c7_02bb03c1,
        64'h00c2e633_0156561b,
        64'h013fc903_00b6129b,
        64'h408000c2_863b9ea1,
        64'h94aa00e2_c2b3048a,
        64'h00f8073b_0083a403,
        64'h9e210107_683301c8,
        64'h581b0048_171b012f,
        64'hc4830107_083b4080,
        64'h9e2194aa_048a0043,
        64'ha4039f21_011fc483,
        64'h9f254000_00c2c4b3,
        64'h942a040a_00d7c2b3,
        64'h0003a703_010fc403,
        64'h13838393_00005397,
        64'h8ffa1c2f_0f130000,
        64'h5f17f255_99e300e4,
        64'h07bb0004_069b0003,
        64'h861b000f_081b8f5d,
        64'h0147171b_00c7579b,
        64'h9f3d0077_473301e7,
        64'h77330083_c7339fb9,
        64'h00d3843b_8ec14098,
        64'h0126d69b_9fb900e6,
        64'h941b94aa_048affcf,
        64'ha7039eb9_0fc101e6,
        64'hc6b3fff5_c4838efd,
        64'h007f46b3_05919f35,
        64'h00cf03bb_00c3e633,
        64'h40189eb9_0176561b,
        64'h0096139b_008fa703,
        64'h9e398e3d_8e7501e7,
        64'hc6339f31_00f80f3b,
        64'h010f6833_0003a703,
        64'h01b8581b_9e390058,
        64'h1f1b010f_083b004f,
        64'ha70300ef_0f3b942a,
        64'h040a4318_972a070a,
        64'h93aa038a_0005c703,
        64'h00ef0f3b_0025c403,
        64'h0015c383_000faf03,
        64'h01e6c733_00cf7f33,
        64'h00d7cf33_2ac28293,
        64'h00005297_1e4f8f93,
        64'h00005f97_2ac58593,
        64'h00005597_f45f17e3,
        64'h00e387bb_0003869b,
        64'h0005881b_0f418f5d,
        64'h0167171b_00a7579b,
        64'h9f3d8f2d_9fa10077,
        64'h77338f2d_0007061b,
        64'h00d703bb_ffcfa403,
        64'h9fa100d3_e6b30116,
        64'h969b00f6_d39b0076,
        64'h86bb8ebd_00cf2403,
        64'h8ef900b7_c6b300d3,
        64'h83bb00c5_873b0083,
        64'h83bb8e59_0146561b,
        64'h00c6171b_9e39008f,
        64'h23838e35_8e6d00f6,
        64'hc6339f31_00f805bb,
        64'h0077073b_0105e833,
        64'h0198581b_0078159b,
        64'h0105883b_004f2703,
        64'hff4fa383_9db90075,
        64'h85bb0fc1_008fa403,
        64'h000f2583_000fa383,
        64'h00b64733_8dfd00c6,
        64'hc5b326af_8f930000,
        64'h5f978876_87f2869a,
        64'h86460405_02938f2a,
        64'he44ae826_ec221101,
        64'h05c52883_05852303,
        64'h05452e03_05052e83,
        64'hbf89eaf7_1de30e50,
        64'h07930181_4703f8d7,
        64'h71e30007_869b0200,
        64'h06134729_93811782,
        64'hf4c7e5e3_05850685,
        64'h00e58023_f91780e3,
        64'hb751842a_bf1900e7,
        64'h85a34721_6786ae5f,
        64'hd0ef082c_462d6506,
        64'hb07fd0ef_45810200,
        64'h06136506_f4450005,
        64'h041ba55f_e0ef1028,
        64'hdbd50181_478302f5,
        64'h1b634791_b7c10005,
        64'h041b8fef_e0ef00f5,
        64'h02234785_752200f5,
        64'h00235795_a8850785,
        64'h00c68023_00fe06b3,
        64'hb7cdffe8_1be30608,
        64'h05630005_48030505,
        64'hbfcdf36d_80826125,
        64'h644660e6_85224419,
        64'h00eef863_a8210007,
        64'h0f1b7125_05130000,
        64'h65179341_17423701,
        64'h00a36c63_91411542,
        64'hf9f7051b_27850006,
        64'hc70348b1_07f00e93,
        64'h43658e2e_4781082c,
        64'hfeb706e3_00074703,
        64'h97369301_02079713,
        64'hfff6079b_bf45863e,
        64'hb74d2605_a06100e7,
        64'h8ca30007_8ba30007,
        64'h8b230460_071300e7,
        64'h8c230210_07136786,
        64'hbc7fd0ef_082c462d,
        64'hc3dd6506_01814783,
        64'he1792501_abbfe0ef,
        64'h10284585_e8410005,
        64'h041bbd6f_e0efda02,
        64'h10284581_ea290200,
        64'h0593eba1_0007c783,
        64'h97b69381_02061793,
        64'h46010001_0c2366a2,
        64'hec550005_041bee3f,
        64'hd0efec86_e8a21028,
        64'h002c4605_e42a711d,
        64'hb7d5842a_bf550004,
        64'h802300f5_15634791,
        64'h80826125_690664a6,
        64'h644660e6_852200a9,
        64'h2023c29f_d0ef953e,
        64'h03478793_02700793,
        64'h00e68463_00054683,
        64'h04300793_470d6562,
        64'he0150005_041be69f,
        64'hd0ef510c_65620209,
        64'h0a63fec7_83e3177d,
        64'h0007c783_97a69381,
        64'h17820007_869bfff6,
        64'h879bce89_00070023,
        64'h02000613_46ad00b4,
        64'h8713ca1f_d0ef8526,
        64'h462d75c2_e93d2501,
        64'hb8ffe0ef_08284585,
        64'he5592501_ca8fe0ef,
        64'hd2020828_4581c4b9,
        64'he0510005_041bf9bf,
        64'hd0efec86_e8a20828,
        64'h4601002c_893284ae,
        64'he42ae0ca_e4a6711d,
        64'h80826125_644660e6,
        64'h2501ad6f_e0ef00f5,
        64'h02234785_00e78ca3,
        64'h0087571b_00e78c23,
        64'h00445703_00e78ba3,
        64'h0087571b_00e78b23,
        64'h75220064_5703cb85,
        64'h6786eb95_0207f793,
        64'h00b7c783_451967a6,
        64'he1292501_9abfe0ef,
        64'he4be1028_083c65a2,
        64'he9292501_810fe0ef,
        64'hec861028_002c4605,
        64'h842ee42a_e8a2711d,
        64'hbfcd47a1_8082614d,
        64'h853e64ea_740a70aa,
        64'h0005079b_b50fe0ef,
        64'h6506e791_0005079b,
        64'he24fe0ef_008800f7,
        64'h022306d7_07a34785,
        64'h06f704a3_0086d69b,
        64'h0106d69b_0087d79b,
        64'h0107d79b_0107979b,
        64'h06f70423_27810107,
        64'hd79b06f7_07230107,
        64'h969b57d6_02f69d63,
        64'h05574683_02e00793,
        64'h6706efb1_0005079b,
        64'hfc3fd0ef_8522c5a5,
        64'h47890005_059bcaef,
        64'he0ef8522_0005059b,
        64'hf2dfd0ef_85a60004,
        64'h450306f7_086357d6,
        64'h4736cbbd_8bc100b4,
        64'hc78300f4_02234785,
        64'h00f485a3_0207e793,
        64'h64060281_4783e0df,
        64'hd0ef00d4_851302a1,
        64'h0593464d_648aefc5,
        64'h0005079b_dc5fe0ef,
        64'h10a80ce7_93634711,
        64'hcbf90005_079baadf,
        64'he0ef10a8_65820c05,
        64'h4d6347ad_f05fd0ef,
        64'h850ae49f_d0ef10a8,
        64'h008c0280_0613e55f,
        64'hd0ef1028_05ad4655,
        64'h0e058e63_479165e6,
        64'h10071263_02077713,
        64'h479900b7_c7037786,
        64'h10079a63_0005079b,
        64'haf7fe0ef_f0be083c,
        64'hf4be0088_65a26786,
        64'h12079663_0005079b,
        64'h964fe0ef_ed26f122,
        64'hf5060088_002c4605,
        64'he02ee42a_71718082,
        64'h616564e6_740670a6,
        64'h2501c9ef_e0ef00f5,
        64'h02234785_008705a3,
        64'h8c3d0274_74138c65,
        64'h8cbd7522_00b74783,
        64'hc30d6706_e39d0207,
        64'hf79300b7_c7834519,
        64'h67a6e915_2501b65f,
        64'he0efe4be_1028083c,
        64'h65a2e131_25019caf,
        64'he0eff486_10284605,
        64'h002c8432_84aee42a,
        64'heca6f0a2_7159b7c5,
        64'h44218082_614d6d46,
        64'h6ce67c06_7ba67b46,
        64'h7ae66a0a_69aa694a,
        64'h64ea740a_70aa8522,
        64'hf25fe0ef_85ca7522,
        64'h441db749_8c6a0ffb,
        64'hfb93f61f_d0ef3bfd,
        64'h85524581_20000613,
        64'hec090005_041b8dcf,
        64'he0ef0195_02230385,
        64'h2823001c_0d1b7522,
        64'ha82d0005_041bd5af,
        64'he0ef00f5_02234785,
        64'h00978aa3_01678a23,
        64'h01378da3_01578d23,
        64'h00e78ca3_00078ba3,
        64'h00078b23_04600713,
        64'h00e78c23_02100713,
        64'h00e785a3_75224741,
        64'h6786e835_0005041b,
        64'hf59fe0ef_1028040b,
        64'h99634c85_00274b83,
        64'h06f404a3_06d407a3,
        64'h0087d79b_0086d69b,
        64'h0107d79b_0106d69b,
        64'h0107979b_06f40423,
        64'h27810107_d79b0107,
        64'h969b06f4_07234781,
        64'h00f69363_571400d6,
        64'h166357d2_00074603,
        64'h468d0574_0aa37722,
        64'h80efe0ef_05440513,
        64'h85d20494_04a30564,
        64'h04230534_07a30554,
        64'h07230404_05a30404,
        64'h05230374_0a230200,
        64'h061304f4_06a30084,
        64'hd49b0089_d99b0460,
        64'h07930ff9_7a9304f4,
        64'h062302e0_0b930104,
        64'hd49b0210_07930109,
        64'hd99b02f4_0fa30104,
        64'h949b0109_199b0ff4,
        64'hfb1347c1_248188cf,
        64'he0ef8552_02000593,
        64'h462d898f_e0ef8552,
        64'h00050c1b_45812000,
        64'h06130344_0a13f6ef,
        64'he0ef8522_0109549b,
        64'h85ca7422_16041463,
        64'h0005041b_a98fe0ef,
        64'h752216f9_0b634405,
        64'h57fd16f9_0f634409,
        64'h47851809_02630005,
        64'h091bb45f_e0ef4581,
        64'h75221807_9f630207,
        64'hf79300b7_c7834419,
        64'h67a61af4_17634791,
        64'h1c040963_0005041b,
        64'hd67fe0ef_e4be1028,
        64'h083c65a2_1c041463,
        64'h0005041b_bd0fe0ef,
        64'he8eaece6_f0e2f4de,
        64'hf8dafcd6_e152e54e,
        64'he94aed26_f506f122,
        64'h1028002c_4605e42a,
        64'h7171b769_d5752501,
        64'h91cff0ef_85a27502,
        64'hbf612501_f20fe0ef,
        64'h7502e411_f1552501,
        64'h9f5fe0ef_1008faf5,
        64'h18e34791_d94d2501,
        64'h836ff0ef_00a84581,
        64'hf1612501_951fe0ef,
        64'hcaa200a8_458996cf,
        64'he0ef00a8_100c0280,
        64'h0613fc87_8de30149,
        64'h2783c89d_88c1cc0d,
        64'h0005041b_ad8fe0ef,
        64'h00094503_79028082,
        64'h61497946_74e6640a,
        64'h60aa451d_cb810014,
        64'hf79300b5_c483c599,
        64'h75e2eb89_0207f793,
        64'h00b7c783_45196786,
        64'he1052501_e3bfe0ef,
        64'he0be1008_081c65a2,
        64'he9052501_ca0fe0ef,
        64'hf8cafca6_e122e506,
        64'h1008002c_4605e42a,
        64'h7175b7b1_00f40523,
        64'hfbf7f793_00a44783,
        64'hf55d2501_648040ef,
        64'h03040593_0017c503,
        64'h46854c50_601cdba5,
        64'h0407f793_00a44783,
        64'hfcf96ae3_4d1c6008,
        64'hfcf900e3_45094785,
        64'hb769449d_b7e12501,
        64'ha1cff0ef_85ca6008,
        64'hf9792501_b37fe0ef,
        64'h167d1000_06374c0c,
        64'hb7dd4505_02f91463,
        64'h57fd0005_091b94df,
        64'he0ef4c0c_bf7d84aa,
        64'h00a405a3_c5390004,
        64'h2a232501_a58ff0ef,
        64'h484cef01_600800f4,
        64'h0523c818_0207e793,
        64'hfed772e3_48144458,
        64'hcf390027_f71300a4,
        64'h47838082_610564a2,
        64'h69028526_644260e2,
        64'h0007849b_cb9100b4,
        64'h4783e491_0005049b,
        64'hbc4fe0ef_842ae04a,
        64'hec06e426_e8221101,
        64'hbfad8a2a_bfbd4a09,
        64'hb7494a05_b7c539f1,
        64'h09112485_e1116582,
        64'h01557533_2501abcf,
        64'he0efe02e_854ab745,
        64'hfc0c94e3_3cfd39f9,
        64'h09092485_e3918fd9,
        64'h0087979b_00094703,
        64'h00194783_038b9163,
        64'h20000993_03440913,
        64'h85cee921_2501d10f,
        64'he0ef0015_899b8522,
        64'h00099e63_1afd4c09,
        64'h44814981_49011000,
        64'h0ab7504c_b74d009b,
        64'h202300f4_02a30017,
        64'he793c804_00544783,
        64'hfef963e3_29054c1c,
        64'h2485e111_09550863,
        64'h09350863_2501a55f,
        64'he0ef8522_85ca4a85,
        64'h59fd4481_490902fb,
        64'h9f634785_00044b83,
        64'h80826165_6ce27c02,
        64'h7ba27b42_7ae26a06,
        64'h69a66946_64e68552,
        64'h740670a6_00fb2023,
        64'h02f76263_ffec871b,
        64'h481c0184_2c836000,
        64'h000a1c63_00050a1b,
        64'he7cfe0ef_ec66f062,
        64'hf45efc56_e4cee8ca,
        64'heca6f486_e0d28522,
        64'h002c4601_8b2ee42a,
        64'hf85a8432_f0a27159,
        64'hbfcd4419_80826165,
        64'h64e67406_70a68522,
        64'hc10fe0ef_102885a6,
        64'hc489cf81_6786e801,
        64'h0005041b_872ff0ef,
        64'he4be1028_083c65a2,
        64'he00d0005_041bedaf,
        64'he0eff486_f0a21028,
        64'h002c4601_84aee42a,
        64'heca67159_bf6584aa,
        64'hd16dbf7d_00042a23,
        64'h00f51663_47912501,
        64'hf8bfe0ef_85224581,
        64'hc68fe0ef_852285ca,
        64'h00042a23_02f51363,
        64'h47912501_b32ff0ef,
        64'h85224581_02243023,
        64'h80826145_64e26942,
        64'h85267402_70a20005,
        64'h049bc5ff_e0ef8522,
        64'h45810009_1f63e889,
        64'h0005049b_d98fe0ef,
        64'h892e842a_f406e84a,
        64'hec26f022_71798082,
        64'h01416402_60a20004,
        64'h3023e119_2501dbaf,
        64'he0ef842a_e406e022,
        64'h1141b7c1_fcf501e3,
        64'h4791bfdd_45258082,
        64'h61217442_70e2f971,
        64'hfcf50be3_47912501,
        64'hcbdfe0ef_00f41423,
        64'h0067d783_85224581,
        64'h67e2c448_e30fe0ef,
        64'h0007c503_67e2a02d,
        64'h00043023_4515e789,
        64'h8bc100b5_c783cd99,
        64'h6c0ce529_250197cf,
        64'hf0eff01c_101ce01c,
        64'h852265a2_67e2e115,
        64'h2501fe6f_e0ef0828,
        64'h002c4601_842ac52d,
        64'he42ef822_fc067139,
        64'hb7bdc45c_013787bb,
        64'h413484bb_cc0c445c,
        64'hfaf5fae3_4f9c601c,
        64'hfabafee3_fd4588e3,
        64'h0005059b_c4bfe0ef,
        64'hbf6984ce_e5990005,
        64'h059bfddf_e0efcb81,
        64'h8b896008_00a44783,
        64'hb765cc0c_c84cb5ed,
        64'h490500f4_05a34785,
        64'h00f59763_57fdbded,
        64'h490900f4_05a34789,
        64'h00f59763_47850005,
        64'h059b814f_f0efe595,
        64'h484cbfb1_9ca90094,
        64'hd49bcd11_2501c87f,
        64'he0ef6008_d7b51ff4,
        64'hf793c45c_9fa5445c,
        64'h0499ea63_4a855a7d,
        64'hd1c19c9d_c45c2781,
        64'h4c0c8ff9_413007bb,
        64'h02c6ed63_0337563b,
        64'h0336d6bb_fff4869b,
        64'h377dc729_0097999b,
        64'h00254783_6008bf59,
        64'hcc44ed35_25012190,
        64'h40ef85ce_0017c503,
        64'h86264685_601c00f4,
        64'h0523fbf7_f79300a4,
        64'h4783ed51_250126b0,
        64'h40ef0017_c50385ce,
        64'h4685601c_c3850407,
        64'hf7930304_099300a4,
        64'h4783fc96_0ee34c50,
        64'hd3e51ff7_f793445c,
        64'h4481bf7d_00f40523,
        64'h0207e793_00a44783,
        64'hc81cfcf7_78e34818,
        64'h445ce4bd_00042623,
        64'h445884ba_e3918b89,
        64'h00a44783_00977763,
        64'h48188082_61216aa2,
        64'h6a4269e2_790274a2,
        64'h854a7442_70e20007,
        64'h891bcf89_00b44783,
        64'h00091763_0005091b,
        64'hfb4fe0ef_84ae842a,
        64'he456e852_ec4efc06,
        64'hf04af426_f8227139,
        64'hb709fe94_65e3fee7,
        64'h8fa32405_07850007,
        64'h47039736_92810204,
        64'h16936722_0789bddd,
        64'h4545b7e9_00c68023,
        64'h377dfc96_4603962a,
        64'h10889201_02071613,
        64'hb7c12785_b7319c3d,
        64'h01368023_fff7c793,
        64'h01271a63_96b29201,
        64'h66a20206_961300e5,
        64'h86bb40f4_05bbfff7,
        64'h871b04e4_62630037,
        64'h871beb05_fc974703,
        64'h97361094_93010207,
        64'h97134781_f5cfe0ef,
        64'h1828100c_b7594509,
        64'hf8e516e3_67a24711,
        64'hdd612501_a9eff0ef,
        64'h18284581_01450e63,
        64'h25018a7f_e0ef0007,
        64'hc50365c6_77e2e105,
        64'h2501e48f_f0ef1828,
        64'h4581f949_2501f63f,
        64'he0ef1828_4581c2aa,
        64'h8cdfe0ef_0007c503,
        64'h65c677e2_f5552501,
        64'he6eff0ef_18284581,
        64'hfd452501_f89fe0ef,
        64'h18284585_80826149,
        64'h7a0679a6_794674e6,
        64'h640a60aa_00078023,
        64'h078d00e7_812302f0,
        64'h07130e94_186300e7,
        64'h80a303a0_071300e7,
        64'h80230307_071b14e7,
        64'h47030000_8717e505,
        64'h67a24501_040a1263,
        64'h4a16c2be_02f00993,
        64'h4bdc597d_842677e2,
        64'hecbe081c_e5292501,
        64'hacdfe0ef_1828002c,
        64'h460184ae_00050023,
        64'hf0d2f4ce_f8cae122,
        64'he506e42a_fca67175,
        64'hbfd94415_fcf41ee3,
        64'h4791b7c5_c8c897bf,
        64'he0ef0004_c50374a2,
        64'hcb998bc1_00b5c783,
        64'h80826165_64e67406,
        64'h70a68522_cbd85752,
        64'h77a2e991_6586e41d,
        64'h0005041b_cd2ff0ef,
        64'he4be1028_083c65a2,
        64'hec190005_041bb3bf,
        64'he0efeca6_f486f0a2,
        64'h1028002c_4601e42a,
        64'h7159bfe5_452d8082,
        64'h610560e2_450120a7,
        64'h83230000_87970005,
        64'h4a6395bf_e0efec06,
        64'h0028e42a_11018082,
        64'h01416402_60a20004,
        64'h3023e119_25019cbf,
        64'he0ef8522_e9012501,
        64'heffff0ef_842ae406,
        64'he0221141_80820141,
        64'h640260a2_4505ebbf,
        64'he06f0141_60a26402,
        64'h00f50223_478500f4,
        64'h0523fdf7_f7936008,
        64'h00a44783_000789a3,
        64'h00078923_00e78ca3,
        64'h00d78da3_04600713,
        64'h0086d69b_00e78c23,
        64'h02100713_0106d69b,
        64'h00e78aa3_0087571b,
        64'h0107571b_0107171b,
        64'h00e78a23_27010107,
        64'h571b0107_169b00e7,
        64'h8d230007_8ba30007,
        64'h8b234858_00e78fa3,
        64'h00d78f23_0187571b,
        64'h0107569b_00d78ea3,
        64'h00e78e23_0086d69b,
        64'h0106d69b_0107169b,
        64'h481800e7_85a30207,
        64'h671300b7_c703741c,
        64'he15d2501_b77fe0ef,
        64'h6008500c_00f40523,
        64'hfbf7f793_00a44783,
        64'hed552501_5e1040ef,
        64'h03040593_0017c503,
        64'h46854c50_601cc395,
        64'h0407f793_cf690207,
        64'hf71300a4_4783e175,
        64'h2501acff_e0ef842a,
        64'he406e022_1141bd2d,
        64'h499db5f9_c81cbf41,
        64'h00f40523_0407e793,
        64'h00a44783_9dbfe0ef,
        64'h952285d2_86260305,
        64'h05130007_849b0127,
        64'hf46340ab_87bb1ff5,
        64'h75130009_049b4448,
        64'h01a42e23_fd092501,
        64'h623040ef_85da4685,
        64'h001dc503_00e7fa63,
        64'h445c4818_00c78e63,
        64'h4c5cbdd1_00faa023,
        64'h9fa5000a_a783c45c,
        64'h9fa54099_093b445c,
        64'h9a3e9381_02049793,
        64'h0094949b_00f40523,
        64'hfbf7f793_00a44783,
        64'ha4ffe0ef_855a95d2,
        64'h20000613_91811582,
        64'h0097959b_0297f263,
        64'h41a587bb_4c4cf151,
        64'h25016bf0_40ef85d2,
        64'h86a6001d_c5034197,
        64'h04bb00f7_74639fb5,
        64'h002dc703_c4b58d32,
        64'h0007849b_00a6863b,
        64'h0099579b_000c869b,
        64'hd1592501_97cff0ef,
        64'h856e4c0c_00043d83,
        64'h00f40523_fbf7f793,
        64'h00a44783_f9692501,
        64'h70d040ef_85da0017,
        64'hc5034685_4c50601c,
        64'hc38d0407_f79300a4,
        64'h4783c85c_e311cc1c,
        64'h4858bf99_498500f4,
        64'h05a34785_01879763,
        64'hb79500f4_05230207,
        64'he79300a4_478312f7,
        64'h6a634818_445cf3fd,
        64'h0005079b_d86ff0ef,
        64'h4c0cb759_498900f4,
        64'h05a34789_02e79863,
        64'h4705cb91_4581485c,
        64'hef01040c_9a630ffc,
        64'hfc930197_fcb337fd,
        64'h00254783_00975c9b,
        64'h60081407_93631ff7,
        64'h77930409_04634458,
        64'h5c7d0304_0b132000,
        64'h0b9304f7_6c630127,
        64'h873b445c_18078f63,
        64'h8b8900a4_47838082,
        64'h61656da2_6d426ce2,
        64'h7c027ba2_7b427ae2,
        64'h6a0669a6_694664e6,
        64'h854e7406_70a60007,
        64'h899bc39d_00b44783,
        64'h00099763_0005099b,
        64'hcb5fe0ef_8ab68932,
        64'h8a2e842a_0006a023,
        64'he46ee86a_ec66f062,
        64'hf45ef85a_eca6f486,
        64'hfc56e0d2_e4cee8ca,
        64'hf0a27159_b59d499d,
        64'hbf9dbd1f_e0ef8552,
        64'h95a28626_03058593,
        64'h0007849b_0127f463,
        64'h40bb87bb_1ff5f593,
        64'h0009049b_444c01a4,
        64'h2e23f115_25010180,
        64'h50ef85da_0017c503,
        64'h863a4685_601c00f4,
        64'h0523fbf7_f7936722,
        64'h00a44783_f1392501,
        64'h06c050ef_e43a85da,
        64'h4685001d_c503c38d,
        64'h0407f793_00a44783,
        64'h04e60163_4c50b705,
        64'h00faa023_9fa5000a,
        64'ha783c45c_9fa54099,
        64'h093b445c_9a3e9381,
        64'h02049793_0094949b,
        64'hc5ffe0ef_955285da,
        64'h20000613_91011502,
        64'h0097951b_0097fc63,
        64'h41a507bb_4c48c385,
        64'h0407f793_00a44783,
        64'hf94d2501_0a6050ef,
        64'h85d2863a_86a6001d,
        64'hc5034196_84bb00f6,
        64'hf4639fb1_002dc683,
        64'hc4b58d3a_0007849b,
        64'h00a6073b_0099579b,
        64'h000c861b_d5792501,
        64'hb98ff0ef_856e4c0c,
        64'h00043d83_cc08b7a5,
        64'h498500f4_05a34785,
        64'h01851763_b7e52501,
        64'hbd6ff0ef_4c0cb741,
        64'h498900f4_05a34789,
        64'h00a7ec63_47854848,
        64'heb11020c_99630ffc,
        64'hfc930197_fcb337fd,
        64'h00254783_00975c9b,
        64'h60081207_90631ff7,
        64'h77934458_fa090ce3,
        64'h5c7d0304_0b132000,
        64'h0b930006_091b00f6,
        64'h7463893e_40f907bb,
        64'h445c0104_29031607,
        64'h89638b85_00a44783,
        64'h80826109_6de27d02,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e67906,
        64'h74a6854e_744670e6,
        64'h0007899b_c39d6622,
        64'h00b44783_00099863,
        64'h0005099b_e91fe0ef,
        64'h8ab6e432_8a2e842a,
        64'h0006a023_ec6ef06a,
        64'hf466f862_fc5ee0da,
        64'hf0caf4a6_fc86e4d6,
        64'he8d2ecce_f8a27119,
        64'hb7d5491d_b7e54911,
        64'h80826149_6b466ae6,
        64'h7a0679a6_794674e6,
        64'h854a640a_60aa00f4,
        64'h94230134_b0230004,
        64'hae230004_a623c888,
        64'h0069d783_dbbfe0ef,
        64'h01c40513_c8c8f33f,
        64'he0ef0009_c5030004,
        64'h85a3d09c_01448523,
        64'hf4800309_a78385a2,
        64'h79a2020a_6a13c399,
        64'h008a7793_e3ad8b85,
        64'h00098463_0029f993,
        64'he72d0107_f71300b4,
        64'h4783f565_a0854921,
        64'hf60981e3_0049f993,
        64'he3d98bc5_00b44783,
        64'ha895892a_c90d2501,
        64'h83aff0ef_01352623,
        64'h85da39fd_7522e911,
        64'h2501e3ff_f0ef030a,
        64'hab038556_85ce0409,
        64'h8b6300fa_82230005,
        64'h099b0004_0aa30004,
        64'h0a230004_0da30004,
        64'h0d234785_fc9fe0ef,
        64'h85a2000a_c5030004,
        64'h0fa30004_0f230004,
        64'h0ea30004_0e230004,
        64'h05a300e4_0c230004,
        64'h0ba30004_0b2300e4,
        64'h08230004_07a30004,
        64'h072300f4_0ca300f4,
        64'h08a30210_07130460,
        64'h07937aa2_cfcd008a,
        64'h77936406_e949008a,
        64'h6a132501_e75ff0ef,
        64'h102800f5_16634791,
        64'hc54dc3e1_01f9fa13,
        64'h01c9f793_4519e011,
        64'he1196406_2501b6df,
        64'hf0efe4be_1028083c,
        64'h65a21409_10630005,
        64'h091b9d6f_f0ef1028,
        64'h002c8a79_84aa89b2,
        64'h00053023_14050d63,
        64'h4925e42e_e8daecd6,
        64'hf0d2f4ce_fca6e122,
        64'he506f8ca_7175bfe5,
        64'h452d8082_612170e2,
        64'h2501a0ef_f0ef0828,
        64'h080c4601_00f61863,
        64'h4785cb11_4501e398,
        64'h97aa0007_0023c319,
        64'h67620007_0023c319,
        64'h66226318_00a78733,
        64'h050e8da7_87930000,
        64'h97970405_426383ef,
        64'hf0eff42e_e432e82e,
        64'hfc061028_ec2a7139,
        64'hb7594505_bf5d0009,
        64'h049b00f4_02a30017,
        64'he7930054_4783c81c,
        64'h27850137_8a63481c,
        64'hf15d2501_8afff0ef,
        64'h852285a6_46010339,
        64'h0763fb49_0ce3bf75,
        64'h45010009_14630005,
        64'h091bec8f_f0ef8522,
        64'h85a600f4_fa634c1c,
        64'h59fd4a05_fcf5fde3,
        64'h84ae842a_e052e44e,
        64'he84af406_ec26f022,
        64'h71794d1c_80826145,
        64'h6a0269a2_694264e2,
        64'h740270a2_45098082,
        64'h450900b7_ed634785,
        64'h80826105_64a28526,
        64'h644260e2_00e78223,
        64'h4705601c_82aff0ef,
        64'h462d6c08_700c84cf,
        64'hf0ef4581_02000613,
        64'h6c08e085_0005049b,
        64'ha42ff0ef_6008484c,
        64'he49d0005_049bfa9f,
        64'hf0ef842a_ec06e426,
        64'he8221101_80826105,
        64'h64a26442_60e2451d,
        64'h00f51363_4791dd79,
        64'h2501bcdf_f0ef8522,
        64'h4585cb99_00978d63,
        64'h0007c783_6c1ced09,
        64'h2501a8cf_f0ef6008,
        64'h484c0e50_0493e50d,
        64'h250188ff_f0ef842a,
        64'he426ec06_e8224581,
        64'h1101bfe5_4511b7cd,
        64'h00042a23_d9452501,
        64'hc13ff0ef_85224581,
        64'h80826145_69a26942,
        64'h64e27402_70a24501,
        64'h00979a63_0017b793,
        64'h17e18bfd_03378063,
        64'h03270263_03f7f793,
        64'h00b7c783_c3210007,
        64'hc7036c1c_e1292501,
        64'hafaff0ef_6008a0b1,
        64'hc90de199_484c49bd,
        64'h0e500913_451184ae,
        64'hf406842a_e44ee84a,
        64'hec26f022_7179bdf9,
        64'h0ff77713_0017e793,
        64'h3701eea8_66e30ff5,
        64'h7513f9f7_051beea8,
        64'h7ae30ff5_7513fbf7,
        64'h051bbd6d_4519f117,
        64'h10e30008_86630005,
        64'h4883cfa5_05130000,
        64'h85170005_4c634185,
        64'h551b0187_151b02b6,
        64'hf263fd37_0ae3f957,
        64'h04e3f947_06e3f4e3,
        64'h74e30007_47039722,
        64'h93011702_0017061b,
        64'h873245ad_46a10ff7,
        64'hf7930027_979b0565,
        64'h9a63bdb9_c4c8af2f,
        64'hf0ef0007_c503609c,
        64'hdbe58bc1_00b5c783,
        64'h6c8cfbf5_8b91b73d,
        64'h4515fb0d_bf154501,
        64'he80703e3_0004bc23,
        64'h0004a623_cb890207,
        64'hf7930047_f713f4e5,
        64'h18e34711_c50500b7,
        64'hc783709c_4511bf65,
        64'h4701bdfd_00e905a3,
        64'h94329201_16020087,
        64'h671300d7_94634691,
        64'h8bb10107_671300b6,
        64'h94634585_0037f693,
        64'h0ff7f793_0027979b,
        64'h01659663_00d90023,
        64'h469500d5_15630e50,
        64'h06930009_4503c6ed,
        64'h4711a06d_268500e5,
        64'h0023954a_91010206,
        64'h95130027_e793a8dd,
        64'h0505a0d1_48650200,
        64'h03134781_45a14701,
        64'h4681b7ad_02400793,
        64'h943a12f6_e0630200,
        64'h0693f757_8be3bf95,
        64'h4709bf1d_04058082,
        64'h61216b02_6aa26a42,
        64'h69e27902_74a27442,
        64'h70e20004_bc232501,
        64'ha85ff0ef_85264581,
        64'hb791c55c_4bdc611c,
        64'hbf75dfdf_f0ef8526,
        64'h4581fed6_08e3fff7,
        64'hc683fff7_46030785,
        64'h07050cb7_8d6300b7,
        64'h8593709c_ef918ba1,
        64'h00b74783_c7e50007,
        64'h47836c98_e96d2501,
        64'hcdaff0ef_608848cc,
        64'h10051063_2501adbf,
        64'hf0ef8526_458100f9,
        64'h05a30200_0793943a,
        64'h09479763_470d1b37,
        64'h8e630024_478300f9,
        64'h00a302e0_07930b37,
        64'h90630014_47830139,
        64'h00230d37_92630004,
        64'h4783b40f_f0ef854a,
        64'h02000593_462d0204,
        64'hb9030d57_80630d47,
        64'h82630004_47834b21,
        64'h02e00993_05c00a93,
        64'h02f00a13_0ae7fc63,
        64'h47fd0004_47030004,
        64'ha6230405_0ce79063,
        64'h05c00713_00e78663,
        64'h842e84aa_02f00713,
        64'h0005c783_e05ae456,
        64'he852ec4e_f04afc06,
        64'hf426f822_7139b7e9,
        64'hdb1c2785_5b1c2a85,
        64'h6018f141_2501d1cf,
        64'hf0ef0145_0223b7b9,
        64'hc848a83f_f0ef85a6,
        64'hc8046008_d91c4157,
        64'h87bb591c_00faed63,
        64'h00254783_60084a05,
        64'h02aa2823_aa5ff0ef,
        64'h855285a6_00043a03,
        64'hbeeff0ef_03450513,
        64'h45812000_06136008,
        64'hf5792501_dd8ff0ef,
        64'h6008fcf4_8de357fd,
        64'hfcf48be3_4785d4bd,
        64'h451d0005_049be81f,
        64'hf0ef480c_f60a0ee3,
        64'h06f4e063_4d1c6008,
        64'hb7614505_00f49463,
        64'h57fdbf49_45090097,
        64'he4634785_0005049b,
        64'hb27ff0ef_fc0a9fe3,
        64'h0157fab3_37fd0049,
        64'h5a9b0025_4783bf5d,
        64'h4501ec1c_97ce0347,
        64'h87930124_15230996,
        64'h601cfcf7_75e30009,
        64'h071b0085_5783e18d,
        64'hc85c6108_2785480c,
        64'h00099d63_842a8a2e,
        64'h00f97993_d7ed495c,
        64'h80826121_6aa26a42,
        64'h69e27902_74a27442,
        64'h70e24511_eb9993c1,
        64'he456e852_ec4ef426,
        64'h03091793_2905f822,
        64'hfc0600a5_5903f04a,
        64'h7139bfad_4405f6f5,
        64'h0fe34785_dd612501,
        64'hdbbff0ef_852685ce,
        64'h8622bf49_00f482a3,
        64'h0017e793_0054c783,
        64'hc89c37fd_fae783e3,
        64'h577dc4c0_489c0209,
        64'h9063e905_2501de9f,
        64'hf0ef8526_85a2167d,
        64'h10000637_b76dfb24,
        64'h11e30545_0863fd55,
        64'h07e3c901_2501c05f,
        64'hf0ef8526_85a24409,
        64'hbf554905_b7d5faf4,
        64'h7ee3894e_4c9c8082,
        64'h61216aa2_6a4269e2,
        64'h790274a2_744270e2,
        64'h8522547d_00f41d63,
        64'h57fd0887_f8634785,
        64'h0005041b_c43ff0ef,
        64'ha8214401_052a6063,
        64'h04f46363_24054c9c,
        64'h5afd4a05_844a04f9,
        64'h77634d1c_04090a63,
        64'h00c52903_e19d89ae,
        64'h84aae456_e852f04a,
        64'hf822fc06_ec4ef426,
        64'h7139bf3d_4989b745,
        64'h012a81a3_00fa8123,
        64'h0189591b_0109579b,
        64'h00fa80a3_0087d79b,
        64'h03240a23_0107d79b,
        64'h94260109_179b0125,
        64'h69338d71_f0000637,
        64'h2501da0f_f0ef8556,
        64'h9aa60344_0a931fc4,
        64'h74130024_141bf809,
        64'h96e30005_099bfd8f,
        64'hf0ef9dbd_0075d59b,
        64'h515cbf79_01448223,
        64'h03240aa3_0089591b,
        64'h0109591b_0109191b,
        64'h03240a23_94261fe4,
        64'h74130014_141bfc09,
        64'h92e30005_099b811f,
        64'hf0ef9dbd_0085d59b,
        64'h515cb7e9_0127e933,
        64'h9bc100f9_79130089,
        64'h591b0347_c7830154,
        64'h87b38082_61216aa2,
        64'h6a4269e2_790274a2,
        64'h854e7442_70e200f4,
        64'h82234785_032a8a23,
        64'h9aa60ff9_79130049,
        64'h591bc40d_1ffafa93,
        64'h00099f63_0005099b,
        64'h86bff0ef_9dbd8526,
        64'h009ad59b_50dc00f4,
        64'h82234785_02fa0a23,
        64'h9a260ff7_f7938fd9,
        64'h8ff50049_179b00f7,
        64'hf71316c1_66850347,
        64'hc7830144_87b3cc19,
        64'h1ffa7a13_0ff97793,
        64'h001a0a9b_88050609,
        64'h96630005_099b8b9f,
        64'hf0ef9dbd_009a559b,
        64'h00ba0a3b_515c0015,
        64'hda1b1547_94630ee7,
        64'h8863470d_0ae78f63,
        64'h842e8932_47090005,
        64'h47830af5_f0634989,
        64'h84aa4d1c_16ba7563,
        64'h4a05e456_ec4ef04a,
        64'hf426f822_fc06e852,
        64'h71398082_610564a2,
        64'h85266442_60e200e7,
        64'h82234705_601c00e7,
        64'h80235715_6c1cf3cf,
        64'hf0ef4581_02000613,
        64'h6c08ec99_0005049b,
        64'h933ff0ef_6008484c,
        64'he4950005_049bf33f,
        64'hf0ef842a_ec06e426,
        64'he8221101_00a55583,
        64'hb78d4505_bfc14134,
        64'h84bbf6f4_76e34f9c,
        64'h00093783_f68afbe3,
        64'h01440c63_0005041b,
        64'he6fff0ef_bf752501,
        64'he59ff0ef_0134f663,
        64'h85a20009_35034a85,
        64'h09925a7d_843a0027,
        64'hc9838722_b75d4501,
        64'h00993c23_00a92a23,
        64'h94be0347_87930496,
        64'h88bd0009_37839d3d,
        64'h0044d79b_d1710089,
        64'h28235788_fce4f7e3,
        64'h0087d703_eb155798,
        64'h00e69463_470d0007,
        64'hc683e021_84aefee4,
        64'h74e34f98_611c8082,
        64'h61216aa2_6a4269e2,
        64'h790274a2_744270e2,
        64'h450900f4_1c63892a,
        64'h478500b5_1523e456,
        64'he852ec4e_f426fc06,
        64'hf04a4540_f8227139,
        64'h8082853e_4785b765,
        64'h17fd2501_100007b7,
        64'h807ff0ef_954a0345,
        64'h05131fc5_75130024,
        64'h151bf935_2501a39f,
        64'hf0ef9dbd_0075d59b,
        64'h515cb759_8fc90087,
        64'h979b0349_45030359,
        64'h47839922_1fe47413,
        64'h0014141b_fd592501,
        64'ha63ff0ef_9dbd0085,
        64'hd59b515c_bf458fe9,
        64'h157d6505_bf658391,
        64'hc0198fc5_0087979b,
        64'h88050349_4783994e,
        64'h1ff9f993_f5792501,
        64'ha93ff0ef_0344c483,
        64'h854a9dbd_94ca1ff4,
        64'hf4930099_d59b0014,
        64'h899b0249_27838082,
        64'h6145853e_69a26942,
        64'h64e27402_70a257fd,
        64'hc9112501_ac7ff0ef,
        64'h9dbd0094_d59b9cad,
        64'h515c0015_d49b00f7,
        64'h1e6308d7_0e63468d,
        64'h06d70c63_842e4689,
        64'h00054703_02e5f963,
        64'h892ae44e_ec26f022,
        64'hf406e84a_71794d18,
        64'h0eb7f763_47858082,
        64'h45018082_9d2d02d5,
        64'h85bb5548_00254583,
        64'h00f6f963_37f9ffe5,
        64'h869b4d1c_80826105,
        64'h64a26442_60e200a0,
        64'h35332501_58d050ef,
        64'h45814601_00144503,
        64'h000402a3_599050ef,
        64'h85a64685_d81022f4,
        64'h01a322e4_012320d4,
        64'h0ca320d4_0c230187,
        64'hd79b0107_d71b2605,
        64'h22e400a3_22f40023,
        64'h07200693_00144503,
        64'h0087571b_0107571b,
        64'h0107971b_501020e4,
        64'h0f23445c_20f40fa3,
        64'h0187d79b_0107d71b,
        64'h20e40ea3_20f40e23,
        64'h0087571b_0107571b,
        64'h0107971b_20e40d23,
        64'h02e40ba3_04100713,
        64'h481c20f4_0da302f4,
        64'h0b230610_079302f4,
        64'h0aa302f4_0a230520,
        64'h079322f4_09a3faa0,
        64'h079322f4_09230550,
        64'h0793a01f_f0ef8526,
        64'h45812000_06130344,
        64'h04930af7_1b634785,
        64'h00544703_0cf71063,
        64'h478d0004_4703ed69,
        64'h2501bfff_f0ef842a,
        64'he426ec06_e8221101,
        64'hbdc59cbd_0017d79b,
        64'h88850297_87bb478d,
        64'hb7010014_949b00f9,
        64'h15634789_d41c9fb5,
        64'he00a05e3_b545a25f,
        64'hf0ef0544_0513b5b9,
        64'h0005099b_a33ff0ef,
        64'h05840513_b3514781,
        64'h00042a23_01240023,
        64'h00f41323_3ef71323,
        64'h00009717_93c117c2,
        64'h27853f47_d7830000,
        64'h9797c448_a63ff0ef,
        64'h22040513_c808a6df,
        64'hf0ef21c4_051300f5,
        64'h1c632727_87932501,
        64'h614177b7_a83ff0ef,
        64'h21840513_02f51763,
        64'h25278793_25014161,
        64'h57b7a99f_f0ef0344,
        64'h051304f7_1263a557,
        64'h07134107_d79b776d,
        64'h0107979b_8fd90087,
        64'h979b0004_02a32324,
        64'h47032334_4783e13d,
        64'h2501ce5f_f0ef8522,
        64'h001a859b_06f71b63,
        64'h47054107_d79b0107,
        64'h979b8fd9_0087979b,
        64'h06444703_06544783,
        64'h08f91963_478d00f4,
        64'h02a3f800_0793c45c,
        64'hc81c57fd_ee99e7e3,
        64'h24810094_d49b1ff4,
        64'h849b0024_949bd408,
        64'hb17ff0ef_06040513,
        64'hf00a15e3_10e91263,
        64'h470dd05c_03542023,
        64'hcc04d458_015787bb,
        64'h248900ea_873b490d,
        64'h00b67363_09051655,
        64'h00b93933_66411955,
        64'h6905dd8d_84ae0364,
        64'hd5bb40c5_04bbf4c5,
        64'h64e38732_00d7063b,
        64'h9f3d004a_571b2781,
        64'h033906bb_dfb18fd9,
        64'h0087979b_25010424,
        64'h47030434_47831405,
        64'h0e638d45_0085151b,
        64'h04744483_04844503,
        64'hf3c100fa_77930144,
        64'h142300fa_6a33008a,
        64'h1a1b0454_47830464,
        64'h4a03ffc9_00fb77b3,
        64'hfffb079b_fa0b03e3,
        64'h01640123_04144b03,
        64'hfaf769e3_0ff7f793,
        64'h012401a3_fff9079b,
        64'h47050134_2e230444,
        64'h49032981_1a098663,
        64'h00f9e9b3_0089999b,
        64'h04a44783_04b44983,
        64'hfef711e3_20000713,
        64'h4107d79b_0107979b,
        64'h8fd90087_979b03f4,
        64'h47030404_4783bfb9,
        64'h47b5c119_4a81f6e5,
        64'h04e34785_470db7bd,
        64'h00e51963_4785470d,
        64'hfe9915e3_0491c10d,
        64'he9dff0ef_852285d6,
        64'h000a8763_45090004,
        64'haa830104_8913ff2a,
        64'h14e30991_094100a9,
        64'ha0232501_c5bff0ef,
        64'h854ac789_4501ffc9,
        64'h478389a6_23a40a13,
        64'h1fa40913_848a04f5,
        64'h1a634785_ee1ff0ef,
        64'h85224581_f5698911,
        64'h00090463_fb71478d,
        64'h00157713_050060ef,
        64'h00a400a3_00040023,
        64'h0ff4f513_80826161,
        64'h853e6b42_6ae27a02,
        64'h79a27942_74e26406,
        64'h60a647a9_c1118911,
        64'h00090563_e38d0015,
        64'h779313e0_60ef0014,
        64'h4503cb85_00044783,
        64'h0089b023_c01547b1,
        64'h84aa6380_97ba66e7,
        64'h87930000_97970035,
        64'h17130205_4e6347ad,
        64'hdd9ff0ef_8932852e,
        64'h89aa0005_3023e85a,
        64'hec56f052_fc26e0a2,
        64'he486f44e_f84a715d,
        64'hbfcd450d_80826105,
        64'h690264a2_644260e2,
        64'h00a03533_8d050125,
        64'h75332501_d33ff0ef,
        64'h08640513_00978c63,
        64'h45010127_f7b31465,
        64'h04930054_4537fff5,
        64'h09130100_05370005,
        64'h079bd59f_f0ef06a4,
        64'h051302f7_1f63a557,
        64'h07134107_d79b776d,
        64'h0107979b_8fd90087,
        64'h979b4509_23244703,
        64'h23344783_e52d2501,
        64'hfa3ff0ef_842ad91c,
        64'h00050223_57fde04a,
        64'he426ec06_e8221101,
        64'h80826105_690264a2,
        64'h644260e2_85220324,
        64'ha823597d_4405c119,
        64'h25011f40_60ef0344,
        64'h8593864a_46850014,
        64'hc503ec19_0005041b,
        64'hfddff0ef_892e84aa,
        64'h02b78763_4401e04a,
        64'he426ec06_e8221101,
        64'h591c8082_4501f8df,
        64'hf06fc399_00454783,
        64'hb7f94505_b7e5397d,
        64'h26c060ef_85ce8626,
        64'h9cbd4685_00144503,
        64'h4c5cff2a_74e34a05,
        64'h00344903_80826145,
        64'h6a0269a2_694264e2,
        64'h740270a2_450100e7,
        64'heb6340f4_87bb0004,
        64'h02234c58_505ce131,
        64'h25012ae0_60ef85ce,
        64'h86264685_00154503,
        64'h842a0345_0993e052,
        64'he84af406_5904e44e,
        64'hec26f022_71798082,
        64'h853e2781_8fd90107,
        64'h979b8fd5_0087979b,
        64'h0145c683_0155c783,
        64'h00d51d63_0007079b,
        64'h8f5d0087_979b468d,
        64'h01a5c703_01b5c783,
        64'h80824525_80820141,
        64'h60a24525_c3914501,
        64'h00157793_320060ef,
        64'h0017c503_e4061141,
        64'h02e69063_00855703,
        64'h0067d683_c70d0007,
        64'hc703cb85_611cc915,
        64'hbfd586a7_47030000,
        64'ha7178082_853ae11c,
        64'h0006871b_078900b6,
        64'h66630ff6_f593fd06,
        64'h869b577d_46050007,
        64'hc683b7dd_0705a00d,
        64'h577d00d7_06630017,
        64'h869300c6_986302d5,
        64'hfc630007_468303a0,
        64'h06130200_0593cf99,
        64'h873e611c_80826105,
        64'h690264a2_644260e2,
        64'h00040023_00f49323,
        64'h8fd90087_979b0169,
        64'h47030179_478300f4,
        64'h92238fd9_0087979b,
        64'h01894703_01994783,
        64'hc088f59f_f0ef00f5,
        64'h842384ae_01c90513,
        64'h00b94783_fcc79ee3,
        64'h06850405_00e40023,
        64'h04050064_00230117,
        64'h95630e50_07130107,
        64'h146300a7_0e632785,
        64'h0006c703_462d02e0,
        64'h031348a5_481586ca,
        64'h02000513_47810185,
        64'h3903cfa5_00958413,
        64'he04ae426_ec06e822,
        64'h1101495c_bfcd0505,
        64'h00b50023_808200f6,
        64'h1363367d_57fdb7f5,
        64'hfee50fa3_05850505,
        64'h0005c703_808200f6,
        64'h1363367d_57fd8082,
        64'h25018d5d_05628fd9,
        64'h07c20035_45030025,
        64'h47838f5d_07a20005,
        64'h47030015_47838082,
        64'h014160a2_30200073,
        64'h0ff0000f_0000100f,
        64'h7ac030ef_bc450513,
        64'h00009517_34179073,
        64'h07fe4785_30079073,
        64'h8fd98807_07136709,
        64'h300027f3_7d0030ef,
        64'hbc850513_00009517,
        64'h7dc030ef_bac50513,
        64'h00009517_8307b583,
        64'h82e7b823_f0070713,
        64'h670580e7_b4238f75,
        64'he40616fd_1141ff80,
        64'h06b78087_b7033000,
        64'h17b7b7d9_14fdb7e9,
        64'hc35ff0ef_bfc1710a,
        64'h84937bf0_50ef4501,
        64'hdff154fd_000a2783,
        64'hbfc5c4ff_f0effc07,
        64'h5de30337_97138309,
        64'h37830207_45630337,
        64'h97138309_3783680b,
        64'h0493f4bf_e0ef8522,
        64'he78d0009_a783e4a9,
        64'ha007ac23_0000a797,
        64'ha207a223_0000a797,
        64'ha207a823_0000a797,
        64'ha207a423_0000a797,
        64'ha2079a23_0000a797,
        64'ha4f70ea3_0000a717,
        64'h00544783_a6f70423,
        64'h0000a717_00444783,
        64'ha6f709a3_0000a717,
        64'h00344783_a6f70f23,
        64'h0000a717_00244783,
        64'ha8f704a3_0000a717,
        64'h30001937_00144783,
        64'ha8f70c23_0000a717,
        64'h00989b37_6a890004,
        64'h47830d70_30efc765,
        64'h05130000_9517aae5,
        64'hc5830000_a597ab76,
        64'h46030000_a617ac06,
        64'hc6830000_a697acb8,
        64'h48030000_a817ad27,
        64'hc7830000_a797ad97,
        64'h47030000_a7171130,
        64'h30ef80e7_b4238f4d,
        64'h91c115c2_adca0a13,
        64'h0000aa17_00800737,
        64'h8087b583_8007b603,
        64'h82e7b423_4721cc65,
        64'h05130000_95178087,
        64'hb7038007_b70380e7,
        64'hb4239341_80a7b023,
        64'h17429101_300017b7,
        64'h15028f55_8f710ff6,
        64'hf69382a1_0086971b,
        64'hf0060613_01000637,
        64'h46b2f4ff_f0efb2e9,
        64'h89930000_a9974481,
        64'h45227d80_50ef0068,
        64'h85a24609_7e2050ef,
        64'hb6f702a3_0000a717,
        64'hb6840413_0000a417,
        64'h0028b745_85930000,
        64'ha59707f0_07934611,
        64'hb8f70223_0000a717,
        64'h578db8f7_06a30000,
        64'ha7174789_b8f70b23,
        64'h0000a717_03e00793,
        64'hbaf700a3_0000a717,
        64'h47e1ba07_85230000,
        64'ha7971e70_30efe85a,
        64'hec56f052_f44ef84a,
        64'hfc26e0a2_e486d765,
        64'h05130000_9517715d,
        64'h80822501_8d5d8d79,
        64'h00ff0737_0085151b,
        64'h8fd98f75_0085571b,
        64'hf0068693_8fd966c1,
        64'h0185579b_0185171b,
        64'h80829141_15428d5d,
        64'h05220085_579b8082,
        64'h614564e2_740270a2,
        64'h85228aef_f0efc165,
        64'h05130000_a5170450,
        64'h0693c0e7_57030000,
        64'ha717c0a8_88930000,
        64'ha89785a6_862247b2,
        64'h0007a803_c2478793,
        64'h0000a797_0cb050ef,
        64'hf4060068_c6c58593,
        64'h0000a597_461184ae,
        64'h8432ec26_f0227179,
        64'hbfc14785_eb9ff0ef,
        64'h80826105_64a26442,
        64'h60e2c3c0_0c2007b7,
        64'h2ad030ef_e1450513,
        64'h00009517_e7990206,
        64'hc1630337_16938304,
        64'hb7033000_14b74781,
        64'h2401ec06_e42643c0,
        64'he8220c20_07b71101,
        64'hb7e1ff06_bc2306a1,
        64'h26050008_380300d7,
        64'h88338082_61010113,
        64'h5f813483_85266001,
        64'h34036081_30838287,
        64'hb8233000_17b70405,
        64'haa1ff0ef_862602e6,
        64'h446397c2_85b63000,
        64'h08378f95_868a83f5,
        64'h02d7473b_17822705,
        64'h46a10077_67139fad,
        64'h377d8005_859b6585,
        64'h02d51a63_80668693,
        64'h6685c691_8005069b,
        64'h00015503_00d10023,
        64'h0086d69b_0106d69b,
        64'h0106969b_00d100a3,
        64'h872646d4_96aa068e,
        64'h9ebd8006_869b7007,
        64'hf7930084_179bea25,
        64'h4390d427_87930000,
        64'ha797cfb5_27818ff1,
        64'hfff7c793_00c5963b,
        64'h10100593_8a1d08b8,
        64'h696335b9_5f200813,
        64'hffc5849b_25816011,
        64'h34235e91_3c23630c,
        64'h8387b783_972a3000,
        64'h05379f2d_8406871b,
        64'h03877593_66850034,
        64'h171b00f6_74132601,
        64'h60813023_9f010113,
        64'h8307b603_300017b7,
        64'hbba54601_3e9030ef,
        64'hf3850513_00009517,
        64'h85aab369_00f41623,
        64'h60800793_00f41f23,
        64'h0024d783_00f41e23,
        64'h0004d783_02f41423,
        64'h01e45783_02f41323,
        64'h02a00613_01c45783,
        64'h277050ef_852285ca,
        64'h46192810_50ef0064,
        64'h0513e0a5_85930000,
        64'ha5974619_293050ef,
        64'h854ee1a5_85930000,
        64'ha5974619_2a3050ef,
        64'h854a85ce_461900f5,
        64'h9a230165_89930205,
        64'h89132000_0793eaf7,
        64'h19e3e5c7_d7830000,
        64'ha7970285_d703ecf7,
        64'h11e3e6a4_84930000,
        64'ha497e727_d7830000,
        64'ha7970265_d703b1e1,
        64'hfb050513_00009517,
        64'hb9c9fa25_05130000,
        64'h9517b9f1_f7c50513,
        64'h00009517_b1ddf665,
        64'h05130000_9517b9c5,
        64'hf5850513_00009517,
        64'hb9edf3a5_05130000,
        64'h9517b311_f3450513,
        64'h00009517_b339f1e5,
        64'h05130000_9517bb21,
        64'hf1050513_00009517,
        64'hb30defa5_05130000,
        64'h9517b335_ef450513,
        64'h00009517_b7993550,
        64'h50ef0868_ef458593,
        64'h0000a597_4611f4f7,
        64'h0de30204_5703f6f7,
        64'h01e317fd_67c101e4,
        64'h5703f6e7_87e35fe0,
        64'h0713bf95_ca0ff0ef,
        64'h02a40513_85ca53b0,
        64'h30eff1a5_05130000,
        64'h9517cb6f_f0ef8522,
        64'h85a654f0_30eff1e5,
        64'h05130000_951702e7,
        64'h98634d20_0713b765,
        64'hd61fe0ef_02a40513,
        64'hf3858593_0000a597,
        64'hf3460613_0000a617,
        64'hf3868693_0000a697,
        64'hf7e9439c_f4478793,
        64'h0000a797_c799439c,
        64'hf5478793_0000a797,
        64'hf4f72823_0000a717,
        64'h47e204e6_94630430,
        64'h07138082_616179a2,
        64'h794274e2_640660a6,
        64'h508060ef_450102a4,
        64'h0593ff89_061bf667,
        64'h87930000_a79766a2,
        64'h47624290_50efe436,
        64'hf8f72823_0000a717,
        64'hf9050513_0000a517,
        64'hf8858593_0000a597,
        64'h461947e2_fad79823,
        64'h0000a797_04e79b63,
        64'h01c15683_04500713,
        64'h00e10e23_02344703,
        64'h00e10ea3_01c11903,
        64'h02244703_00e10e23,
        64'h27810274_470300e1,
        64'h0ea301c1_178300f1,
        64'h0e230254_478300f1,
        64'h0ea30264_47030244,
        64'h4783bdb5_00450513,
        64'h00009517_b559ff65,
        64'h05130000_9517bd41,
        64'hfe850513_00009517,
        64'ha06ddbff_e0ef4501,
        64'h85a202f4_12238626,
        64'h01c15783_00a10e23,
        64'h812100a1_0ea3db9f,
        64'hf0ef00f4_1e230029,
        64'hd78300f4_1d230009,
        64'hd78302f4_10230224,
        64'h0513fde4_859b01c4,
        64'h578300f4_1f230204,
        64'h12230204_012301a4,
        64'h57835090_50ef854a,
        64'h09058593_0000a597,
        64'h46195190_50ef8522,
        64'h85ca4619_10f71c63,
        64'h0c27d783_0000a797,
        64'h02045703_12f71463,
        64'h0d098993_0000a997,
        64'h0d87d783_0000a797,
        64'h01e45703_b73d1e65,
        64'h05130000_9517f0f5,
        64'h9ce30880_079326f5,
        64'h89630ff0_079326f5,
        64'h88630890_0793b73d,
        64'hf4f58ae3_1dc50513,
        64'h00009517_06c00793,
        64'h26f58b63_06700793,
        64'h00b7ef63_28f58663,
        64'h08400793_bf91f6f5,
        64'h8de31ca5_05130000,
        64'h951705e0_079328f5,
        64'h846305c0_0793b7bd,
        64'hf8f58ae3_1b450513,
        64'h00009517_03200793,
        64'h28f58763_02f00793,
        64'h00b7ef63_2af58263,
        64'h03300793_04b7e263,
        64'h2cf58263_06200793,
        64'hb7c91b25_05130000,
        64'h9517faf5_96e30290,
        64'h07932af5_86630210,
        64'h0793bf6d_fef580e3,
        64'h19850513_00009517,
        64'h47d916f5_8a6347c5,
        64'h00b7ed63_2cf58263,
        64'h47f5a431_7c9030ef,
        64'hfef591e3_17c50513,
        64'h00009517_47a118f5,
        64'h82634799_a41d7e30,
        64'h30ef3125_05130000,
        64'h951702f5_83631765,
        64'h05130000_95174789,
        64'h10f58463_478502b7,
        64'he3631af5_83634791,
        64'h04b7e563_1cf58263,
        64'h47b108b7_e76332f5,
        64'h896302e0_07930174,
        64'h45836790_50ef1c65,
        64'h05130000_a5174619,
        64'h85ca0064_091368d0,
        64'h50ef4611_082884b2,
        64'h05e94407_9a638005,
        64'h079b0af5_0e636dd7,
        64'h879367a1_3cf50563,
        64'h842e8067_8793f44e,
        64'hf84afc26_e486e0a2,
        64'h6785715d_bf55943e,
        64'h00e15783_00f10723,
        64'h00d14783_00f107a3,
        64'h34f90909_00c14783,
        64'h6df050ef_00684609,
        64'h85ca8082_61459141,
        64'h694264e2_1542fff5,
        64'h45137402_70a29522,
        64'h01045513_942a9041,
        64'h14420104_55130290,
        64'h44634401_84ae892a,
        64'hf406e84a_ec26f022,
        64'h71798082_1ec50513,
        64'h00009517_bf752365,
        64'h05130000_95178407,
        64'h8793fce6_08e32365,
        64'h05130000_95178387,
        64'h8713bfe9_22450513,
        64'h00009517_82878793,
        64'h00c74963_fee609e3,
        64'h24850513_00009517,
        64'h83078713_8082faf6,
        64'h12e322a5_05130000,
        64'h95178187_879300e6,
        64'h0a6322a5_05130000,
        64'h95178107_87138082,
        64'h01412c25_05130000,
        64'ha51760a2_124040ef,
        64'he4062d25_05130000,
        64'ha5172ca5_85930000,
        64'h95979e3d_11417c07,
        64'h879b77fd_04c7c963,
        64'h2d850513_00009517,
        64'h87f78793_6785c3ad,
        64'h25850513_00009517,
        64'h8006079b_04c74963,
        64'h06e60b63_27c50513,
        64'h00009517_80878713,
        64'h08a74463_862a0ce5,
        64'h07638207_87136785,
        64'h8082953e_057e4505,
        64'h97aa2000_0537e308,
        64'h95360017_86930075,
        64'h6513157d_631c36e7,
        64'h07130000_a7178082,
        64'h40000537_8082057e,
        64'h45058082_853e4785,
        64'hbf990384_04132a05,
        64'h7ed050ef_856a4581,
        64'h864e1f60_40ef8562,
        64'h85ea9d3e_864e40f9,
        64'h89b30184_3d030337,
        64'hf163701c_02843983,
        64'h066060ef_856a85ee,
        64'h864e21e0_40ef8566,
        64'h86ce85ea_866e8082,
        64'h6165853e_6da26d42,
        64'h6ce27c02_7ba27b42,
        64'h7ae26a06_69a66946,
        64'h64e67406_70a6478d,
        64'h24c040ef_2dc50513,
        64'h00009517_864a02ba,
        64'hfa6395ce_00b48db3,
        64'h01843d03_640c0409,
        64'h8d630204_39832720,
        64'h40ef855e_85d2cbc1,
        64'h741c0967_9b63401c,
        64'ha8354781_00fa6463,
        64'h0384d783_33cc8c93,
        64'h00009c97_35cc0c13,
        64'h00009c17_31cb8b93,
        64'h00009b97_4b054a01,
        64'h942a84aa_892e06ea,
        64'he663478d_9722020a,
        64'hda93e46e_e86aec66,
        64'hf062f45e_f85ae0d2,
        64'he4cee8ca_eca6f486,
        64'h02059a93_fc567100,
        64'hf0a202f7_07337159,
        64'h03800793_03855703,
        64'h10e69763_47090045,
        64'h468310e6_9c634789,
        64'h57f70713_464c4737,
        64'h00056683_12b7f463,
        64'h04000793_bfd58f8d,
        64'h25058082_e21c00b7,
        64'hf4634501_918187aa,
        64'h1582bf39_07050107,
        64'h00230005_d4634185,
        64'hd59b0185_959bc519,
        64'h09757513_00054503,
        64'h00bc0533_00074583,
        64'hbfdd4701_bf1d3cfd,
        64'hfe976ae3_27056722,
        64'h04e070ef_e43a855e,
        64'hb75d00c5_80230ff6,
        64'h761300ea_85b30006,
        64'hc603bf65_00c59023,
        64'h92411642_95d60017,
        64'h15930006_d603006d,
        64'h1c63bfc1_e19095d6,
        64'h00371593_6290011d,
        64'h1863bf85_68627882,
        64'h070596d2_73226742,
        64'h66a23ae0_40efe436,
        64'he83aec42_f046f41a,
        64'h855a6582_92011602,
        64'hc1902601_95d60027,
        64'h15934290_030d1b63,
        64'hb795557d_d1350220,
        64'h70ef9936_92811682,
        64'h41b4043b_66a23ea0,
        64'h40effa06_0c23e436,
        64'h46850513_00009517,
        64'h85d6963e_011c0ac5,
        64'hed634157_05bb0006,
        64'h861b02e0_08138756,
        64'h03bd06bb_0d9de663,
        64'h99ba0347_07339301,
        64'h020d9713_05b66c63,
        64'h0007061b_430948a1,
        64'h48114701_86ce000c,
        64'h8d9b008c_f4630004,
        64'h0d9b4460_40ef4ae5,
        64'h05130000_951785ca,
        64'h8082616d_6daa6d4a,
        64'h6cea7c0a_7baa7b4a,
        64'h7aea6a0e_69ae694e,
        64'h64ee740e_70ae4501,
        64'he00d3f2c_0c130000,
        64'h8c1745ab_8b930000,
        64'h9b974f2b_0b130000,
        64'h9b170381_0a93020a,
        64'h5a130017_849be03e,
        64'h020d1a13_001d179b,
        64'h03acdcbb_4cc1000c,
        64'h956302cc_dcbb0400,
        64'h0c9300e7_f6638436,
        64'h8d3289ae_892a0400,
        64'h0793e56e_f162f55e,
        64'hf95afd56_e1d2eda6,
        64'hf586e96a_e5cee9ca,
        64'hf1a202c7_073b8cba,
        64'hed667151_4e80406f,
        64'h610554a5_05130000,
        64'h951764a2_690285a6,
        64'h864a60e2_64425020,
        64'h40ef5425_05130000,
        64'h951785a2_c8015120,
        64'h40ef8932_54c50513,
        64'h00009517_05851459,
        64'h0087f463_00e45433,
        64'h942a47a5_00d41433,
        64'h440503b6_869b02f5,
        64'h053347a9_c10d4401,
        64'h8d7dfff7_c79300e7,
        64'h97b357fd_b7f559e5,
        64'h05130000_951785aa,
        64'hfb079de3_27855620,
        64'h406f6105_5b450513,
        64'h00009517_85aa6902,
        64'h64a260e2_6442e495,
        64'he04ae822_ec060007,
        64'hc483e426_97c21101,
        64'h61080813_0000a817,
        64'h93811782_cd8500e5,
        64'h55b303c6_871b02f8,
        64'h86bb4819_58d94781,
        64'h862eb78d_5d450513,
        64'h00009517_85aa5ba0,
        64'h406f6105_60450513,
        64'h00009517_690264a2,
        64'h85ca8626_60e26442,
        64'h5d4040ef_61450513,
        64'h00009517_85a2c801,
        64'h5e4040ef_84b261e5,
        64'h05130000_9517f861,
        64'h02f45433_bfc102e4,
        64'h5433a039_943e0014,
        64'h44130324_341302e4,
        64'h743302f4_57b30640,
        64'h07130287_74630630,
        64'h0713c705_02f47733,
        64'h47a90287_e6634729,
        64'h3e800793_c02102f5,
        64'h55b302f5_7433bf7d,
        64'h24078793_4685b7d9,
        64'ha0078793_468164a0,
        64'h406f6105_67450513,
        64'h00009517_85aa6902,
        64'h64a260e2_64420209,
        64'h1663e426_e822ec06,
        64'h00074903_e04a9736,
        64'h11017027_07130000,
        64'ha7173e80_07934689,
        64'h0ca7f763_3e700793,
        64'h04a76763_23f78713,
        64'h000f47b7_04a76963,
        64'h862e9ff7_87133b9a,
        64'hd7b78082_612d4501,
        64'h60ee6ae0_40ef6ce5,
        64'h05130000_9517002c,
        64'hfebff0ef_ed864505,
        64'h0c800613_002c7115,
        64'hf73ff06f_4581862e,
        64'h86b28082_614569a2,
        64'h694264e2_854a7402,
        64'h70a227c0_60ef6e65,
        64'h85930000_95970089,
        64'h0533ffd4_841b00f4,
        64'h4463ffe4_879b9c29,
        64'h6c4040ef_954a7166,
        64'h06130000_961786ce,
        64'h40a485bb_00955d63,
        64'h00098f63_842a6e20,
        64'h40ef854a_85a672e6,
        64'h06130000_9617c167,
        64'h07130000_97177366,
        64'h86930000_9697c509,
        64'hfd868693_0000a697,
        64'h893289ae_84b6f022,
        64'hf406e44e_e84aec26,
        64'h7179bfdd_760040ef,
        64'h8562b7e9_090576a0,
        64'h40ef8566_00fbe763,
        64'h0ff7f793_fe05879b,
        64'h0007c583_012a07b3,
        64'hb7810485_240578a0,
        64'h40ef2c25_05130000,
        64'ha51700f4_5b630009,
        64'h079bff04_79137a20,
        64'h40ef855a_ff2dcce3,
        64'h2d857ae0_40ef8556,
        64'ha02900f9_79134d81,
        64'hfffd4913_028d1d63,
        64'h7c4040ef_7bc50513,
        64'h00009517_0104c583,
        64'hdbe5b7c5_7d8040ef,
        64'h8562a031_7e0040ef,
        64'h85567e60_40ef31e5,
        64'h05130000_a517ffb9,
        64'h12e30905_7f8040ef,
        64'h856602fb_e2630ff7,
        64'hf793fe05_879b0007,
        64'hc5830124_87b34dc1,
        64'h49010170_40ef855a,
        64'he7a9c429_00f47793,
        64'h80826165_6da26d42,
        64'h6ce27c02_7ba27b42,
        64'h7ae26a06_69a66946,
        64'h64e67406_70a60334,
        64'h4163fff5_8d1b82ec,
        64'h8c930000_ac9783ec,
        64'h0c130000_ac170600,
        64'h0b93832b_0b130000,
        64'hab1754aa_8a930000,
        64'haa974401_ff050493,
        64'h89ae8a2a_e46ee8ca,
        64'hf486e86a_ec66f062,
        64'hf45ef85a_fc56e0d2,
        64'he4ceeca6_f0a27159,
        64'hb7cd0970_40efa007,
        64'hab230000_b79785e5,
        64'h05130000_a5178082,
        64'h61516412_60b28522,
        64'h0b5040ef_84450513,
        64'h0000a517_81c58593,
        64'h0000a597_860ac10d,
        64'h842adedf_f0ef8522,
        64'h0d5040ef_83c50513,
        64'h0000a517_83c58593,
        64'h0000a597_842a0005,
        64'h46030015_46830025,
        64'h47030035_47830045,
        64'h48030055_4883e222,
        64'he606716d_80827f01,
        64'h01137c81_39837d01,
        64'h39037d81_34837e01,
        64'h34034501_7e813083,
        64'h61658e9f_f0ef86c6,
        64'h85a61808_56326882,
        64'hfd4ff0ef_03e10513,
        64'h863e86c2_85a267c2,
        64'h6822fa4f_f0efd64e,
        64'h05210513_85a2864a,
        64'h86ba943e_7fc40413,
        64'h6762747d_97ba8107,
        64'h87931018_67857bc0,
        64'h60efd602_e83eec3a,
        64'he4428936_89b2e046,
        64'h05a10513_84aa7159,
        64'h7d313423_7d213823,
        64'h7c913c23_7e813023,
        64'h7e113423_81010113,
        64'h19d0406f_8ec50513,
        64'h0000a517_85aa8082,
        64'h61257aa2_7a4279e2,
        64'h690664a6_64464501,
        64'h60e6911a_6305985f,
        64'hf0ef85ce_86a61008,
        64'h465286ff_f0ef4601,
        64'h56fd02e1_051385a2,
        64'h83bff0ef_04400613,
        64'h04300693_04210513,
        64'h85a2943e_1451978a,
        64'h020a8793_12f11c23,
        64'h35378793_679912f1,
        64'h1b232637_879377e1,
        64'h05f060ef_04f10623,
        64'h06610513_46414799,
        64'h85ce04f1_15231010,
        64'h07930270_60efca3e,
        64'h04a10513_45810f00,
        64'h06130fc0_079308d0,
        64'h60ef0001_07a31541,
        64'h022314f1_01a31451,
        64'h05134605_85ca57fd,
        64'h0a7060ef_13f10513,
        64'h461195be_ff040593,
        64'h978a020a_879312f1,
        64'h0f234791_12f10ea3,
        64'h03700793_0cb060ef,
        64'h014107a3_1a684605,
        64'h85ca993e_978a020a,
        64'h879312f1_1d231350,
        64'h0793c83e_4a05fef4,
        64'h0913439c_b1c78793,
        64'h0000b797_0a9060ef,
        64'h852655fd_461994be,
        64'hff840493_978a020a,
        64'h8793747d_2c1040ef,
        64'hca026a85_9fc50513,
        64'h0000a517_911a89aa,
        64'hf456f852_fc4ee0ca,
        64'he4a6e8a2_ec86711d,
        64'h737db3c1_2e9040ef,
        64'h9e850513_0000a517,
        64'hbf459e25_05130000,
        64'ha51795be_978ad004,
        64'h05933507_87936785,
        64'h30d040ef_9dc50513,
        64'h0000a517_319040ef,
        64'h9d850513_0000a517,
        64'h00fa2023_4785e007,
        64'h93e3000a_2783b531,
        64'h335040ef_9e450513,
        64'h0000a517_bd293430,
        64'h40ef9e25_05130000,
        64'ha51795be_978af004,
        64'h05933504_879335b0,
        64'h40ef9ea5_05130000,
        64'ha51795be_e0040593,
        64'h978a3504_87933730,
        64'h40efd4f7_1e230000,
        64'hb7170121_5783d6f7,
        64'h13230000_b7179fe5,
        64'h05130000_a51755c2,
        64'h01015783_399040ef,
        64'h9f050513_0000a517,
        64'h01014583_01114603,
        64'h01214683_01314703,
        64'h3b5040ef_9ec50513,
        64'h0000a517_01814583,
        64'h01914603_01a14683,
        64'h01b14703_3d1040ef,
        64'h00b14703_dcf71323,
        64'h0000b717_9ec50513,
        64'h0000a517_00814583,
        64'h35215783_dcf71e23,
        64'h0000b717_00914603,
        64'h00a14683_35015783,
        64'h405040ef_9ec50513,
        64'h0000a517_35014583,
        64'h35114603_35214683,
        64'h35314703_273060ef,
        64'h01490593_4611953e,
        64'hcb840513_978a3504,
        64'h87936485_28b060ef,
        64'h0e880109_05934611,
        64'h445040ef_a1c50513,
        64'h0000a517_00fa2023,
        64'h47851007_9d63000a,
        64'h2783b311_d00d0023,
        64'h2b7060ef_9d228562,
        64'h866ab759_cc048513,
        64'hbb29cef4_2023401c,
        64'h00f40023_ce344783,
        64'h00f400a3_ce244783,
        64'h00f40123_ce144783,
        64'h00f401a3_ce044783,
        64'h2ef060ef_4611953e,
        64'hce048513_978a3507,
        64'h87936785_bfdd855a,
        64'h4611bbb1_30b060ef,
        64'h85564611_b39df00d,
        64'h00233190_60ef9d22,
        64'h953e866a_f0048513,
        64'h978a3507_87936785,
        64'ha00d953e_978a3507,
        64'h87936785_4611cd04,
        64'h85138082_3b010113,
        64'h35013d03_35813c83,
        64'h36013c03_36813b83,
        64'h37013b03_37813a83,
        64'h38013a03_38813983,
        64'h39013903_39813483,
        64'h3a013403_3a813083,
        64'h911a6305_cebff0ef,
        64'h0e8885de_86ca5672,
        64'hbd5ff0ef_35e10513,
        64'h85a24601_56fdba1f,
        64'hf0ef3721_051385a2,
        64'h04400613_04300693,
        64'h943ecec4_0413978a,
        64'h350a8793_46f11423,
        64'h35378793_679946f1,
        64'h13232637_879377e1,
        64'h3c7060ef_36f10e23,
        64'h39610513_85de4799,
        64'h464136f1_1d231010,
        64'h079338f0_60efde3e,
        64'h37a10513_45810f00,
        64'h06131020_07933f50,
        64'h60ef4731_0d230001,
        64'h03a346f1_0ca347b1,
        64'h051385a6_460557fd,
        64'h40f060ef_47410a23,
        64'h47510513_461195be,
        64'hcf440593_978a350a,
        64'h879346f1_09a30360,
        64'h07934310_60ef4741,
        64'h072346f1_05134611,
        64'h4a1195be_cf040593,
        64'h978a350a_879346f1,
        64'h06a30320_07934550,
        64'h60efc0d2_46c10513,
        64'h85a64605_94becb74,
        64'h0493c2a6_978a350a,
        64'h879346f1_15231350,
        64'h079300f1_03a3478d,
        64'h42d060ef_854a55fd,
        64'h4619993e_cf840913,
        64'h978a350a_87936430,
        64'h40efde02_54e25a52,
        64'hc0850513_0000a517,
        64'h4a7060ef_953e4611,
        64'h01490593_ce840513,
        64'h978a350a_87934bd0,
        64'h60ef013c_a023953e,
        64'h46110109_0593ce44,
        64'h05134985_978a350a,
        64'h87936a85_16079263,
        64'h000ca783_3ae79063,
        64'h470936e7_84634719,
        64'h24e78163_0007859b,
        64'h747d4715_00614783,
        64'hf8e79ce3_0ff00713,
        64'h24e78563_03800713,
        64'haad94605_cb648513,
        64'hfae798e3_03500713,
        64'h22e78063_03300713,
        64'h00f76e63_22e78363,
        64'h03600713_b759e00d,
        64'h00235390_60ef9d22,
        64'h953e866a_e0048513,
        64'h978a3507_87936785,
        64'hfee794e3_473d22e7,
        64'h85634731_b77d70b0,
        64'h40efe225_05130000,
        64'ha51785b6_22e78963,
        64'hcc848513_470d2ae7,
        64'h89634705_02f76263,
        64'h24e78163_471904f7,
        64'h6b6326e7_8d630007,
        64'h869b01a9_89bb0589,
        64'h02a00713_29890f07,
        64'hc7830015_cd030139,
        64'h07b395ca_0f098593,
        64'h9c3a9b3a_49818a36,
        64'h8cb28bae_d0048c13,
        64'hcb848b13_970a3507,
        64'h87139aba_cd848a93,
        64'h970a3507_871374fd,
        64'h678526f7_11634789,
        64'h00054703_a0017930,
        64'h40efd325_05130000,
        64'ha51785aa_00e7ea63,
        64'h892a5800_073797aa,
        64'hd0040023_f0040023,
        64'he0040023_ca040b23,
        64'hce042023_d00007b7,
        64'h943e747d_978a911a,
        64'h35078793_35a13823,
        64'h35913c23_37813023,
        64'h37713423_37613823,
        64'h37513c23_39413023,
        64'h39313423_38913c23,
        64'h3a113423_39213823,
        64'h3a813023_6785737d,
        64'hc5010113_fadff06f,
        64'h614564e2_00e4859b,
        64'h70a27402_852200f4,
        64'h162347a1_673060ef,
        64'h85b64619_852266a2,
        64'h67f060ef_e436f406,
        64'h46190519_84b2842a,
        64'hec26f022_71798082,
        64'h01416402_60a28522,
        64'hfa5ff0ef_e4064501,
        64'h85aa8622_0005841b,
        64'he0221141_bff105a1,
        64'h25050116_b02396ba,
        64'h010686bb_0035169b,
        64'h0005b883_808280c7,
        64'h3823973e_678500f5,
        64'h47636805_450102d7,
        64'hc7bb2785_0077e793,
        64'hfff6079b_8007bc23,
        64'h97ba46a1_67856398,
        64'h13878793_0000b797,
        64'h80826145_740270a2,
        64'h00f41523_fff7c793,
        64'h9fb94107_d71b9fb9,
        64'h93411742_4107579b,
        64'hfed79ce3_9f31ffe7,
        64'hd6030789_470187a2,
        64'h01440693_733060ef,
        64'h01040513_002c4611,
        64'h73f060ef_00c40513,
        64'h00041523_006c4611,
        64'h00f404a3_47c57550,
        64'h60efec3e_00840513,
        64'h00041323_082c4621,
        64'h47c17690_60ef0044,
        64'h05130161_05934609,
        64'h777060ef_00f11b23,
        64'hc4360509_084c57fd,
        64'h460900f1_1a238fd9,
        64'h0087979b_0ff77713,
        64'h0087d713_c632842a,
        64'h419c00f5_10230457,
        64'h879b6785_c19c27d1,
        64'hf022f406_7179419c,
        64'h80820005_132300f5,
        64'h122300d5_112300c5,
        64'h10238fd9_0087979b,
        64'h0ff77713_c19c0087,
        64'hd7138ed9_06a20086,
        64'hd71b8e59_27a10622,
        64'h0086571b_419cc19c,
        64'h2785c319_0017f713,
        64'h419cbfcd_fda00513,
        64'h80826121_74a27442,
        64'h70e29782_85a66562,
        64'h701ce509_c39ff0ef,
        64'h842a0830_65a2c105,
        64'hc7dff0ef_84b2e42e,
        64'hf822fc06_f4267139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2655c,
        64'h862686ca_6562e519,
        64'hc75ff0ef_083065a2,
        64'hc115cb7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2615c,
        64'h862686ca_6562e519,
        64'hcb5ff0ef_083065a2,
        64'hc115cf7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hb7e16522_f569cdbf,
        64'hf0ef8526_85ce0030,
        64'hbfc90284_8493c501,
        64'h689060ef_854a608c,
        64'h27c050ef_855285ca,
        64'h60908082_61216a42,
        64'h69e27902_74a27442,
        64'h70e24501_00849b63,
        64'h942602f4_043302ea,
        64'h0a130000_aa1789ae,
        64'h892afc06_e852ec4e,
        64'hf04a0280_079302f4,
        64'h043b840d_8c053a24,
        64'h84930000_b4973aa4,
        64'h04130000_b417f426,
        64'hf822639c_26478793,
        64'h0000b797_7139bfdd,
        64'h45018082_61056442,
        64'h60e2fda0_05138302,
        64'h610560e2_65a26442,
        64'h85220003_0e630205,
        64'h3303c919_db9ff0ef,
        64'he42eec06_4108842a,
        64'he8221101_bfc56562,
        64'hf96dd97f_f0ef0830,
        64'h80826145_70a24501,
        64'he50965a2_de1ff0ef,
        64'hf406e42e_7179bfc1,
        64'h5479fcf7_1be30ff0,
        64'h079300c7_c70367a2,
        64'h034080ef_6522f565,
        64'h842adcff_f0ef85a6,
        64'h00308522_80826145,
        64'h64e27402_70a28522,
        64'h54350600_80ef0ee5,
        64'h05130000_a51700f4,
        64'hcf63445c_380050ef,
        64'h0f050513_0000a517,
        64'h85a6842a_c11dfda0,
        64'h0413e47f_f0ef84ae,
        64'hf406ec26_f0227179,
        64'h80826145_694264e2,
        64'h740270a2_852209a0,
        64'h80ef6522_3b8050ef,
        64'h11850513_0000a517,
        64'h864a608c_ed01842a,
        64'he45ff0ef_84aa85ca,
        64'h0030c11d_fda00413,
        64'he8dff0ef_892eec26,
        64'hf406e84a_f0227179,
        64'hb7d92405_0d8080ef,
        64'h65223f60_50ef854e,
        64'h85a20127_896300c7,
        64'hc78367a2_ed09e83f,
        64'hf0ef8526_85a20030,
        64'h80826121_69e27902,
        64'h74a27442_70e200f4,
        64'h496344dc_17498993,
        64'h0000a997_0ff00913,
        64'h440184aa_cd01eebf,
        64'hf0efec4e_f04af426,
        64'hf822fc06_7139bfd5,
        64'h54798082_61457402,
        64'h70a28522_13e080ef,
        64'h00f70963_00c54703,
        64'h0ff00793_6562e911,
        64'h842aee7f_f0ef0830,
        64'h65a2c105_fda00413,
        64'hf2dff0ef_e42ef406,
        64'hf0227179_b7c1fda0,
        64'h0513bf65_24051780,
        64'h80ef4981_652249a0,
        64'h50ef8552_00099563,
        64'h2485cb99_0087c783,
        64'h67a2ed19_f29ff0ef,
        64'h854a85a2_00308082,
        64'h61216a42_69e27902,
        64'h74a27442_70e24501,
        64'hc0915535_00f44d63,
        64'h00c92783_00ca0a13,
        64'h0000ba17_44014481,
        64'h4985892a_cd31f9bf,
        64'hf0efe852_ec4ef04a,
        64'hf426f822_fc067139,
        64'hbfe54501_80820141,
        64'h60a26108_c509fbbf,
        64'hf0efe406_1141b7f5,
        64'h02870713_fea68de3,
        64'h47148082_853a4701,
        64'h00e79563_97ba02d7,
        64'h87b30280_069302d7,
        64'h87bb878d_8f9961a7,
        64'h87930000_b7976294,
        64'h62470713_0000b717,
        64'h4d868693_0000b697,
        64'hb7edfda0_07138302,
        64'h853e85b2_00030563,
        64'h01853303_8082853a,
        64'he21c97b6_470102a7,
        64'h87b30a00_051300b7,
        64'hd963454c_0005cc63,
        64'h5735c285_87ae6914,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h000a2e2e_2e746e65,
        64'h6d6f6d20_61207469,
        64'h61772065_7361656c,
        64'h50202165_6e616972,
        64'h41206d6f_7266206f,
        64'h6c6c6548_ffdff06f,
        64'h10500073_34102373,
        64'h342022f3_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_45e090ef,
        64'hfec5c6e3_02058593,
        64'h0005bc23_0005b823,
        64'h0005b423_0005b023,
        64'hd9060613_0000c617,
        64'h83058593_0000c597,
        64'h30579073_09078793,
        64'h00000797_00078067,
        64'h40b787b3_00d787b3,
        64'h01478793_00000797,
        64'hfcc5cce3_02068693,
        64'h02058593_00e6bc23,
        64'h0185b703_00e6b823,
        64'h0105b703_00e6b423,
        64'h0085b703_00e6b023,
        64'h0005b703_0006b703,
        64'hff810113_01b11113,
        64'h0110011b_fe0e9ae3,
        64'h0085b703_fffe8e93,
        64'h0005b703_240e8e9b,
        64'h000f4eb7_01169693,
        64'h3ff6869b_000046b7,
        64'h81c60613_0000c617,
        64'hfc058593_00000597,
        64'h000280e7_13050513,
        64'h00000517_07a28293,
        64'h00008297_000280e7,
        64'h05428293_00008297,
        64'h01111113_3ff1011b,
        64'h00004137_11249463,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
