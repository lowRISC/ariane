/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'h01111113fff1011b0000613711249463, /*    1 */
128'h00008297000280e708c2829300008297, /*    2 */
128'h000280e713050513000005170b228293, /*    3 */
128'h9c5606130000c617fc05859300000597, /*    4 */
128'h000f4eb701169693fff6869b000066b7, /*    5 */
128'h0085b703fffe8e930005b703240e8e9b, /*    6 */
128'hff81011301b111130110011bfe0e9ae3, /*    7 */
128'h0085b70300e6b0230005b7030006b703, /*    8 */
128'h0185b70300e6b8230105b70300e6b423, /*    9 */
128'hfcc5cce3020686930205859300e6bc23, /*   10 */
128'h40b787b300d787b30147879300000797, /*   11 */
128'h30579073090787930000079700078067, /*   12 */
128'h1c8606130000c617a30585930000c597, /*   13 */
128'h0005bc230005b8230005b4230005b023, /*   14 */
128'h020004b767a090effec5c6e302058593, /*   15 */
128'h02000937004484930124a02300100913, /*   16 */
128'h3440297310500073ff24c6e34009091b, /*   17 */
128'hf1402973020004b7fe090ae300897913, /*   18 */
128'h0004a903000920230099093300291913, /*   19 */
128'h4009091b0200093700448493fe091ee3, /*   20 */
128'h1050007334102373342022f3ff24c6e3, /*   21 */
128'h41206d6f7266206f6c6c6548ffdff06f, /*   22 */
128'h617720657361656c502021656e616972, /*   23 */
128'h000a2e2e2e746e656d6f6d2061207469, /*   24 */
128'h00000000000000000000000000000000, /*   25 */
128'h00000000000000000000000000000000, /*   26 */
128'h00000000000000000000000000000000, /*   27 */
128'h00000000000000000000000000000000, /*   28 */
128'h00000000000000000000000000000000, /*   29 */
128'h00000000000000000000000000000000, /*   30 */
128'h00000000000000000000000000000000, /*   31 */
128'hd963454c0005cc635735c28587ae6914, /*   32 */
128'he21c97b6470102a787b30a00051300b7, /*   33 */
128'h853e85b200030563018533038082853a, /*   34 */
128'h708686930000b697b7edfda007138302, /*   35 */
128'h87930000b79762947d0707130000b717, /*   36 */
128'h87b30280069302d787bb878d8f997c67, /*   37 */
128'h47148082853a470100e7956397ba02d7, /*   38 */
128'hf0efe4061141b7f502870713fea68de3, /*   39 */
128'hbfe545018082014160a26108c509fbbf, /*   40 */
128'hf0efe852ec4ef04af426f822fc067139, /*   41 */
128'h0000ba17440144814985892acd31f9bf, /*   42 */
128'he091450100f44d6300c9278328ca0a13, /*   43 */
128'h61216a4269e2790274a2744270e25535, /*   44 */
128'h67a2ed19f29ff0ef854a85a200308082, /*   45 */
128'h50ef8552000995632485cb990087c783, /*   46 */
128'h0513bf652405222080ef498165224720, /*   47 */
128'hf2dff0efe42ef406f0227179b7c1fda0, /*   48 */
128'h842aee7ff0ef083065a2c105fda00413, /*   49 */
128'h00f7096300c547030ff007936562e911, /*   50 */
128'h547980826145740270a285221e8080ef, /*   51 */
128'hf0efec4ef04af426f822fc067139bfd5, /*   52 */
128'h0000a9970ff00913440184aacd01eebf, /*   53 */
128'h74a2744270e200f4496344dc3a498993, /*   54 */
128'hf0ef852685a200308082612169e27902, /*   55 */
128'h85a20127896300c7c78367a2ed09e83f, /*   56 */
128'hb7d92405182080ef65223ce050ef854e, /*   57 */
128'he8dff0ef892eec26f406e84af0227179, /*   58 */
128'he45ff0ef84aa85ca0030c11dfda00413, /*   59 */
128'h348505130000a517864a608ced01842a, /*   60 */
128'h740270a28522144080ef6522390050ef, /*   61 */
128'hf406ec26f022717980826145694264e2, /*   62 */
128'h85a6842ac11dfda00413e47ff0ef84ae, /*   63 */
128'hcf63445c358050ef320505130000a517, /*   64 */
128'h543510a080ef31e505130000a51700f4, /*   65 */
128'h003085228082614564e2740270a28522, /*   66 */
128'h0de080ef6522f565842adcfff0ef85a6, /*   67 */
128'h5479fcf71be30ff0079300c7c70367a2, /*   68 */
128'he50965a2de1ff0eff406e42e7179bfc1, /*   69 */
128'hf96dd97ff0ef08308082614570a24501, /*   70 */
128'he42eec064108842ae8221101bfc56562, /*   71 */
128'h852200030e6302053303c919db9ff0ef, /*   72 */
128'h60e2fda005138302610560e265a26442, /*   73 */
128'h0000b7977139bfdd4501808261056442, /*   74 */
128'h04130000b417f426f822639c49478793, /*   75 */
128'h043b840d8c0554e484930000b4975564, /*   76 */
128'h892afc06e852ec4ef04a0280079302f4, /*   77 */
128'h942602f4043325ea0a130000aa1789ae, /*   78 */
128'h69e2790274a2744270e2450100849b63, /*   79 */
128'h254050ef855285ca6090808261216a42, /*   80 */
128'hbfc902848493c501681060ef854a608c, /*   81 */
128'hb7e16522f569cdbff0ef852685ce0030, /*   82 */
128'h84b68432e42efc06f04af426f8227139, /*   83 */
128'hcb5ff0ef083065a2c115cf7ff0ef893a, /*   84 */
128'h70e2978285a2615c862686ca6562e519, /*   85 */
128'hbfc5fda0051380826121790274a27442, /*   86 */
128'h84b68432e42efc06f04af426f8227139, /*   87 */
128'hc75ff0ef083065a2c115cb7ff0ef893a, /*   88 */
128'h70e2978285a2655c862686ca6562e519, /*   89 */
128'hbfc5fda0051380826121790274a27442, /*   90 */
128'hc7dff0ef84b2e42ef822fc06f4267139, /*   91 */
128'h701ce509c39ff0ef842a083065a2c105, /*   92 */
128'h8082612174a2744270e2978285a66562, /*   93 */
128'h2785c3190017f713419cbfcdfda00513, /*   94 */
128'hd71b8e5927a106220086571b419cc19c, /*   95 */
128'h0ff77713c19c0087d7138ed906a20086, /*   96 */
128'h122300d5112300c510238fd90087979b, /*   97 */
128'hf022f4067179419c80820005132300f5, /*   98 */
128'h419c00f510230457879b6785c19c27d1, /*   99 */
128'h0087979b0ff777130087d713c632842a, /*  100 */
128'hc4360509084c57fd460900f11a238fd9, /*  101 */
128'h051301610593460976b060ef00f11b23, /*  102 */
128'h00041323082c462147c175d060ef0044, /*  103 */
128'h00f404a347c5749060efec3e00840513, /*  104 */
128'h733060ef00c4051300041523006c4611, /*  105 */
128'h01440693727060ef01040513002c4611, /*  106 */
128'hfed79ce39f31ffe7d6030789470187a2, /*  107 */
128'h9fb94107d71b9fb9934117424107579b, /*  108 */
128'h80826145740270a200f41523fff7c793, /*  109 */
128'h97b64721678563942b8787930000b797, /*  110 */
128'hc7bb27850077e793fff6079b8007bc23, /*  111 */
128'h678500f747630005071b6805450102e7, /*  112 */
128'h00e588b300351713808280c6b82396be, /*  113 */
128'hbfe1050501173023973697420008b883, /*  114 */
128'he406450185aa86220005841be0221141, /*  115 */
128'h717980820141640260a28522fa1ff0ef, /*  116 */
128'he436f4064619051984b2842aec26f022, /*  117 */
128'h663060ef85b64619852266a266f060ef, /*  118 */
128'h00e4859b70a27402852200f4162347a1, /*  119 */
128'h6785737dc5010113fadff06f614564e2, /*  120 */
128'h38913c233a113423392138233a813023, /*  121 */
128'h3761382337513c233941302339313423, /*  122 */
128'h35a1382335913c233781302337713423, /*  123 */
128'hd00007b7943e747d978a911a35078793, /*  124 */
128'hf0040023e0040023ca040b23ce042023, /*  125 */
128'h00e7ea63892a5800073797aad0040023, /*  126 */
128'ha001767040eff5e505130000a51785aa, /*  127 */
128'h871374fd678524f71d63478900054703, /*  128 */
128'h970a350787139abacd848a93970a3507, /*  129 */
128'h49818a368cb28baed0048c13cb848b13, /*  130 */
128'hcd03013907b395ca0f0985939c3a9b3a, /*  131 */
128'h89bb058902a0071329890f07c7830015, /*  132 */
128'h22e78f63471904f76b6326e78b6301a9, /*  133 */
128'hcc848513470d2ae78963470502f76263, /*  134 */
128'h40ef062505130000a51785be22e78763, /*  135 */
128'hfee794e3473d22e783634731bf4d6e30, /*  136 */
128'h953e866ae0048513978a350787936785, /*  137 */
128'h03600713b769e00d002352d060ef9d22, /*  138 */
128'h20e78e630330071300f76e6322e78163, /*  139 */
128'haac94605cb648513fae798e303500713, /*  140 */
128'hf8e79ce30ff0071324e7856303800713, /*  141 */
128'h8363479924f58363747d479500614583, /*  142 */
128'h16079263000ca7833af59f63478938f5, /*  143 */
128'h0593ce4405134985978a350a87936a85, /*  144 */
128'h87934b5060ef013ca023953e46110109, /*  145 */
128'h953e461101490593ce840513978a350a, /*  146 */
128'h54e25a52e3c505130000a51749f060ef, /*  147 */
128'hcf840913978a350a879361f040efde02, /*  148 */
128'h03a3478d429060ef854a55fd4619993e, /*  149 */
128'h978a350a879346f115231350079300f1, /*  150 */
128'h46c1051385a6460594becb740493c2a6, /*  151 */
128'h879346f106a30320079344d060efc0d2, /*  152 */
128'h051346114a1195becf040593978a350a, /*  153 */
128'h09a303600793429060ef4741072346f1, /*  154 */
128'h461195becf440593978a350a879346f1, /*  155 */
128'h460557fd407060ef47410a2347510513, /*  156 */
128'h0d23000103a346f10ca347b1051385a6, /*  157 */
128'h45810f000613102007933ed060ef4731, /*  158 */
128'h1d231010079338b060efde3e37a10513, /*  159 */
128'h36f10e233961051385de4799464136f1, /*  160 */
128'h679946f113232637879377e13bf060ef, /*  161 */
128'h0413978a350a879346f1142335378793, /*  162 */
128'h051385a20440061304300693943ecec4, /*  163 */
128'h35e1051385a2460156fdba5ff0ef3721, /*  164 */
128'hcf3ff0ef0e8885de86ca5672bd9ff0ef, /*  165 */
128'h398134833a0134033a813083911a6305, /*  166 */
128'h37813a8338013a033881398339013903, /*  167 */
128'h35813c8336013c0336813b8337013b03, /*  168 */
128'h4611cd04851380823b01011335013d03, /*  169 */
128'h87936785a00d953e978a350787936785, /*  170 */
128'h60ef9d22953e866af0048513978a3507, /*  171 */
128'h303060ef85564611b3bdf00d00233110, /*  172 */
128'h978a350787936785bfdd855a4611b395, /*  173 */
128'hce0457832e7060ef4611953ece048513, /*  174 */
128'h578300f411238fd90087979b0087d71b, /*  175 */
128'h00f410238fd90087979b0087d71bce24, /*  176 */
128'h866ab749cc048513bb39cef42023401c, /*  177 */
128'h2783b321d00d00232ab060ef9d228562, /*  178 */
128'h0000a51700fa2023478512079a63000a, /*  179 */
128'h0e8801090593461141d040efc4c50513, /*  180 */
128'hcb840513978a35048793648527f060ef, /*  181 */
128'h35314703267060ef014905934611953e, /*  182 */
128'h0000a517350145833511460335214683, /*  183 */
128'h00a14683350157833dd040efc1c50513, /*  184 */
128'h35215783fcf71e230000b71700914603, /*  185 */
128'h0000b717c1c505130000a51700814583, /*  186 */
128'h01b147033a9040ef00b14703fcf71323, /*  187 */
128'h0000a517018145830191460301a14683, /*  188 */
128'h012146830131470338d040efc1c50513, /*  189 */
128'hc20505130000a5170101458301114603, /*  190 */
128'h05130000a51755c201015783371040ef, /*  191 */
128'hb71701215783f6f713230000b717c2e5, /*  192 */
128'hf6bb02f5d63b03c00793f4f71e230000, /*  193 */
128'h02f5d5bbe107879b678502f6763b02f5, /*  194 */
128'h95bee0040593978a35048793331040ef, /*  195 */
128'h35048793319040efc08505130000a517, /*  196 */
128'hc00505130000a51795be978af0040593, /*  197 */
128'h40efc0a505130000a517bbf5301040ef, /*  198 */
128'h20234785de0794e3000a2783b3fd2f30, /*  199 */
128'ha5172d7040efbfe505130000a51700fa, /*  200 */
128'h3507879367852cb040efc02505130000, /*  201 */
128'hc08505130000a51795be978ad0040593, /*  202 */
128'hb34d2a7040efc0e505130000a517bf45, /*  203 */
128'hf852fc4ee0cae4a6e8a2ec86711d737d, /*  204 */
128'h6a85c22505130000a517911a89aaf456, /*  205 */
128'h0493978a020a8793747d27f040efca02, /*  206 */
128'hb797087060ef852655fd461994beff84, /*  207 */
128'hc83e4a05fef40913439cc82787930000, /*  208 */
128'h993e978a020a879312f11d2313500793, /*  209 */
128'h07930a5060ef014107a31a68460585ca, /*  210 */
128'h020a879312f10f23479112f10ea30370, /*  211 */
128'h60ef13f10513461195beff040593978a, /*  212 */
128'h14f101a314510513460585ca57fd0810, /*  213 */
128'h0fc00793067060ef000107a315410223, /*  214 */
128'h005060efca3e04a1051345810f000613, /*  215 */
128'h05134641479985ce04f1152310100793, /*  216 */
128'h2637879377e1039060ef04f106230661, /*  217 */
128'h879312f11c2335378793679912f11b23, /*  218 */
128'h06930421051385a2943e1451978a020a, /*  219 */
128'h02e1051385a2821ff0ef044006130430, /*  220 */
128'h85ce86a610084652855ff0ef460156fd, /*  221 */
128'h64a66446450160e6911a630596fff0ef, /*  222 */
128'ha51785aa808261257aa27a4279e26906, /*  223 */
128'hf0a2f486715915b0406fb12505130000, /*  224 */
128'h05a1051384aa81010113e4cee8caeca6, /*  225 */
128'h60efd602e83eec3ae442893689b2e046, /*  226 */
128'h6762747d97ba81078793101867857a00, /*  227 */
128'h0521051385a2864a86ba943e7fc40413, /*  228 */
128'h863e86c285a267c26822f94ff0efd64e, /*  229 */
128'h85a6180856326882fc4ff0ef03e10513, /*  230 */
128'h7406450170a67f0101138ddff0ef86c6, /*  231 */
128'he222e606716d8082616569a6694664e6, /*  232 */
128'h00254703003547830045480300554883, /*  233 */
128'h85930000a597842a0005460300154683, /*  234 */
128'h85220a7040efa76505130000a517a765, /*  235 */
128'h85930000a597860ac10d842ae01ff0ef, /*  236 */
128'h8522087040efa7e505130000a517a565, /*  237 */
128'ha98505130000a51780826151641260b2, /*  238 */
128'h7159b7cd069040efc007a8230000b797, /*  239 */
128'hec66f062f45ef85afc56e0d2e4ceeca6, /*  240 */
128'h44818aae89aae46ee8caf0a2f486e86a, /*  241 */
128'ha70b0b130000ab17740a0a130000aa17, /*  242 */
128'h0000ac97a7cc0c130000ac1706000b93, /*  243 */
128'h035441630004841bfff58d1ba6cc8c93, /*  244 */
128'h7b427ae26a0669a6694664e6740670a6, /*  245 */
128'hc01d808261656da26d426ce27c027ba2, /*  246 */
128'hff0489137e8040ef855ae39d00f47793, /*  247 */
128'h5b0505130000a51702879d630009079b, /*  248 */
128'hc583009987b37ca040ef85527d0040ef, /*  249 */
128'h12637b6040efa16505130000a5170007, /*  250 */
128'h87b3a80500f979134d81fffd4913068d, /*  251 */
128'he7630ff7f793fe05879b0007c5830129, /*  252 */
128'h40ef8562b75d090578c040ef856600fb, /*  253 */
128'hff2dcce32d8577a040ef8552bfdd7820, /*  254 */
128'h079b4124093b76a040ef00f4f913855a, /*  255 */
128'h40ef532505130000a51700f45a630009, /*  256 */
128'h879b0007c583012987b3bf1504857520, /*  257 */
128'h734040ef856600fbe7630ff7f793fe05, /*  258 */
128'hec267179bfdd72a040ef8562b7f10905, /*  259 */
128'ha697893289ae84b6f022f406e44ee84a, /*  260 */
128'h968686930000a697c5091ba686930000, /*  261 */
128'h960606130000a617e187071300009717, /*  262 */
128'h5d6300098f63842a6ac040ef854a85a6, /*  263 */
128'h948606130000a61786ce40a485bb0095, /*  264 */
128'h00f44463ffe4879b9c2968e040ef954a, /*  265 */
128'h918585930000a59700890533ffd4841b, /*  266 */
128'h69a2694264e2854a740270a226a060ef, /*  267 */
128'h7115f73ff06f4581862e86b280826145, /*  268 */
128'h002cfebff0efed8645050c800613002c, /*  269 */
128'h450160ee678040ef900505130000a517, /*  270 */
128'h6963862e9ff787133b9ad7b78082612d, /*  271 */
128'h079304a7676323f78713000f47b704a7, /*  272 */
128'h0000b7173e80079346890ca7fc633e70, /*  273 */
128'hec0600074903e04a9736110187470713, /*  274 */
128'h690264a260e2644202091663e426e822, /*  275 */
128'h6140406f61058a6505130000a51785aa, /*  276 */
128'hbf7d240787934685b7d9a00787934681, /*  277 */
128'h47293e800793c81502f555b302f57433, /*  278 */
128'h0713cf3902f4773346a547a90687e263, /*  279 */
128'h743302f457b30640071300877d630630, /*  280 */
128'h0000a517943e001444130324341302e4, /*  281 */
128'ha51785a2c8015ba040ef84b285c50513, /*  282 */
128'h862660e264425aa040ef852505130000, /*  283 */
128'h6105842505130000a517690264a285ca, /*  284 */
128'hf46302f45733bf6102e454335900406f, /*  285 */
128'h0000951785aabf554401bf51843a0086, /*  286 */
128'h86bb459958d94701862ebfa17fc50513, /*  287 */
128'h1702cf8500f557b3883e03c6879b02e8, /*  288 */
128'he426972e1101776585930000a5979301, /*  289 */
128'h60e26442e495e04ae822ec0600074483, /*  290 */
128'h61057da505130000951785aa690264a2, /*  291 */
128'h0000951785aafab71ce327055200406f, /*  292 */
128'hfff7471301071733577db7f57c450513, /*  293 */
128'h03b6869b02e505334729c10d44018d79, /*  294 */
128'h746301045433942a472500d414334405, /*  295 */
128'h770505130000951785be078514590087, /*  296 */
128'h05130000951785a2c8014ce040ef8932, /*  297 */
128'h690285a6864a60e264424be040ef7665, /*  298 */
128'h4a40406f610576e505130000951764a2, /*  299 */
128'hf54ef94ae1a202c7073b8cbafce67155, /*  300 */
128'he162e55ee95aed56f152fd26e586f8ea, /*  301 */
128'hf66384368d3289ae892a04000793f4ee, /*  302 */
128'h4cc1000c956302ccdcbb04000c9300e7, /*  303 */
128'h001a849b020d1a13001d1a9b03acdcbb, /*  304 */
128'h00009b9771cb0b1300009b17020a5a13, /*  305 */
128'h4501e00d5dcc0c1300008c17684b8b93, /*  306 */
128'h6b4a6aea7a0a79aa794a74ea640e60ae, /*  307 */
128'h85ca808261697da67d467ce66c0a6baa, /*  308 */
128'h00040d9b408040ef6d85051300009517, /*  309 */
128'h482146914781874e000c8d9b008cf463, /*  310 */
128'h9381020d979305b66b630007861b4889, /*  311 */
128'h083803bd06bb0d9de56399be034787b3, /*  312 */
128'h0b079c630006881b02e0089385ba4781, /*  313 */
128'h8c23e036694505130000951797ba1098, /*  314 */
128'h9281168241b4043b66823ae040effa07, /*  315 */
128'h02dd1963b79d557dd13d0b8070ef9936, /*  316 */
128'h1602c19095aa26010828002795934310, /*  317 */
128'h6702376040efe03ae43e855a85d69201, /*  318 */
128'h1963bf9d4691482107859752488967a2, /*  319 */
128'hbfd1e19095aa0828003795936310010d, /*  320 */
128'h164208280017959300075603011d1d63, /*  321 */
128'h082c00074603bf6d00c5902395aa9241, /*  322 */
128'he03e855eb76500c580230ff6761395be, /*  323 */
128'hbf253cfdfe97eae3278567820e4070ef, /*  324 */
128'h0005450300cc053300074603bfdd4781, /*  325 */
128'h54634186561b0186161bc51909757513, /*  326 */
128'h87aa1582b70d07052785011700230006, /*  327 */
128'h8f8d25058082e21c00b7f46345019181, /*  328 */
128'h0088458189aa04000613fd4e7115bfd5, /*  329 */
128'hed5ef15af556f952e1cae5a6e9a2ed86, /*  330 */
128'h07130000a71767869982e16ae566e962, /*  331 */
128'h440106e79d63557983e107e2631848e7, /*  332 */
128'h9b9756ab0b1300009b174a8503800a13, /*  333 */
128'h9d1708000cb780000c375a2b8b930000, /*  334 */
128'h656600f464630781578357ad0d130000, /*  335 */
128'h9dbd0028038006137786028a05bba091, /*  336 */
128'h855a85a2cfbd77c20957926347a29982, /*  337 */
128'h018487b37482040908637922240040ef, /*  338 */
128'h40ef51a505130000951785a60397e863, /*  339 */
128'h7a4a79ea690e64ae644e60ee55752220, /*  340 */
128'h8082612d6d0a6caa6c4a6bea7b0a7aaa, /*  341 */
128'h061b45c21f8040ef856a86ca85a66642, /*  342 */
128'h79020097ff6377a274c2998285260009, /*  343 */
128'h86261d6040ef855e85ca993e86268c9d, /*  344 */
128'h057e4505bfb124057ed050ef854a4581, /*  345 */
128'h580707130000a7178082400005378082, /*  346 */
128'he30895360017869300756513157d631c, /*  347 */
128'h67858082953e057e450597aa20000537, /*  348 */
128'h871308a74463862a0ce5076382078713, /*  349 */
128'h496306e60b634c650513000095178087, /*  350 */
128'hc3ad4a250513000095178006079b04c7, /*  351 */
128'hc963522505130000951787f787936785, /*  352 */
128'h000095979e3d11417c07879b77fd04c7, /*  353 */
128'h40efe4064e4505130000a51751458593, /*  354 */
128'h808201414d4505130000a51760a210e0, /*  355 */
128'h00e60a63474505130000951781078713, /*  356 */
128'hfaf612e3474505130000951781878793, /*  357 */
128'h09e34925051300009517830787138082, /*  358 */
128'h0513000095178287879300c74963fee6, /*  359 */
128'h480505130000951783878713bfe946e5, /*  360 */
128'h480505130000951784078793fce608e3, /*  361 */
128'hf022717980824365051300009517bf75, /*  362 */
128'h07bb00a5893b440184aaf406e84aec26, /*  363 */
128'h942a904114420104551302f044634099, /*  364 */
128'h1542fff54513740270a2952201045513, /*  365 */
128'h0068460985a6808261459141694264e2, /*  366 */
128'h979b0087d71b048900c157836df050ef, /*  367 */
128'hbf45943e93c117c200f117238fd90087, /*  368 */
128'h8793f44ef84afc26e486e0a26785715d, /*  369 */
128'h0e636dd7879367a13cf50463842e8067, /*  370 */
128'h082884b205e9440799638005079b0af5, /*  371 */
128'ha517461985ca0064091368d050ef4611, /*  372 */
128'h079301744583679050ef3d2505130000, /*  373 */
128'h1cf5816347b108b7e76332f5886302e0, /*  374 */
128'h478502b7e3631af58263479104b7e563, /*  375 */
128'h83633ba5051300009517478910f58463, /*  376 */
128'ha4157c7030ef556505130000951702f5, /*  377 */
128'h3c0505130000951747a118f581634799, /*  378 */
128'h2cf5816347f5a4297ad030effef591e3, /*  379 */
128'h0000951747d916f5896347c500b7ed63, /*  380 */
128'h856302100793bf6dfef580e33dc50513, /*  381 */
128'h051300009517faf596e3029007932af5, /*  382 */
128'h04b7e2632cf5816306200793b7c93f65, /*  383 */
128'h02f0079300b7ef632af5816303300793, /*  384 */
128'h3f850513000095170320079328f58663, /*  385 */
128'h079328f5836305c00793b7bdf8f58ae3, /*  386 */
128'hbf91f6f58de340e505130000951705e0, /*  387 */
128'h0670079300b7ef6328f5856308400793, /*  388 */
128'h420505130000951706c0079326f58a63, /*  389 */
128'h079326f5876308900793b73df4f58ae3, /*  390 */
128'h9517f0f59ce30880079326f588630ff0, /*  391 */
128'h0000a79701e45703b73d42a505130000, /*  392 */
128'h12f713632dc989930000a9972e47d783, /*  393 */
128'h10f71b632ce7d7830000a79702045703, /*  394 */
128'h0000a5974619519050ef852285ca4619, /*  395 */
128'h012301a45783509050ef854a29c58593, /*  396 */
128'h859b01c4578300f41f23020412230204, /*  397 */
128'h1d230009d78302f4102302240513fde4, /*  398 */
128'h579bdb3ff0ef00f41e230029d78300f4, /*  399 */
128'h862602a4122300a11e238d5d05220085, /*  400 */
128'h051300009517a06ddcdfe0ef450185a2, /*  401 */
128'h9517b56123c5051300009517bd4922e5, /*  402 */
128'h0264470302444783bdbd24a505130000, /*  403 */
128'h01c1178300f10e230254478300f10ea3, /*  404 */
128'h470300e10e2327810274470300e10ea3, /*  405 */
128'h0e230234470300e10ea301c119030224, /*  406 */
128'ha79704e79b6301c156830450071300e1, /*  407 */
128'h85930000a597461947e21ad79f230000, /*  408 */
128'h2f230000a71719e505130000a5171965, /*  409 */
128'h0000a79766a2476242b050efe43618f7, /*  410 */
128'h60ef450102a40593ff89061b17478793, /*  411 */
128'h8082616179a2794274e2640660a654e0, /*  412 */
128'h2f230000a71747e204e6946304300713, /*  413 */
128'ha797c799439c162787930000a79714f7, /*  414 */
128'h86930000a697f7e9439c152787930000, /*  415 */
128'h85930000a597142606130000a6171466, /*  416 */
128'h4d200713b765d73fe0ef02a405131465, /*  417 */
128'h535030ef164505130000951702e79863, /*  418 */
128'h1605051300009517ccaff0ef852285a6, /*  419 */
128'hbf95cb4ff0ef02a4051385ca521030ef, /*  420 */
128'h17fd67c101e45703f6e787e35fe00713, /*  421 */
128'ha5974611f4f70de302045703f6f701e3, /*  422 */
128'h9517b799357050ef0868102585930000, /*  423 */
128'h1405051300009517b33d13a505130000, /*  424 */
128'h00009517bb291565051300009517b315, /*  425 */
128'hb31917a5051300009517bb0116450513, /*  426 */
128'h051300009517b9f51805051300009517, /*  427 */
128'h9517b1e51ac5051300009517b9cd19e5, /*  428 */
128'h1e85051300009517b9f91c2505130000, /*  429 */
128'h0265d703b1e91f65051300009517b9d1, /*  430 */
128'h078484930000a4970807d7830000a797, /*  431 */
128'h06a7d7830000a7970285d703ecf711e3, /*  432 */
128'h016589930205891320000793eaf719e3, /*  433 */
128'h46192a5050ef854a85ce461900f59a23, /*  434 */
128'h4619295050ef854e028585930000a597, /*  435 */
128'h283050ef00640513018585930000a597, /*  436 */
128'h061301c45783279050ef852285ca4619, /*  437 */
128'hd78302f4142301e4578302f4132302a0, /*  438 */
128'h079300f41f230024d78300f41e230004, /*  439 */
128'h05130000951785aab36900f416236080, /*  440 */
128'hb603300017b7bba546013cf030ef17e5, /*  441 */
128'h00f674132601608130239f0101138307, /*  442 */
128'h879b0387f5930034179b66858387b703, /*  443 */
128'h5e913c23639c97ae300005b79fad8406, /*  444 */
128'h849b5f200513fee7881b278160113423, /*  445 */
128'h00c5163b101005138a1d09056c63ffc7, /*  446 */
128'h07130000a717c34927018f71fff74713, /*  447 */
128'h871b700776130084171beb3d4318f4e7, /*  448 */
128'h969b00d100a345d495ba070e9f318006, /*  449 */
128'h550300d100230086d69b0106d69b0106, /*  450 */
128'h1e63806686936685c6918005069b0001, /*  451 */
128'h30000837860a27850077e79337ed02d5, /*  452 */
128'h983a00369813974285b246814037d79b, /*  453 */
128'h0006881bff063c230621068500083803, /*  454 */
128'h300017b70405a9bff0ef8626fef845e3, /*  455 */
128'h3483852660013403608130838287b823, /*  456 */
128'he8220c2007b711018082610101135f81, /*  457 */
128'hb703300014b747812401ec06e42643c0, /*  458 */
128'h00009517e7990206c163033716938304, /*  459 */
128'h60e2c3c00c2007b729d030ef06450513, /*  460 */
128'hbfc14785ec3ff0ef8082610564a26442, /*  461 */
128'h0000a597461184ae8432ec26f0227179, /*  462 */
128'h0000a7970d7050eff4060068e8458593, /*  463 */
128'ha89785a6862247b20007a803e3c78793, /*  464 */
128'h0693e26757030000a717e22888930000, /*  465 */
128'h85228e0ff0efe2e505130000a5170450, /*  466 */
128'h05220085579b8082614564e2740270a2, /*  467 */
128'h0185579b0185171b8082914115428d5d, /*  468 */
128'h8fd98f750085571bf00686938fd966c1, /*  469 */
128'h808225018d5d8d7900ff07370085151b, /*  470 */
128'h4585460100740207879b070007b7715d, /*  471 */
128'hf052f44ef84afc26e0a2e48604b00513, /*  472 */
128'h0513000095178a2a047070efc63eec56, /*  473 */
128'h89930000a9975ae144011bf030eff9e5, /*  474 */
128'h028a863b4499f969091300009917da69, /*  475 */
128'h0286061b0405854a0004059b013407b3, /*  476 */
128'h185030ef00c780230ff6761300ca5633, /*  477 */
128'h0048d6c585930000a5974611fc941ee3, /*  478 */
128'h0028d5a585930000a59746097de050ef, /*  479 */
128'h010006374722f43ff0ef45127ce050ef, /*  480 */
128'h0ff777138ff183210087179bf0060613, /*  481 */
128'h80a6b02317c29101300016b78fd91502, /*  482 */
128'h60a68086b7838006b78380f6b42393c1, /*  483 */
128'h7a0279a2794274e282f6b42347a16406, /*  484 */
128'hb5838007b603300017b7808261616ae2, /*  485 */
128'hfc068f4d91c115c20080073771398087, /*  486 */
128'hb423e05ae456e852ec4ef04af426f822, /*  487 */
128'ha7170d7030efede505130000951780e7, /*  488 */
128'ha817cbe7c7830000a797cc5747030000, /*  489 */
128'ha617cac6c6830000a697cb7848030000, /*  490 */
128'h9517c9a5c5830000a597ca3646030000, /*  491 */
128'h04130000a41709b030efeb2505130000, /*  492 */
128'hc60989930000a997448100044783c864, /*  493 */
128'h0000aa1700144783c6f70c230000a717, /*  494 */
128'h4783c6f701a30000a7176a89c54a0a13, /*  495 */
128'h08230000a7173000193700262b370024, /*  496 */
128'h4783c4f702a30000a71700344783c4f7, /*  497 */
128'ha71700544783c2f70d230000a7170044, /*  498 */
128'ha797c00793230000a797c2f707a30000, /*  499 */
128'ha797c007a1230000a797be07ad230000, /*  500 */
128'he4a9be07a5230000a797be07ab230000, /*  501 */
128'h5a0b0493f23fe0ef8522e78d0009a783, /*  502 */
128'h83093783020745630337971383093783, /*  503 */
128'h2783bfc5c13ff0effc075de303379713, /*  504 */
128'h710a84937c9050ef4501dff154fd000a, /*  505 */
128'h00154783b7d914fdb7e9bf9ff0efbfc1, /*  506 */
128'h00354503002547838f5d07a200054703, /*  507 */
128'h871b4781808225018d5d05628fd907c2, /*  508 */
128'h0007468300f58733808200e613630007, /*  509 */
128'h079b9e29b7d500d70023078500f50733, /*  510 */
128'hbfc5feb50fa30505808200f613630005, /*  511 */
128'h00958413e04ae426ec06e8221101495c, /*  512 */
128'h4821451502000613478101853903cfb5, /*  513 */
128'h00630007470300f9073346ad02e00893, /*  514 */
128'h15630007831b0e50071300a7146302c7, /*  515 */
128'h0785040500e400230405011400230103, /*  516 */
128'h842384ae01c9051300b94783fcd79be3, /*  517 */
128'h0189470301994783c088f4bff0ef00f5, /*  518 */
128'h47030179478300f492238fd90087979b, /*  519 */
128'h0004002300f493238fd90087979b0169, /*  520 */
128'h873e611c80826105690264a2644260e2, /*  521 */
128'hfc630007468303a0061302000593cf99, /*  522 */
128'h577d00d706630017869300c6986302d5, /*  523 */
128'h869b577d46050007c683b7dd0705a00d, /*  524 */
128'h0006871b078900b666630ff6f593fd06, /*  525 */
128'hbfd5aa2747030000a7178082853ae11c, /*  526 */
128'h0067d683c70d0007c703cb85611cc915, /*  527 */
128'h0017c503e406114102e6906300855703, /*  528 */
128'h60a24525c391450100157793402060ef, /*  529 */
128'h01a5c68301b5c7838082452580820141, /*  530 */
128'h00e51d630006879b8edd0087979b470d, /*  531 */
128'h979b8fd10087179b0145c6030155c703, /*  532 */
128'hec26f02271798082853e27818fd50107, /*  533 */
128'h842a03450993e052e84af4065904e44e, /*  534 */
128'h2501390060ef85ce8626468500154503, /*  535 */
128'heb6340f487bb000402234c58505ce131, /*  536 */
128'h6a0269a2694264e2740270a2450100e7, /*  537 */
128'h4c5cff2a74e34a050034490380826145, /*  538 */
128'h34e060ef85ce86269cbd468500144503, /*  539 */
128'hf06fc39900454783b7f94505b7e5397d, /*  540 */
128'he426ec06e8221101591c80824501f8df, /*  541 */
128'hfddff0ef892e84aa02b787634401e04a, /*  542 */
128'h8593864a46850014c503ec190005041b, /*  543 */
128'ha823597d4405c11925012d6060ef0344, /*  544 */
128'h80826105690264a2644260e285220324, /*  545 */
128'h0005022357fde04ae426ec06e8221101, /*  546 */
128'h23344783e52d2501fa3ff0ef842ad91c, /*  547 */
128'h0107979b8fd90087979b450923244703, /*  548 */
128'h051302e79f63a55707134107d79b776d, /*  549 */
128'h0913010005370005079bd4bff0ef06a4, /*  550 */
128'h45010127f7b31465049300544537fff5, /*  551 */
128'h75332501d25ff0ef0864051300978c63, /*  552 */
128'h690264a2644260e200a035338d050125, /*  553 */
128'he486f44ef84a715dbfcd450d80826105, /*  554 */
128'h852e89aa00053023ec56f052fc26e0a2, /*  555 */
128'h0035171302054e6347adddbff0ef8932, /*  556 */
128'h47b184aa638097ba8a8787930000a797, /*  557 */
128'h00144503c79d000447830089b023c015, /*  558 */
128'h891100090563e38500157793222060ef, /*  559 */
128'h7a0279a2794274e2640660a647a9c111, /*  560 */
128'h000400230ff4f51380826161853e6ae2, /*  561 */
128'hfb79478d00157713136060ef00a400a3, /*  562 */
128'hee5ff0ef85224581f571891100090463, /*  563 */
128'h23a40a131fa40913848a04f51a634785, /*  564 */
128'hc51ff0ef854ac7894501ffc9478389a6, /*  565 */
128'h8913ff2a14e30991094100a9a0232501, /*  566 */
128'h852285d2000a076345090004aa030104, /*  567 */
128'h4785470dfe9915e30491c10dea1ff0ef, /*  568 */
128'h4a01f6e505e34785470dbf8500e51963, /*  569 */
128'h979b03f4470304044783b78547b5c119, /*  570 */
128'h200007134107d79b0107979b8fd90087, /*  571 */
128'h0089999b04a4478304b44983fee791e3, /*  572 */
128'h2e230444448329811a09876300f9e9b3, /*  573 */
128'h0ff7f793009401a3fff4879b47050134, /*  574 */
128'hfa0903e30124012304144903faf769e3, /*  575 */
128'h04644a83ffc100f977b3fff9079b2901, /*  576 */
128'h0154142300faeab3008a9a9b04544783, /*  577 */
128'h151b0474478304844503ffbd00faf793, /*  578 */
128'h042447030434478314050e638d5d0085, /*  579 */
128'h2781033486bbdfa98fd90087979b2501, /*  580 */
128'hf4c563e3873200d7063b9f3d004ad71b, /*  581 */
128'h6605f3266ce384ae032655bb40c5063b, /*  582 */
128'h00b939331955694100b6776349051655, /*  583 */
128'hcc04d458014787bb24890147073b0909, /*  584 */
128'hf00a93e310e91163470dd05c03442023, /*  585 */
128'h849b0024949bd408b09ff0ef06040513, /*  586 */
128'hc45cc81c57fdee99e6e30094d49b1ff4, /*  587 */
128'h478308f91963478d00f402a3f8000793, /*  588 */
128'h0107979b8fd90087979b064447030654, /*  589 */
128'h8522001a059b06e79b6347054107d79b, /*  590 */
128'h2324470323344783e13d2501ce7ff0ef, /*  591 */
128'h776d0107979b8fd90087979b000402a3, /*  592 */
128'h0344051304e79263a55707134107d79b, /*  593 */
128'h1763252787932501416157b7a8dff0ef, /*  594 */
128'h2501614177b7a77ff0ef2184051302f5, /*  595 */
128'ha61ff0ef21c4051300f51c6327278793, /*  596 */
128'h00009797c448a57ff0ef22040513c808, /*  597 */
128'h10230000971793c117c2278562e7d783, /*  598 */
128'h478100042a230124002300f4132362f7, /*  599 */
128'hb5b10005099ba27ff0ef05840513b351, /*  600 */
128'h9fb5e00a84e3b545a19ff0ef05440513, /*  601 */
128'h478db7090014949b00f915634789d41c, /*  602 */
128'h1101bdcd9cbd0017d79b8885029787bb, /*  603 */
128'hed692501c01ff0ef842ae426ec06e822, /*  604 */
128'h4785005447030cf71063478d00044703, /*  605 */
128'h8526458120000613034404930af71b63, /*  606 */
128'hfaa0079322f40923055007939fdff0ef, /*  607 */
128'h02f40aa302f40a230520079322f409a3, /*  608 */
128'h0713481c20f40da302f40b2306100793, /*  609 */
128'h571b0107971b20e40d2302e40ba30410, /*  610 */
128'hd71b20e40ea320f40e230087571b0107, /*  611 */
128'h20e40f23445c20f40fa30187d79b0107, /*  612 */
128'h45030087571b0107571b0107971b5010, /*  613 */
128'h260522e400a322f40023072006930014, /*  614 */
128'h20d40ca320d40c230187d79b0107d71b, /*  615 */
128'h50ef85a64685d81022f401a322e40123, /*  616 */
128'h50ef4581460100144503000402a367d0, /*  617 */
128'h610564a2644260e200a0353325016710, /*  618 */
128'h00e7f963377985beffe5879b4d188082, /*  619 */
128'h450180829d3d02b787bb554800254783, /*  620 */
128'hf406e84a71794d180eb7f56347858082, /*  621 */
128'h0005470302e5f963892ae44eec26f022, /*  622 */
128'h1e6308d70d63468d06d70b63842e4689, /*  623 */
128'h9dbd0094d59b9cad515c0015d49b00f7, /*  624 */
128'h64e2740270a257fdc9112501ac7ff0ef, /*  625 */
128'h899b0249278380826145853e69a26942, /*  626 */
128'h854a9dbd94ca1ff4f4930099d59b0014, /*  627 */
128'h1ff9f993f5792501a93ff0ef0344c483, /*  628 */
128'hc0198fc50087979b880503494783994e, /*  629 */
128'h0085d59b515cbf4d93d117d2bf658391, /*  630 */
128'h74130014141bf1452501a65ff0ef9dbd, /*  631 */
128'h0087979b034945030359478399221fe4, /*  632 */
128'ha3bff0ef9dbd0075d59b515cb7618fc9, /*  633 */
128'h034505131fc575130024151bf93d2501, /*  634 */
128'h4785bfb9024557931512ffaff0ef954a, /*  635 */
128'hf822fc06f04a4544f42671398082853e, /*  636 */
128'h9c63892a478500b51523e456e852ec4e, /*  637 */
128'h6a4269e2790274a2744270e2450900f4, /*  638 */
128'h842efee4f4e34f98611c808261216aa2, /*  639 */
128'heb0d579800e69463470d0007c683e0a9, /*  640 */
128'hd171009928235788fce477e30087d703, /*  641 */
128'h883d0009378300f92a239fa90044579b, /*  642 */
128'hb75d450100893c23943e034787930416, /*  643 */
128'h0009350309924a855a7d0027c98384ba, /*  644 */
128'hf0efbf7d2501e5dff0ef0134766385a6, /*  645 */
128'h3783f69afce301448c630005049be75f, /*  646 */
128'h4505bfc14134043bf6f4f7e34f9c0009, /*  647 */
128'h842aec06e426e822110100a55583b795, /*  648 */
128'hf0ef6008484ce4950005049bf35ff0ef, /*  649 */
128'h4581020006136c08ec990005049b939f, /*  650 */
128'h4705601c00e7802357156c1cf3cff0ef, /*  651 */
128'h8082610564a28526644260e200e78223, /*  652 */
128'he456f04af426f822fc06e852ec4e7139, /*  653 */
128'hf0634a0984aa4d1c0ab9f5634a094985, /*  654 */
128'h0ae78f63842e89324709000547830af5, /*  655 */
128'h515c0015d99b093794630ee78863470d, /*  656 */
128'h0a1b8bdff0ef9dbd0099d59b00b989bb, /*  657 */
128'h0ff9779300198a9b8805060a16630005, /*  658 */
128'h66850347c783013487b3cc191ff9f993, /*  659 */
128'hf7938fd98ff50049179b00f7f71316c1, /*  660 */
128'h50dc00f48223478502f98a2399a60ff7, /*  661 */
128'h00050a1b86fff0ef9dbd8526009ad59b, /*  662 */
128'h79130049591bc40d1ffafa93000a1f63, /*  663 */
128'h70e200f482234785032a8a239aa60ff9, /*  664 */
128'h61216aa26a4269e2790274a285527442, /*  665 */
128'h79130089591b0347c783015487b38082, /*  666 */
128'h0085d59b515cb7e90127e9339bc100f9, /*  667 */
128'h141bfc0a12e300050a1b815ff0ef9dbd, /*  668 */
128'h0109191b03240a2394261fe474130014, /*  669 */
128'h0134822303240aa30089591b0109591b, /*  670 */
128'h0a1bfdcff0ef9dbd0075d59b515cbf79, /*  671 */
128'h0a931fc474130024141bf80a16e30005, /*  672 */
128'hf00006372501d96ff0ef85569aa60344, /*  673 */
128'hd79b94260109179b2901012569338d71, /*  674 */
128'h579b00fa80a30087d79b03240a230107, /*  675 */
128'hbf79012a81a300fa81230189591b0109, /*  676 */
128'he456e852f04af822fc06ec4ef4267139, /*  677 */
128'h4d1c0009056300c52903e99189ae84aa, /*  678 */
128'h0005041bc5bff0efa815490502f96d63, /*  679 */
128'h74a2744270e2852244050087ed634785, /*  680 */
128'h026357fd808261216aa26a4269e27902, /*  681 */
128'h5afd4a05844afef461e3894e4c9c08f4, /*  682 */
128'hb7e94401012a646300f4676324054c9c, /*  683 */
128'h0a63c9012501c0dff0ef852685a24409, /*  684 */
128'h10000637b7cdfd241de3fb450ae30555, /*  685 */
128'h9063e9052501debff0ef852685a2167d, /*  686 */
128'hc89c37fdf8e788e3577dc4c0489c0209, /*  687 */
128'h8622bfb500f482a30017e7930054c783, /*  688 */
128'h14e34785dd612501dbdff0ef852685ce, /*  689 */
128'hfc0600a55903f04a7139b795547df6f5, /*  690 */
128'he456e852ec4ef426030917932905f822, /*  691 */
128'h69e2790274a2744270e24511eb9993c1, /*  692 */
128'h00f97993d7ed495c808261216aa26a42, /*  693 */
128'hc85c61082785480c00099d63842a8a2e, /*  694 */
128'h601cfcf775e30009071b00855783e18d, /*  695 */
128'h4501ec1c97ce03478793012415230996, /*  696 */
128'h0157fab337fd00495a9b00254783bf5d, /*  697 */
128'he46347850005049bb2fff0effc0a9fe3, /*  698 */
128'hb761450500f4946357fdbf4945090097, /*  699 */
128'hf0ef480cf60a0ee306f4e0634d1c6008, /*  700 */
128'hfcf48be34785d4bd451d0005049be83f, /*  701 */
128'hf5792501de0ff0ef6008fcf48de357fd, /*  702 */
128'hbf0ff0ef034505134581200006136008, /*  703 */
128'h02aa2823aabff0ef855285a600043a03, /*  704 */
128'h87bb591c00faed630025478360084a05, /*  705 */
128'hc848a89ff0ef85a6c8046008d91c4157, /*  706 */
128'h6018f1412501d24ff0ef01450223b7b9, /*  707 */
128'hf426f8227139b7e9db1c27855b1c2a85, /*  708 */
128'h0005c783e05ae456e852ec4ef04afc06, /*  709 */
128'h05c0071300e78663842e84aa02f00713, /*  710 */
128'h47fd000447030004a62304050ce79463, /*  711 */
128'h02e0099305c00a9302f00a130ce7f063, /*  712 */
128'hb9030d5784630d478663000447834b21, /*  713 */
128'h4783b42ff0ef854a02000593462d0204, /*  714 */
128'h946300144783013900230d3796630004, /*  715 */
128'h89630024478300f900a302e007930b37, /*  716 */
128'h05a302000793943a09479b63470d1d37, /*  717 */
128'h100519632501adfff0ef8526458100f9, /*  718 */
128'h100511632501ce0ff0ef608848cc492d, /*  719 */
128'h8ba100b7478312078063000747836c98, /*  720 */
128'hc68300f58633078500f706b3708cef89, /*  721 */
128'hf0ef852645810cd60a63fff646030006, /*  722 */
128'hbf35c55c4bdc611ca0e1dd5d2501df9f, /*  723 */
128'h70e20004bc232501a81ff0ef85264581, /*  724 */
128'h61216b026aa26a4269e2790274a27442, /*  725 */
128'h0693f75787e3b7b54709b73d04058082, /*  726 */
128'h4681b78d02400793943a12f6e7630200, /*  727 */
128'h0505a8c948e502000313478145a14701, /*  728 */
128'h0023954a9101020695130027e793a211, /*  729 */
128'h94320200051392011602a865268500e5, /*  730 */
128'h071300094683c6e5460100e573634611, /*  731 */
128'h01659f6300e90023471500e695630e50, /*  732 */
128'h00e7946347118bb10ff7f7930027979b, /*  733 */
128'h46850037f713bded00c905a300866613, /*  734 */
128'h709cf1279de3b7c501066613fed714e3, /*  735 */
128'h0047f713f4e513e34711c51500b7c783, /*  736 */
128'h0ae30004bc230004a623cb990207f793, /*  737 */
128'hb7054515f315bfd94511b72d4501e607, /*  738 */
128'h609cdbe58bc100b5c7836c8cfbe58b91, /*  739 */
128'h05659a63b5a1c4c8ae4ff0ef0007c503, /*  740 */
128'h061b873245ad46a10ff7f7930027979b, /*  741 */
128'hf2e37de3000747039722930117020017, /*  742 */
128'h02b6f263fd370ae3f35709e3f3470be3, /*  743 */
128'h0000851700054c634185551b0187151b, /*  744 */
128'hef0719e30008066300054803f1450513, /*  745 */
128'heea8f3e30ff57513fbf7051bb5754519, /*  746 */
128'he7933701eca8efe30ff57513f9f7051b, /*  747 */
128'he84aec26f0227179bdc10ff777130017, /*  748 */
128'h49bd0e500913451184aef406842ae44e, /*  749 */
128'h2501aecff0ef6008a0b1c90de199484c, /*  750 */
128'hf79300b7c783c3210007c7036c1ce129, /*  751 */
128'hb79317e18bfd033780630327026303f7, /*  752 */
128'h694264e2740270a2450100979a630017, /*  753 */
128'h2501bfdff0ef852245818082614569a2, /*  754 */
128'h45811101bfe54511b7cd00042a23d945, /*  755 */
128'he50d250187dff0ef842ae426ec06e822, /*  756 */
128'hed092501a7eff0ef6008484c0e500493, /*  757 */
128'h85224585cb9900978d630007c7836c1c, /*  758 */
128'h451d00f513634791dd792501bb7ff0ef, /*  759 */
128'he426e82211018082610564a2644260e2, /*  760 */
128'h484ce49d0005049bfa9ff0ef842aec06, /*  761 */
128'h06136c08e0850005049ba34ff0ef6008, /*  762 */
128'hf0ef462d6c08700c838ff0ef45810200, /*  763 */
128'h8526644260e200e782234705601c80ef, /*  764 */
128'h71794d1c08b7f06347858082610564a2, /*  765 */
128'h892e842ae052e44eec26f406e84af022, /*  766 */
128'hed6ff0ef852285ca59fd4a0506f5f063, /*  767 */
128'h694264e2740270a24501e8910005049b, /*  768 */
128'h03348c6303448c63808261456a0269a2, /*  769 */
128'h481cfd7125018abff0ef852285ca4601, /*  770 */
128'h0017e79300544783c81c278501378a63, /*  771 */
128'hbf65faf4e7e30004891b4c1c00f402a3, /*  772 */
128'hec2a713980824509bf4d4505bf5d4509, /*  773 */
128'h4263832ff0eff42ee432e82efc061028, /*  774 */
128'h00a78733050eb0678793000097970405, /*  775 */
128'h0023c319676200070023c31966226318, /*  776 */
128'h00f618634785cb114501e39897aa0007, /*  777 */
128'h612170e22501a02ff0ef0828080c4601, /*  778 */
128'hf8cafca6e122e5067175bfe5452d8082, /*  779 */
128'h0005302316050c63e42eecd6f0d2f4ce, /*  780 */
128'h25019ceff0ef1028002c8a7984aa8932, /*  781 */
128'h2501b61ff0efe4be1028083c65a2e91d, /*  782 */
128'h01f9799301c977934519e011e1196406, /*  783 */
128'hf0ef102800f517634791c11510078e63, /*  784 */
128'h79a6794674e6640a60aac9052501e7df, /*  785 */
128'h8bc5451d00b44783808261496ae67a06, /*  786 */
128'h0a6300897913fff9452100497793f3fd, /*  787 */
128'h046007937a220089e9936406a0210809, /*  788 */
128'h0004072300f40ca300f408a302100713, /*  789 */
128'h00040ba300040b2300e40823000407a3, /*  790 */
128'h00040ea300040e23000405a300e40c23, /*  791 */
128'he0ef85a2000a450300040fa300040f23, /*  792 */
128'h00040a2300040da300040d234785f9bf, /*  793 */
128'h0209036300fa02230005091b00040aa3, /*  794 */
128'hfd212501e1fff0ef030a2a83855285ca, /*  795 */
128'h250180cff0ef0125262385d6397d7522, /*  796 */
128'h85a279220209e993c3990089f793f139, /*  797 */
128'h000485a3d09c01348523f48003092783, /*  798 */
128'he0ef01c40513c8c8f35fe0ef00094503, /*  799 */
128'h0004ae230004a623c88800695783daff, /*  800 */
128'hee051de3bdf5450100f494230124b023, /*  801 */
128'h7913ee0716e30107f713451100b44783, /*  802 */
128'hbf51ec079ee3451d8b85fa0900e30029, /*  803 */
128'hfc86e4d6e8d2eccef8a27119bdd14525, /*  804 */
128'hec6ef06af466f862fc5ee0daf0caf4a6, /*  805 */
128'he85fe0ef8ab6e4328a2e842a0006a023, /*  806 */
128'hc39d662200b44783000998630005099b, /*  807 */
128'h69e6790674a6854e744670e60007899b, /*  808 */
128'h6de27d027ca27c427be26b066aa66a46, /*  809 */
128'h290316078c638b8500a4478380826109, /*  810 */
128'h091b00f67463893e40f907bb445c0104, /*  811 */
128'h5cfd03040b131ff00c1320000b930006, /*  812 */
128'h6008120791631ff777934458fa090ae3, /*  813 */
128'h7d1301a7fd3337fd0025478300975d1b, /*  814 */
128'h00a7ec6347854848eb11020d19630ffd, /*  815 */
128'hbc6ff0ef4c0cbfb5498900f405a34789, /*  816 */
128'h498500f405a3478501951763b7e52501, /*  817 */
128'hb86ff0efe43e853e4c0c601ccc08b795, /*  818 */
128'h67a28dc200a6083b000d061bd5792501, /*  819 */
128'h00c4873b0099549b0027c683072c7a63, /*  820 */
128'h864286a60017c50341a684bb00e6f463, /*  821 */
128'hf79300a44783f9452501176050ef85d2, /*  822 */
128'h951b0097fc6341b507bb4c48c3850407, /*  823 */
128'he0ef955285da20000613910115020097, /*  824 */
128'h445c9a3e9381020497930094949bc3ff, /*  825 */
128'ha0239fa5000aa783c45c9fa54099093b, /*  826 */
128'h771300a44703050601634c50bf3900fa, /*  827 */
128'h50efe44285da46850017c503c30d0407, /*  828 */
128'hfbf7f793682200a44783f131250113c0, /*  829 */
128'h85da0017c50386424685601c00f40523, /*  830 */
128'h049b444c01b42e23f10d25010e8050ef, /*  831 */
128'h049b0127746340bb873b1ff5f5930009, /*  832 */
128'hbb1fe0ef855295a28626030585930007, /*  833 */
128'he8d2eccef0caf8a27119b585499dbf9d, /*  834 */
128'hf06af466f862fc5ee0daf4a6fc86e4d6, /*  835 */
128'he0ef8ab689328a2e842a0006a023ec6e, /*  836 */
128'hc39d00b44783000997630005099bca3f, /*  837 */
128'h69e6790674a6854e744670e60007899b, /*  838 */
128'h6de27d027ca27c427be26b066aa66a46, /*  839 */
128'h445c1a0782638b8900a4478380826109, /*  840 */
128'h1ff00c1320000b9304f76e630127873b, /*  841 */
128'h1ff777930409046344585cfd03040b13, /*  842 */
128'h37fd0025478300975d1b600814079463, /*  843 */
128'h485cef01040d1a630ffd7d1301a7fd33, /*  844 */
128'h00f405a3478902e798634705cb914581, /*  845 */
128'hf3fd0005079bd6aff0ef4c0cb7494989, /*  846 */
128'h0207e79300a4478312f76b634818445c, /*  847 */
128'h00f405a3478501979763b78500f40523, /*  848 */
128'h00a44783c85ce311cc1c4858bf894985, /*  849 */
128'h0017c50346854c50601cc38d0407f793, /*  850 */
128'hf79300a44783f96925017d9040ef85da, /*  851 */
128'hf0efe43e853e4c0c601c00f40523fbf7, /*  852 */
128'h8db200a8063b000d081bd1592501964f, /*  853 */
128'h873b0099549b0027c683072c7a6367a2, /*  854 */
128'h86a60017c50341a684bb00e6f4630104, /*  855 */
128'h41b587bb4c4cf1492501789040ef85d2, /*  856 */
128'h20000613918115820097959b0297f263, /*  857 */
128'hfbf7f79300a44783a29fe0ef855a95d2, /*  858 */
128'h9a3e9381020497930094949b00f40523, /*  859 */
128'h9fa5000aa783c45c9fa54099093b445c, /*  860 */
128'h4458481400c70e634c58bdc900faa023, /*  861 */
128'h6ed040ef85da46850017c50300d77a63, /*  862 */
128'h75130009049b444801b42e23fd012501, /*  863 */
128'h05130007049b0127746340ab873b1ff5, /*  864 */
128'h00a447839b5fe0ef952285d286260305, /*  865 */
128'h499db5f1c81cbf4100f405230407e793, /*  866 */
128'h2501ab7fe0ef842ae406e0221141bd15, /*  867 */
128'h0407f793cf610207f71300a44783e16d, /*  868 */
128'h030405930017c50346854c50601cc395, /*  869 */
128'hfbf7f79300a44783ed4d25016ab040ef, /*  870 */
128'he1552501b5ffe0ef6008500c00f40523, /*  871 */
128'h481800e785a30207671300b7c703741c, /*  872 */
128'h00e78e230086d69b0106d69b0107169b, /*  873 */
128'h00d78f230187571b0107569b00d78ea3, /*  874 */
128'h8d2300078ba300078b23485800e78fa3, /*  875 */
128'h171b00e78a230107571b0107169b00e7, /*  876 */
128'hd69b00e78aa30087571b0107571b0107, /*  877 */
128'h07130086d69b00e78c23021007130106, /*  878 */
128'h89a30007892300e78ca300d78da30460, /*  879 */
128'h00f40523fdf7f793600800a447830007, /*  880 */
128'hea3fe06f014160a2640200f502234785, /*  881 */
128'he406e022114180820141640260a24505, /*  882 */
128'h9b5fe0ef8522e9012501f01ff0ef842a, /*  883 */
128'h80820141640260a200043023e1192501, /*  884 */
128'h00054a63945fe0efec060028e42a1101, /*  885 */
128'h8082610560e2450142a7842300008797, /*  886 */
128'hf0a21028002c4601e42a7159bfe5452d, /*  887 */
128'h65a2ec190005041bb25fe0efeca6f486, /*  888 */
128'he41d0005041bcb4ff0efe4be1028083c, /*  889 */
128'h740670a68522cbd8575277a2e9916586, /*  890 */
128'h74a2cb998bc100b5c7838082616564e6, /*  891 */
128'h1ee34791b7c5c8c8965fe0ef0004c503, /*  892 */
128'he122e506e42afca67175bfd94415fcf4, /*  893 */
128'h1828002c460184ae00050023f4cef8ca, /*  894 */
128'h842677e2ecbe081ce5212501ab9fe0ef, /*  895 */
128'h4501040991634996c2be4bdc02f00913, /*  896 */
128'h0307071b3747470300008717e50567a2, /*  897 */
128'h0e94156300e780a303a0071300e78023, /*  898 */
128'h60aa00078023078d00e7812302f00713, /*  899 */
128'h182845858082614979a6794674e6640a, /*  900 */
128'he6cff0ef18284581fd4d2501f75fe0ef, /*  901 */
128'h8bdfe0ef0007c50365c677e2f55d2501, /*  902 */
128'h4581f9512501f4ffe0ef18284581c2aa, /*  903 */
128'hc50365c677e2e1052501e46ff0ef1828, /*  904 */
128'h1828458101350e632501897fe0ef0007, /*  905 */
128'hf6e512e367a24711dd612501a86ff0ef, /*  906 */
128'h97134781f48fe0ef1828100cb7614509, /*  907 */
128'h871be705fc9747039736109493010207, /*  908 */
128'h9713662236fd86a285be04e460630037, /*  909 */
128'h01260023fff7c793e989963a93010206, /*  910 */
128'h0007059bfff5871bb7e12785bf199c3d, /*  911 */
128'h00e60023fc974703972a108893011702, /*  912 */
128'h92810204169367220789bdf54545b7e9, /*  913 */
128'h65e3fee78fa324050785000747039736, /*  914 */
128'hec4efc06f04af426f8227139b721fe94, /*  915 */
128'h0005091bfa8fe0ef84ae842ae456e852, /*  916 */
128'h70e20007891bcf8900b4478300091763, /*  917 */
128'h61216aa26a4269e2790274a2854a7442, /*  918 */
128'he3918b8900a447830097776348188082, /*  919 */
128'h78e34818445ce4bd00042623445884ba, /*  920 */
128'h00f405230207e79300a44783c81cfcf7, /*  921 */
128'h0ee34c50d3e51ff7f793445c4481bf7d, /*  922 */
128'hc3850407f7930304099300a44783fc96, /*  923 */
128'h2501341040ef0017c50385ce4685601c, /*  924 */
128'h601c00f40523fbf7f79300a44783ed51, /*  925 */
128'h25012ef040ef85ce0017c50386264685, /*  926 */
128'h0097999b002547836008bf59cc44ed35, /*  927 */
128'h0337563b0336d6bbfff4869b377dc729, /*  928 */
128'hc45c27814c0c8ff9413007bb02c6ed63, /*  929 */
128'h9fa5445c0499ea634a855a7dd1c19c9d, /*  930 */
128'h2501c79fe0ef6008d7b51ff4f793c45c, /*  931 */
128'hf0efe595484cbfb19ca90094d49bcd11, /*  932 */
128'h05a3478900f5976347850005059b802f, /*  933 */
128'h05a3478500f5976357fdbded490900f4, /*  934 */
128'h00a44783b765cc0cc84cb5ed490500f4, /*  935 */
128'he5990005059bfcbfe0efcb818b896008, /*  936 */
128'hfd4588e30005059bc3ffe0efbf6984ce, /*  937 */
128'hcc0c445cfaf5fae34f9c601cfabafee3, /*  938 */
128'hfc067139b7bdc45c013787bb413484bb, /*  939 */
128'he0ef0828002c4601842ac52de42ef822, /*  940 */
128'h101ce01c852265a267e2e1152501fdaf, /*  941 */
128'hc783cd996c0ce5292501968ff0eff01c, /*  942 */
128'h67e2a02d000430234515e7898bc100b5, /*  943 */
128'h8522458167e2c448e24fe0ef0007c503, /*  944 */
128'h47912501cadfe0ef00f414230067d783, /*  945 */
128'h452580826121744270e2f971fcf50be3, /*  946 */
128'he406e0221141b7c1fcf501e34791bfdd, /*  947 */
128'h60a200043023e1192501daefe0ef842a, /*  948 */
128'hf406e84aec26f0227179808201416402, /*  949 */
128'h1f63e8890005049bd8cfe0ef892e842a, /*  950 */
128'h70a20005049bc4ffe0ef852245810009, /*  951 */
128'h022430238082614564e2694285267402, /*  952 */
128'h02f5136347912501b34ff0ef85224581, /*  953 */
128'h85224581c58fe0ef852285ca00042a23, /*  954 */
128'h00042a2300f5166347912501f77fe0ef, /*  955 */
128'h84aee42aeca67159bf6584aad16dbf7d, /*  956 */
128'h041becefe0eff486f0a21028002c4601, /*  957 */
128'h85eff0efe4be1028083c65a2e00d0005, /*  958 */
128'h102885a6c489cf816786e8010005041b, /*  959 */
128'h8082616564e6740670a68522c00fe0ef, /*  960 */
128'h8b2ee42af85a8432f0a27159bfcd4419, /*  961 */
128'he4cee8caeca6f486e0d28522002c4601, /*  962 */
128'h00050a1be70fe0efec66f062f45efc56, /*  963 */
128'hffec871b481c01842c836000000a1c63, /*  964 */
128'h64e68552740670a600fb202302f76263, /*  965 */
128'h6ce27c027ba27b427ae26a0669a66946, /*  966 */
128'h490902fb9f63478500044b8380826165, /*  967 */
128'h2501a49fe0ef852285ca4a8559fd4481, /*  968 */
128'h29054c1c2485e1110955086309350863, /*  969 */
128'h02a30017e793c80400544783fef963e3, /*  970 */
128'h490110000ab7504cb74d009b202300f4, /*  971 */
128'h899b852200099e631afd4c0944814981, /*  972 */
128'h0344091385cee9212501d04fe0ef0015, /*  973 */
128'h0009470300194783038b916320000993, /*  974 */
128'h3cfd39f909092485e3918fd90087979b, /*  975 */
128'h2501aa2fe0efe02e854ab745fc0c94e3, /*  976 */
128'hb7c539f109112485e111658201557533, /*  977 */
128'he8221101bfad8a2abfbd4a09b7494a05, /*  978 */
128'h0005049bbb8fe0ef842ae04aec06e426, /*  979 */
128'h644260e20007849bcb9100b44783e491, /*  980 */
128'hf71300a447838082610564a269028526, /*  981 */
128'h0207e793fed772e348144458cf390027, /*  982 */
128'ha5aff0ef484cef01600800f40523c818, /*  983 */
128'hbf7d84aa00a405a3c53900042a232501, /*  984 */
128'h02f9146357fd0005091b941fe0ef4c0c, /*  985 */
128'hb25fe0ef167d100006374c0cb7dd4505, /*  986 */
128'hb7e12501a1eff0ef85ca6008f9792501, /*  987 */
128'h4d1c6008fcf900e345094785b769449d, /*  988 */
128'h601cdba50407f79300a44783fcf96ae3, /*  989 */
128'h71e040ef030405930017c50346854c50, /*  990 */
128'h00f40523fbf7f79300a44783f55d2501, /*  991 */
128'he122e5061008002c4605e42a7175b7b1, /*  992 */
128'h081c65a2e9052501c94fe0eff8cafca6, /*  993 */
128'h45196786e1052501e27fe0efe0be1008, /*  994 */
128'hc483c59975e2eb890207f79300b7c783, /*  995 */
128'h74e6640a60aa451dcb810014f79300b5, /*  996 */
128'haccfe0ef000945037902808261497946, /*  997 */
128'h8de301492783c89d88c1cc0d0005041b, /*  998 */
128'h4589952fe0ef00a8100c02800613fc87, /*  999 */
128'h00a84581f1612501941fe0efcaa200a8, /* 1000 */
128'h1008faf518e34791d94d2501838ff0ef, /* 1001 */
128'hf12fe0ef7502e411f15525019e3fe0ef, /* 1002 */
128'hf551250191eff0ef85a27502bf612501, /* 1003 */
128'hf506f1221028002c4605e42a7171b7ed, /* 1004 */
128'hf0e2f4def8dafcd6e152e54ee94aed26, /* 1005 */
128'h1c0412630005041bbc4fe0efe8eaece6, /* 1006 */
128'h0005041bd53fe0efe4be1028083c65a2, /* 1007 */
128'hc783441967a61af4156347911c040763, /* 1008 */
128'he0ef4581752218079d630207f79300b7, /* 1009 */
128'h440975224785180480630005049bb33f, /* 1010 */
128'ha8cfe0ef16f48863440557fd16f48c63, /* 1011 */
128'h0104d91b85a67422160412630005041b, /* 1012 */
128'h45812000061303440b13f60fe0ef8522, /* 1013 */
128'h02000593462d886fe0ef855a00050c1b, /* 1014 */
128'h0104999b0ff97a9347c187afe0ef855a, /* 1015 */
128'h021007930109d99b02f40fa30109191b, /* 1016 */
128'h0ff4fa1304f4062302e00b930109591b, /* 1017 */
128'h04f406a30089591b0089d99b04600793, /* 1018 */
128'h040405a30404052303740a2302000613, /* 1019 */
128'h052404a305540423053407a305440723, /* 1020 */
128'h05740aa37722ff7fd0ef0544051385da, /* 1021 */
128'h9363571400d6166357d200074603468d, /* 1022 */
128'h0107d79b0107969b06f40723478100f6, /* 1023 */
128'h0107d79b0106d69b0107979b06f40423, /* 1024 */
128'h06f404a306d407a30087d79b0086d69b, /* 1025 */
128'hf5ffe0ef1028040b99634c8500274b83, /* 1026 */
128'h00e785a3752247416786e8350005041b, /* 1027 */
128'h00078b230460071300e78c2302100713, /* 1028 */
128'h01378da301478d2300e78ca300078ba3, /* 1029 */
128'he0ef00f50223478501278aa301578a23, /* 1030 */
128'h2823001c0d1b7522a82d0005041bd50f, /* 1031 */
128'hec090005041b8d4fe0ef019502230385, /* 1032 */
128'hfb93f53fd0ef3bfd855a458120000613, /* 1033 */
128'hf2bfe0ef85a67522441db7498c6a0ffb, /* 1034 */
128'h7ae66a0a69aa694a64ea740a70aa8522, /* 1035 */
128'h44218082614d6d466ce67c067ba67b46, /* 1036 */
128'h002c843284aee42aeca6f0a27159b7c5, /* 1037 */
128'h65a2e13125019c2fe0eff48610284605, /* 1038 */
128'h67a6e9152501b55fe0efe4be1028083c, /* 1039 */
128'hc30d6706e39d0207f79300b7c7834519, /* 1040 */
128'h8c3d027474138c658cbd752200b74783, /* 1041 */
128'h2501c94fe0ef00f502234785008705a3, /* 1042 */
128'he02ee42a71718082616564e6740670a6, /* 1043 */
128'h95cfe0efed26f122f5060088002c4605, /* 1044 */
128'hf4be008865a26786120795630005079b, /* 1045 */
128'h100799630005079bae7fe0eff0be083c, /* 1046 */
128'h1007116302077713479900b7c7037786, /* 1047 */
128'hd0ef102805ad46550e058d63479165e6, /* 1048 */
128'h850ae33fd0ef10a8008c02800613e3ff, /* 1049 */
128'he0ef10a865820c054c6347adefdfd0ef, /* 1050 */
128'h10a80ce792634711cbf10005079ba9df, /* 1051 */
128'h0593464d648aebdd0005079bdcbfe0ef, /* 1052 */
128'h640602814783df7fd0ef00d4851302a1, /* 1053 */
128'hc78300f40223478500f485a30207e793, /* 1054 */
128'h450306f7076357d64736cbb58bc100b4, /* 1055 */
128'he0ef85220005059bf25fd0ef85a60004, /* 1056 */
128'hfbbfd0ef8522c1bd47890005059bca4f, /* 1057 */
128'h0557468302e007936706efa90005079b, /* 1058 */
128'hd79b06f707230107969b57d602f69c63, /* 1059 */
128'hd79b0107d79b0107979b06f704230107, /* 1060 */
128'h478506f704a30086d69b0106d69b0087, /* 1061 */
128'h079be18fe0ef008800f7022306d707a3, /* 1062 */
128'h70aa0005079bb48fe0ef6506e7910005, /* 1063 */
128'h711dbfcd47a18082614d853e64ea740a, /* 1064 */
128'he0efec861028002c4605842ee42ae8a2, /* 1065 */
128'he0efe4be1028083c65a2e929250180af, /* 1066 */
128'hf79300b7c783451967a6e129250199df, /* 1067 */
128'h8b23752200645703cb856786eb950207, /* 1068 */
128'h8c230044570300e78ba30087571b00e7, /* 1069 */
128'h00f50223478500e78ca30087571b00e7, /* 1070 */
128'h711d80826125644660e62501acefe0ef, /* 1071 */
128'h08284601002c893284aee42ae0cae4a6, /* 1072 */
128'hc4b9e0510005041bf95fd0efec86e8a2, /* 1073 */
128'h4585e5592501c9efe0efd20208284581, /* 1074 */
128'h8526462d75c2e93d2501b97fe0ef0828, /* 1075 */
128'h00230200061346ad00b48713c8dfd0ef, /* 1076 */
128'h938117820007869bfff6879bce890007, /* 1077 */
128'h02090a63fec783e3177d0007c78397a6, /* 1078 */
128'h6562e0150005041be63fd0ef510c6562, /* 1079 */
128'h079300e684630005468304300793470d, /* 1080 */
128'h00a92023c15fd0ef953e034787930270, /* 1081 */
128'h479180826125690664a6644660e68522, /* 1082 */
128'h711db7d5842abf550004802300f51563, /* 1083 */
128'heddfd0efec86e8a21028002c4605e42a, /* 1084 */
128'h9713478100010c236522e4710005041b, /* 1085 */
128'h02000613eb2900074703972a93010207, /* 1086 */
128'h0005041bbccfe0efda0210284581ebb1, /* 1087 */
128'h100515632501ac3fe0ef10284585e045, /* 1088 */
128'hbb1fd0ef082c462dc7e5650601814783, /* 1089 */
128'h8b230460071300e78c23021007136786, /* 1090 */
128'hb7452785a0e900e78ca300078ba30007, /* 1091 */
128'h96aa928102071693fff7871bb77d87ba, /* 1092 */
128'h06b3432d48e54701fec686e30006c683, /* 1093 */
128'h92c1030596930017061b0006c58300e5, /* 1094 */
128'h36810108ec63030858131842f9f6881b, /* 1095 */
128'h00068e1b92c585930000759792c116c2, /* 1096 */
128'h4419feb045e34185d59b0185959ba831, /* 1097 */
128'h0005c803058580826125644660e68522, /* 1098 */
128'h082cfe6702e3b7ddffc81be300080563, /* 1099 */
128'hf8f6e9e30007069b00d58023070595ba, /* 1100 */
128'h0007869b020006134729938102061793, /* 1101 */
128'hf0f713e30e5007930181470300d77963, /* 1102 */
128'h5795b7c5078500c6802396be0834b77d, /* 1103 */
128'h8b2fe0ef00f502234785752200f50023, /* 1104 */
128'h0181478302f51b634791b7710005041b, /* 1105 */
128'h6506f8350005041ba19fe0ef1028d3c1, /* 1106 */
128'h082c462d6506ab7fd0ef458102000613, /* 1107 */
128'h842abdd100e785a347216786a8dfd0ef, /* 1108 */
128'h28830585230305452e0305052e83bf81, /* 1109 */
128'h040502938f2ae44ae826ec22110105c5, /* 1110 */
128'h488f8f9300005f97887687f2869a8646, /* 1111 */
128'h2583000fa38300b647338dfd00c6c5b3, /* 1112 */
128'ha3839db9007585bb0fc1008fa403000f, /* 1113 */
128'h581b0078159b0105883b004f2703ff4f, /* 1114 */
128'h9f3100f805bb0077073b0105e8330198, /* 1115 */
128'h171b9e39008f23838e358e6d00f6c633, /* 1116 */
128'h00c5873b008383bb8e590146561b00c6, /* 1117 */
128'h8ebd00cf24038ef900b7c6b300d383bb, /* 1118 */
128'h00d3e6b30116969b00f6d39b007686bb, /* 1119 */
128'h8f2d0007061b00d703bbffcfa4039fa1, /* 1120 */
128'h171b00a7579b9f3d8f2d9fa100777733, /* 1121 */
128'h87bb0003869b0005881b0f418f5d0167, /* 1122 */
128'h5f974caf0f1300005f17f45f17e300e3, /* 1123 */
128'hc5b34ca2829300005297402f8f930000, /* 1124 */
128'h001f4383000fa58300b6c7338df100d7, /* 1125 */
128'h070a93aa038a000f47039db9002f4403, /* 1126 */
128'h883b004fa7039db9942a040a4318972a, /* 1127 */
128'h0003a70301b8581b9e390058159b0105, /* 1128 */
128'h8e7500b7c6339f3100f805bb0105e833, /* 1129 */
128'h0176561b0096139b008fa7039e398e3d, /* 1130 */
128'h0f119f3500c583bb00c3e63340189eb9, /* 1131 */
128'h9eb90fc18eadffff44838efd0075c6b3, /* 1132 */
128'hd69b9fb900e6941b94aa048affcfa703, /* 1133 */
128'h0083c7339fb900d3843b8ec140980126, /* 1134 */
128'h0147171b00c7579b9f3d007747338f6d, /* 1135 */
128'h07bb0004069b0003861b0005881b8f5d, /* 1136 */
128'h82fe3eaf8f9300005f97f25f1ee300e4, /* 1137 */
128'h0003a7030102c4033603839300005397, /* 1138 */
128'h9f25400000c5c4b3942a040a00d7c5b3, /* 1139 */
128'h9e2194aa048a0043a4039f210112c483, /* 1140 */
128'h581b0048171b0122c4830107083b4080, /* 1141 */
128'h00f8073b0083a4039e210107683301c8, /* 1142 */
128'h00b6159b40809e2d9ea194aa8db9048a, /* 1143 */
128'h00c705bb03c18e4d0156561b0132c903, /* 1144 */
128'h9ea1090a8ead00e7c6b3ffc3a4839c35, /* 1145 */
128'h000924830106d69b9fa50106941b992a, /* 1146 */
128'h8f219fa58f2d0007081b00d5843b8ec1, /* 1147 */
128'h861b02918f5d0177171b0097579b9f3d, /* 1148 */
128'h5297f45f17e300e407bb0004069b0005, /* 1149 */
128'h00d745b38f5dfff647132e2282930000, /* 1150 */
128'hc5839f2d022fc403021fc3830002a703, /* 1151 */
128'h942a040a418c95aa058a93aa038a020f, /* 1152 */
128'h9e2d0068171b0107083b0042a5839f2d, /* 1153 */
128'h00f8073b0107683301a8581b0003a583, /* 1154 */
128'h0082a5839e2d8e3d8e59fff6c6139db1, /* 1155 */
128'h00c3e633400c9ead0166561b00a6139b, /* 1156 */
128'he5b3fff7c593023fc4839ead00c703bb, /* 1157 */
128'h969b048a9db5ffc2a4038db902c10075, /* 1158 */
128'h85bb40809fa18dd50115d59b94aa00f5, /* 1159 */
128'h47339fa18f4dfff747130007081b00b3, /* 1160 */
128'h0f918f5d0157171b00b7579b9f3d0077, /* 1161 */
128'hf3ff1de300e587bb0005869b0003861b, /* 1162 */
128'h863b00d306bb00fe07bb010e883b6462, /* 1163 */
128'h692264c2cd70cd34c97c0505282300c8, /* 1164 */
128'hf44ef84afc26e0a2715d653c80826105, /* 1165 */
128'h97b203f7f413ec56f052e486e45ee85a, /* 1166 */
128'h04000b9304000b13e53c893289ae84aa, /* 1167 */
128'h00f974639381178200078a1b408b07bb, /* 1168 */
128'h853385ce020ada93020a1a9300090a1b, /* 1169 */
128'h415909334a7020ef0144043b86560084, /* 1170 */
128'hb7c997824401852660bc0174176399d6, /* 1171 */
128'h6b426ae27a0279a2794274e2640660a6, /* 1172 */
128'h03f7f793f0227179653c808261616ba2, /* 1173 */
128'h071300178513e84af406e44eec26842a, /* 1174 */
128'h863b449d0400099300e7802397a2f800, /* 1175 */
128'h20ef95224581920116020006091b40a9, /* 1176 */
128'h8522603cfc1c078e643c0124f5633f30, /* 1177 */
128'h694264e2740270a2fd24fde345019782, /* 1178 */
128'h639cf9a78793000077978082614569a2, /* 1179 */
128'h639cf927879300007797e93c04053423, /* 1180 */
128'h11018082e13cb807879300000797ed3c, /* 1181 */
128'h47013e5020efec06850a464105050593, /* 1182 */
128'h3c858593000065971a06869300007697, /* 1183 */
128'hd613070506890007c78300e107b34541, /* 1184 */
128'h0007c78397ae000646038bbd962e0047, /* 1185 */
128'h751760e2fca71de3fef68fa3fec68f23, /* 1186 */
128'h842ae122717580826105162505130000, /* 1187 */
128'h080885a26622f71ff0efe42ee5060808, /* 1188 */
128'hf83ff0ef0808f01ff0ef0808e85ff0ef, /* 1189 */
128'h0d63711c46a1595880826149640a60aa, /* 1190 */
128'h4501cf980200071300d71763469100d7, /* 1191 */
128'he82211018082556dbfe50007ac238082, /* 1192 */
128'h02f5026384ae842a200007b7ec06e426, /* 1193 */
128'h00006597088006130906869300005697, /* 1194 */
128'h1d3030ef33c505130000651732c58593, /* 1195 */
128'he82211018082610564a2644260e2fc24, /* 1196 */
128'h02f4026384ae200007b7ec06e4266100, /* 1197 */
128'h0000659702f006130686869300005697, /* 1198 */
128'h193030ef2fc50513000065172ec58593, /* 1199 */
128'he82211018082610564a2644260e2e004, /* 1200 */
128'h02f4026384ae200007b7ec06e4266100, /* 1201 */
128'h00006597036006130386869300005697, /* 1202 */
128'h153030ef2bc50513000065172ac58593, /* 1203 */
128'he42611018082610564a2644260e2e404, /* 1204 */
128'h02f48263842e200007b7ec06e8226104, /* 1205 */
128'h0000659703e00613e606869300007697, /* 1206 */
128'h113030ef27c505130000651726c58593, /* 1207 */
128'h8082610564a2644260e2e88090011402, /* 1208 */
128'h842e200007b7ec06e8226104e4261101, /* 1209 */
128'h04500613e14686930000769702f48263, /* 1210 */
128'h23850513000065172285859300006597, /* 1211 */
128'h64a2644260e2ec80900114020cf030ef, /* 1212 */
128'h07b7ec06e4266100e822110180826105, /* 1213 */
128'hf80686930000569702f4026384ae2000, /* 1214 */
128'h000065171e4585930000659704c00613, /* 1215 */
128'h64a2644260e2f00408b030ef1f450513, /* 1216 */
128'h07b7ec06e4266100e822110180826105, /* 1217 */
128'hf50686930000569702f4026384ae2000, /* 1218 */
128'h000065171a4585930000659705300613, /* 1219 */
128'h64a2644260e2f40404b030ef1b450513, /* 1220 */
128'hf426f82200053983ec4e713980826105, /* 1221 */
128'h84638436893284ae200007b7fc06f04a, /* 1222 */
128'h659705a00613f16686930000569702f9, /* 1223 */
128'he43a16a505130000651715a585930000, /* 1224 */
128'h191b8b0588090014141b67227fe030ef, /* 1225 */
128'h012464330034949b8c59004979130029, /* 1226 */
128'h790274a2744270e20289b8238c4588a1, /* 1227 */
128'h468147057100e02211418082612169e2, /* 1228 */
128'h45818522f7dff0efe406458185224605, /* 1229 */
128'hf0ef45814605468547058522f35ff0ef, /* 1230 */
128'h4501640260a2d97ff0ef45816008f67f, /* 1231 */
128'h460546814705e022e406114180820141, /* 1232 */
128'hf39ff0ef842a45810405302302053c23, /* 1233 */
128'h4685470545818522ef1ff0ef45818522, /* 1234 */
128'h0141458160a264026008f23ff0ef4605, /* 1235 */
128'h07b7ec06e8226104e4261101d4dff06f, /* 1236 */
128'he40686930000569702f48263842e2000, /* 1237 */
128'h00006517074585930000659706100613, /* 1238 */
128'h60e2fc809041144271a030ef08450513, /* 1239 */
128'he8226104e42611018082610564a26442, /* 1240 */
128'h0000569702f48263842e200007b7ec06, /* 1241 */
128'h030585930000659706800613e0c68693, /* 1242 */
128'h905114526d6030ef0405051300006517, /* 1243 */
128'he82211018082610564a2644260e2e0a0, /* 1244 */
128'h02f4026384ae200007b7ec06e4266100, /* 1245 */
128'h0000659706f00613dd86869300005697, /* 1246 */
128'h692030efffc5051300006517fec58593, /* 1247 */
128'he04a11018082610564a2644260e2e424, /* 1248 */
128'h842a200007b7ec06e426e82200053903, /* 1249 */
128'h0613da2686930000569702f9026384ae, /* 1250 */
128'h051300006517fa658593000065970760, /* 1251 */
128'h644260e2c84404993c2364c030effb65, /* 1252 */
128'heca67100f0a2715980826105690264a2, /* 1253 */
128'hf062f45ef85afc56e0d2e4cef486e8ca, /* 1254 */
128'he03084b2892e0005d783020408a3ec66, /* 1255 */
128'h9c636f6020ef00c9051345814611d01c, /* 1256 */
128'h07b700043983bf7ff0ef458560080e04, /* 1257 */
128'h44810049278316f99a6304043a032000, /* 1258 */
128'h4c1c4485e391448d8b89c7090017f713, /* 1259 */
128'h8b85008a2783000a09638cdd03243c23, /* 1260 */
128'h45814605468147050144e49316078663, /* 1261 */
128'h2583be3ff0ef85224581d73ff0ef8522, /* 1262 */
128'h00095583c55ff0ef00989a3785220089, /* 1263 */
128'hf0ef852285a6c8bff0ef681a0a138522, /* 1264 */
128'h460546854705cffff0ef85224581cc7f, /* 1265 */
128'h24058593000f45b7d31ff0ef85224581, /* 1266 */
128'hb583cdbff0ef85224585e9bff0ef8522, /* 1267 */
128'h0015e593cccc8c9300005c9785220d89, /* 1268 */
128'h6b17e82a8a9300006a97ebbff0ef2581, /* 1269 */
128'h64e6740670a6efe9485ce92b0b130000, /* 1270 */
128'h6ce27c027ba27b427ae26a0669a66946, /* 1271 */
128'hdb9ff0efe024852244cc808261654501, /* 1272 */
128'hee079be38b85449cdf5ff0ef8522488c, /* 1273 */
128'h458163900107e683654100043883603c, /* 1274 */
128'h6e89f005051300ff0e37431147014781, /* 1275 */
128'h183b070500371f1b00064803ec0689e3, /* 1276 */
128'h0067036316fd060527810107e7b301e8, /* 1277 */
128'h981b010767330187971b0187d81bf2e5, /* 1278 */
128'h8fe9010767330087d79b01c878330087, /* 1279 */
128'h9746938183751782170200be873b8fd9, /* 1280 */
128'h869300005697b765470147812585e31c, /* 1281 */
128'h6517db2585930000659714900613bbe6, /* 1282 */
128'h00c4e493bd85458030efdc2505130000, /* 1283 */
128'h5597000b9d633bfd20000c378bd2bd61, /* 1284 */
128'h00efdb25051300006517ba2585930000, /* 1285 */
128'h061386e60189096300043903b7117020, /* 1286 */
128'h485c07093483418030ef855a85d60f20, /* 1287 */
128'h3783020937031404806324818cfd4981, /* 1288 */
128'hcc5cf9200793c7817c1c00f76f630c89, /* 1289 */
128'hb29ff0ef85224581b71ff0ef85224581, /* 1290 */
128'hff397913852201442903c39d0044f793, /* 1291 */
128'h651785cad45ff0ef85ca290100896913, /* 1292 */
128'hc39d0084f79368a000efd52505130000, /* 1293 */
128'h290100496913ff397913852201442903, /* 1294 */
128'hd50505130000651785cad1bff0ef85ca, /* 1295 */
128'h390300043983cfb50014f793660000ef, /* 1296 */
128'h0613b0a686930000569701898c630384, /* 1297 */
128'h2783cba97c1c368030ef855a85d609c0, /* 1298 */
128'h08e69f630037f693470d02043c230049, /* 1299 */
128'h63104591480d468100c9079301898713, /* 1300 */
128'h370301068763c3900086161bff870513, /* 1301 */
128'h90e30791872a2685c3988f518361ff87, /* 1302 */
128'h485cc85c0027e793485ccbb5603cfeb6, /* 1303 */
128'h040439036004cc9d49858889c85c9bf9, /* 1304 */
128'h0ca00613aa4686930000569701848c63, /* 1305 */
128'h00090963040430232ea030ef855a85d6, /* 1306 */
128'h485cb4bff0ef8522ef8d8b8500892783, /* 1307 */
128'h8ce3c43ff0ef8522484cc85c9bf54985, /* 1308 */
128'hb783dbd98b85bd85677020ef4505d809, /* 1309 */
128'hbf41b1bff0ef8522b77100f926230009, /* 1310 */
128'h8913dcd5010964830009398397a667a1, /* 1311 */
128'h3c2020efe43e002c4621854e639c0087, /* 1312 */
128'h717908b041635535b7dd87ca14e109a1, /* 1313 */
128'h84b2e44ef406e84aec26f02204800513, /* 1314 */
128'h551785a2c41d5551842a1dc030ef892e, /* 1315 */
128'h862285aa89aa7b3010efa12505130000, /* 1316 */
128'h00099d63508000efc205051300006517, /* 1317 */
128'h694264e2740270a2557d1f6030ef8522, /* 1318 */
128'h01242423e01c200007b78082614569a2, /* 1319 */
128'hbfe94501c45c4789c7890024f793f404, /* 1320 */
128'h46098082b7f9c45c4785d8f145018885, /* 1321 */
128'h200007b7050ef73ff06f200005374581, /* 1322 */
128'h6380e0221141711c80822501638897aa, /* 1323 */
128'h86930000569702f40263200007b7e406, /* 1324 */
128'h6517b02585930000659734c006139ae6, /* 1325 */
128'he3914505703c1a8030efb12505130000, /* 1326 */
128'h842ae822110180820141640260a2557d, /* 1327 */
128'h6622644285a2501010efe42eec064501, /* 1328 */
128'h2000051371797a00006f6105468560e2, /* 1329 */
128'h0e2030efe052e44ee84aec26f022f406, /* 1330 */
128'hb5031ea030efb76505130000651784aa, /* 1331 */
128'h10ef842a4bf010ef4501479010ef0001, /* 1332 */
128'h00ef638cb5c5051300006517681c2240, /* 1333 */
128'h00efb5a505130000651706f445834020, /* 1334 */
128'h0085d59bb645051300006517546c3f20, /* 1335 */
128'h651706c4458358303dc000ef91c115c2, /* 1336 */
128'h77930106569b0086571bb5a505130000, /* 1337 */
128'h00ef0186561b0ff6f6930ff777130ff6, /* 1338 */
128'h3a4000efb4c50513000065175c0c3b20, /* 1339 */
128'h00006597c789ad65859300006597545c, /* 1340 */
128'h384000efb3c5051300006517ac458593, /* 1341 */
128'h6597744813c030efb485051300006517, /* 1342 */
128'h584c19c42783e01fb0ef14a585930000, /* 1343 */
128'h061300006617e789aa06061300006617, /* 1344 */
128'h4581346000efb265051300006517dfe6, /* 1345 */
128'hb28a0a1300006a174401ed9ff0ef8526, /* 1346 */
128'h01f4779320000913b289899300006997, /* 1347 */
128'h008487b3318000ef8552e7810004059b, /* 1348 */
128'h00ef819100f5f6130405854e0007c583, /* 1349 */
128'h00ef0d25051300006517fd241de33020, /* 1350 */
128'h45016a0269a2694264e2740270a22f20, /* 1351 */
128'h0003b6830083b7830103b70380826145, /* 1352 */
128'h079300d7fe6393811782278540f707b3, /* 1353 */
128'h45050103b78300a7002300f3b8230017, /* 1354 */
128'hb7830083b70380824501808200078023, /* 1355 */
128'h06930003b7038f999201020596130103, /* 1356 */
128'h47819d9dfff7059b00c6f5638e9dfff7, /* 1357 */
128'h0007002300b6e6630103b7030007869b, /* 1358 */
128'h00f506b300d3b823001706938082852e, /* 1359 */
128'h56634301bfd900d7002307850006c683, /* 1360 */
128'hc21906100693430540a0053be6810005, /* 1361 */
128'h089b385986ba4e250ff6f81304100693, /* 1362 */
128'h061b04ae6a630ff5761302b8f53b0005, /* 1363 */
128'h02b8d53bfec68fa306850ff676130306, /* 1364 */
128'h06bb0300059340e0063b8536fcb8ffe3, /* 1365 */
128'h002302d007930003076302f6e96300a6, /* 1366 */
128'h46810015559b9d1900050023050500f5, /* 1367 */
128'h063b808200b7ea630006879bfff5081b, /* 1368 */
128'h40f807bbb7d1feb50fa30505bf4500c8, /* 1369 */
128'h48830007c30300d7063397ba93811782, /* 1370 */
128'h7119b7e1011780230066002306850006, /* 1371 */
128'he4d6e8d2eccef4a6f8a2597d011cf0ca, /* 1372 */
128'hf82af02ef42afc3e843684b2e0dafc86, /* 1373 */
128'h0209591303000a9306c00a1302500993, /* 1374 */
128'h0017079bc52d8f1d0004c50377a27742, /* 1375 */
128'h04850135086304d7ff63938117827682, /* 1376 */
128'h0f630014c503bfe1e71ff0ef02010393, /* 1377 */
128'hcb9d0004c78303551063478104890545, /* 1378 */
128'h478100f6f36346a50ff7f793fd07879b, /* 1379 */
128'heb6306d50f630640069304890014c503, /* 1380 */
128'h09630630079304d50f630580069302a6, /* 1381 */
128'h6a4669e6790674a6744670e6f55d08f5, /* 1382 */
128'h0024c503808261090007051b6b066aa6, /* 1383 */
128'h00a76c6306e50e6307300713b74d048d, /* 1384 */
128'h4685003800840b13f6e51ee307000713, /* 1385 */
128'h0780071302e5006307500713a00d4601, /* 1386 */
128'h4685003800840b13fa850613f6e510e3, /* 1387 */
128'h00840b13f8b50693a81145c100163613, /* 1388 */
128'he31ff0ef400845a946010016b6930038, /* 1389 */
128'ha809dd1ff0ef0028020103930005059b, /* 1390 */
128'hd89ff0ef00840b130201039300044503, /* 1391 */
128'h852201247433600000840b13b5fd845a, /* 1392 */
128'hb7f18522020103930005059b501010ef, /* 1393 */
128'he4c6e0c2fc3ef83aec061034f436715d, /* 1394 */
128'hf032715d8082616160e2e8dff0efe436, /* 1395 */
128'hfc3ef83aec06100005931014862ef436, /* 1396 */
128'h8082616160e2e69ff0efe436e4c6e0c2, /* 1397 */
128'h100005931234862afe36fa32f62e710d, /* 1398 */
128'he436eec6eac2e6bee2baea22ee060808, /* 1399 */
128'h60f28522157020ef0808842ae3fff0ef, /* 1400 */
128'h03630087b303679c691c808261356452, /* 1401 */
128'h469704b7ec63479d8082450183020003, /* 1402 */
128'h1101431c973600259713502686930000, /* 1403 */
128'h08c52483795c878297b6e426e822ec06, /* 1404 */
128'h029454330e7010ef908114827540f55c, /* 1405 */
128'h7d5c8082610545016442e90064a260e2, /* 1406 */
128'h659c95aa058e05e135f1bfe1617cbff1, /* 1407 */
128'he406e02211418082557d8082557db7f1, /* 1408 */
128'hb303679c681c00055e63ff5ff0ef842a, /* 1409 */
128'h8302014160a264028522000307630207, /* 1410 */
128'h47ad8082557d80820141640260a24501, /* 1411 */
128'h817549a7879300004797150200a7eb63, /* 1412 */
128'h808271a505130000551780826108953e, /* 1413 */
128'h102347a1715d83020007b303679c691c, /* 1414 */
128'he83ee42e078517824785d23e47d502f1, /* 1415 */
128'hf0efcc3ed402e486100c200007930030, /* 1416 */
128'he063400407374d148082616160a6fd3f, /* 1417 */
128'h980101f1041322813823dc01011308e6, /* 1418 */
128'hf0ef1a05348322113c232291342385a2, /* 1419 */
128'h00f70d630a0447830a04c703e909fadf, /* 1420 */
128'h228134832301340323813083fb600513, /* 1421 */
128'h11e30dd447830dd4c703808224010113, /* 1422 */
128'hc703fcf71be30c0447830c04c703fef7, /* 1423 */
128'h0d4405934611fcf715e30e0447830e04, /* 1424 */
128'h4501bf654501fd4559b010ef0d448513, /* 1425 */
128'h20eff4063e800513842af02271798082, /* 1426 */
128'hc202c40200011023858a4601852271c0, /* 1427 */
128'h6fe020ef7d000513e509842af21ff0ef, /* 1428 */
128'h10234785717980826145740270a28522, /* 1429 */
128'hc195842ac402c23ef406f022478500f1, /* 1430 */
128'h8ff9f80686934bdc008006b74538691c, /* 1431 */
128'h8fd9400007378fd98f75600006b78ff5, /* 1432 */
128'h47b2e119ec9ff0ef8522858a4601c43e, /* 1433 */
128'h102347b5711d80826145740270a2c43c, /* 1434 */
128'hf852fc4ee0ca07c55783c23e47d500f1, /* 1435 */
128'he4a6e8a26a056989fdf949370107979b, /* 1436 */
128'h09134495c43e842e8b2af456ec86f05a, /* 1437 */
128'h855a858a4601e00a0a13e00989930809, /* 1438 */
128'hf7b3c7891005f79345b2ed15e71ff0ef, /* 1439 */
128'h00005517c7950125f7b3054795630135, /* 1440 */
128'h644660e6fba00513d4dff0ef57450513, /* 1441 */
128'h808261257b027aa27a4279e2690664a6, /* 1442 */
128'h051300805863fff40a9bfe04c5e334fd, /* 1443 */
128'h47e345018456b74d8456608020ef3e80, /* 1444 */
128'h0513d07ff0ef5465051300005517fc80, /* 1445 */
128'h102347c17139e7a919c52783bf6df920, /* 1446 */
128'hf426fc06f822858a460147d5c42e00f1, /* 1447 */
128'h8b891b842783c11ddddff0efc23e842a, /* 1448 */
128'hc901dc7ff0ef8522858a46014495cb91, /* 1449 */
128'h45018082612174a2744270e2f8ed34fd, /* 1450 */
128'he8a2ec86e0cae4a6711d80824501bfd5, /* 1451 */
128'h02c9270347c906d7f66384b6892a4785, /* 1452 */
128'h4755d432cf3108c92783260102f11023, /* 1453 */
128'hca26d23a854a100c47850030cc3ee42e, /* 1454 */
128'h0497f0634785e529842ad6fff0efc83e, /* 1455 */
128'hd402854a100c47f5460102f1102347b1, /* 1456 */
128'h4a05051300005517c11dd4fff0efd23e, /* 1457 */
128'h6125690664a6644660e68522c41ff0ef, /* 1458 */
128'h0004841bb74d02f6063bbf6147c58082, /* 1459 */
128'hf04af426f822fc067139b7c54401b7d5, /* 1460 */
128'h84b28a2e4148842ace05e456e852ec4e, /* 1461 */
128'h852200b44583c11d892a4a4010ef8ab6, /* 1462 */
128'h7a63014485b3681000054d63905fa0ef, /* 1463 */
128'h4481bd7ff0ef456505130000551700b6, /* 1464 */
128'h89a6f96decdff0ef854a08c92583a089, /* 1465 */
128'h86a2844e0089f3630207e40301093783, /* 1466 */
128'h6783fc851ae3f01ff0ef854a85d68652, /* 1467 */
128'h99e39aa2028784339a22408989b308c9, /* 1468 */
128'h6a4269e274a279028526744270e2fc09, /* 1469 */
128'h71390106161b0086969b808261216aa2, /* 1470 */
128'h47f58e5500f11023030006b78e554799, /* 1471 */
128'h4601440dc432c23e84aafc06f426f822, /* 1472 */
128'h85263e800593e919c4dff0ef8526858a, /* 1473 */
128'h347d8082612174a2744270e2d8bff0ef, /* 1474 */
128'h3823bffc07b7db0101134d18bfcdfc79, /* 1475 */
128'h22913c2324813023241134239fb92321, /* 1476 */
128'h04131ce7f36349013ffc073723313423, /* 1477 */
128'h1a63892ac03ff0ef84aa85a2980101f1, /* 1478 */
128'h792020ef20000513e7991a04b7831e05, /* 1479 */
128'h200006131e0505631a04b5031aa4b023, /* 1480 */
128'h1cf76d6347210c04478313d010ef85a2, /* 1481 */
128'h07b753b897ba078a0407071300004717, /* 1482 */
128'h0d44278300e7fd63cc981ff787934004, /* 1483 */
128'h00d773630147d69307a6800707136705, /* 1484 */
128'h8b8506f48f2309b449830a044783f8dc, /* 1485 */
128'h0b344783c7890e244783e7810019f993, /* 1486 */
128'hc7898b890a04478300098a6308f480a3, /* 1487 */
128'h091407130e24478306f48fa309c44783, /* 1488 */
128'h09d405130a844783fcdc07c60c848613, /* 1489 */
128'h979b00074583fff74783e0fc07c64681, /* 1490 */
128'hc39197aeffe745839fad0105959b0087, /* 1491 */
128'h478302f585b30e04458300098c634685, /* 1492 */
128'h14e30621070de21c07ce02b787b30dd4, /* 1493 */
128'h468508d4470308e4478304098f63fce5, /* 1494 */
128'h97ba08c447039fb90087171b0107979b, /* 1495 */
128'h02e787b30dd4478302f707330e044703, /* 1496 */
128'h0187979b08a4470308b44783f8fc07ce, /* 1497 */
128'h9fb90087171b089447039fb90107171b, /* 1498 */
128'hf4fc07a6c319f4fc54d89fb908844703, /* 1499 */
128'he3918bfd09c44783c7898b850a044783, /* 1500 */
128'he0bff0ef852645850af006134685c6b5, /* 1501 */
128'h00a7979b0e0447830af407a34785e141, /* 1502 */
128'h0d44278300098663c79954dc08f4aa23, /* 1503 */
128'h02e787bb0dd447030e044783f8dc07a6, /* 1504 */
128'h08f480230a74478308f4ac2300a7979b, /* 1505 */
128'h390323813483854a2401340324813083, /* 1506 */
128'h0af44783808225010113228139832301, /* 1507 */
128'h8b7d0057d79b00a7d71b50fcf3dd8b85, /* 1508 */
128'hb75d08f4aa2302f707bb278527058bfd, /* 1509 */
128'h1a04b0235f0020efdd4d1a04b503892a, /* 1510 */
128'h3c23dc010113b7655929b7755951bf45, /* 1511 */
128'h47892321302322913423228138232211, /* 1512 */
128'h842eed8554a9468104b7ec6306f58463, /* 1513 */
128'he11d84aad3fff0ef892a45850b900613, /* 1514 */
128'h980101f10413ed91258199f5ffe4059b, /* 1515 */
128'he3990b944783e9159a7ff0ef854a85a2, /* 1516 */
128'h390385262301340323813083df400493, /* 1517 */
128'hffc5879b808224010113228134832201, /* 1518 */
128'hbfd984aab7554685fef760e354a94705, /* 1519 */
128'h08154783f022f406e44ee84aec267179, /* 1520 */
128'h06138edd892e9be10079f6930ff5f993, /* 1521 */
128'h842a57b5c519cc1ff0ef84aa45850b30, /* 1522 */
128'h86dff0ef852685ca00091c6300f51e63, /* 1523 */
128'h70a28522013505a317a010ef8526842a, /* 1524 */
128'hd60101138082614569a2694264e27402, /* 1525 */
128'h29213023289134232881382328113c23, /* 1526 */
128'h27613023275134232741382327313c23, /* 1527 */
128'h25a13023259134232581382325713c23, /* 1528 */
128'hbffc07b74d180ac7ed63478923b13c23, /* 1529 */
128'h84aabfe787933ffc07b79f3dbff7879b, /* 1530 */
128'h00e7eb6305450513000055178a2e8b32, /* 1531 */
128'h051300005517e7b90016f79307e4c683, /* 1532 */
128'h298130838522f8400413f8eff0ef0765, /* 1533 */
128'h27813983280139032881348329013403, /* 1534 */
128'h25813b8326013b0326813a8327013a03, /* 1535 */
128'h23813d8324013d0324813c8325013c03, /* 1536 */
128'h0513000055170984a70380822a010113, /* 1537 */
128'hfe09f99302f109930045aa83db4504e5, /* 1538 */
128'hf7bb0005ac83e79102eaf7bb060a8063, /* 1539 */
128'hf14ff0ef04c5051300005517cb8902ec, /* 1540 */
128'h9c9be3994b8502eadabb54dcb7615429, /* 1541 */
128'h4e0547818956866200ca05138c0a009c, /* 1542 */
128'h8d6302e878bb0017859b000528034311, /* 1543 */
128'hb7c9ed6ff0ef04650513000055170008, /* 1544 */
128'h0116202302e858bbb7f14b814a814c81, /* 1545 */
128'hcb898b850107c78397d2078e02080063, /* 1546 */
128'h0128893b0ffbfb9300fbebb300be17bb, /* 1547 */
128'h8a89000b8963fa6596e387ae06110521, /* 1548 */
128'h852685ceee068de30285051300005517, /* 1549 */
128'hc78309f9c603ee051ae3842af8aff0ef, /* 1550 */
128'h09d9c7839e3d0087979b0106161b09e9, /* 1551 */
128'h020505130000551785ca01267a63963e, /* 1552 */
128'hf7130a79c683008a4783b5c9e50ff0ef, /* 1553 */
128'he913c3990fe6f9138b89c71989360017, /* 1554 */
128'h97d2078e0017861b4591450547810016, /* 1555 */
128'h571b00c517bbc39d8b850017579b4b98, /* 1556 */
128'h4187d79b8b050189191b0187979b0027, /* 1557 */
128'h87b20ff979130127e933c70d4189591b, /* 1558 */
128'hef898b850a69c78302d90263fcb614e3, /* 1559 */
128'hc793b5a939c020effd85051300005517, /* 1560 */
128'hcb898b8509b9c783bfd100f97933fff7, /* 1561 */
128'hb535547ddb8ff0ef0085051300005517, /* 1562 */
128'h06134685e3958b850af9c783e20b05e3, /* 1563 */
128'h87a34785e579a21ff0ef852645850af0, /* 1564 */
128'h4d0108f4aa2300a7979b0e09c7830af9, /* 1565 */
128'hf693f88d061b00dcd6bb003d169b4d91, /* 1566 */
128'h8a2a9edff0ef852645850ff676130ff6, /* 1567 */
128'hd6bb003a169b4c8dfdbd1fe32d05e945, /* 1568 */
128'h45850ff676130ff6f693f8ca061b00da, /* 1569 */
128'h0a13ff9a10e32a05e92d9c5ff0ef8526, /* 1570 */
128'h000c26834c818ad209b00d934d6108f0, /* 1571 */
128'hf0ef85260ff6f6930196d6bb45858656, /* 1572 */
128'hffac90e30ffafa932ca12a85e139999f, /* 1573 */
128'h061386defdba18e30c110ffa7a132a0d, /* 1574 */
128'h0ee34785ed19971ff0ef8526458509c0, /* 1575 */
128'h09b00613468501279b630a79c783d4fb, /* 1576 */
128'h061386cab381842a953ff0ef85264585, /* 1577 */
128'hb335dd79842a941ff0ef852645850a70, /* 1578 */
128'hffdfe0ef842ae406e0221141b325842a, /* 1579 */
128'h000307630187b303679c681c00055e63, /* 1580 */
128'h640260a245058302014160a264028522, /* 1581 */
128'h4791f04af822fc06f426713980820141, /* 1582 */
128'h079304f592635529478500f5866384aa, /* 1583 */
128'h979b4955842e07c4d78300f110230370, /* 1584 */
128'hd44ff0efc43ec24a8526858a46010107, /* 1585 */
128'h00f41f634791c24a00f110234799ed19, /* 1586 */
128'h70e2d26ff0ef8526858a4601c43e4789, /* 1587 */
128'hfef414e3478580826121790274a27442, /* 1588 */
128'hf3630007869b4f5c6918e215b7cdc402, /* 1589 */
128'hf3630007069b0007859b4f1887ae00d5, /* 1590 */
128'hf06f02c50823dd0c0007859b87ba00d5, /* 1591 */
128'h4b9c711910000737691c80828082c18f, /* 1592 */
128'he4d6e8d2eccef0caf4a6fc86f8a2070d, /* 1593 */
128'hf0ef842ac17c8fd9f466f862fc5ee0da, /* 1594 */
128'h02042423eb8d6b9c679c681cc509f07f, /* 1595 */
128'hf8500493b98ff0efe085051300005517, /* 1596 */
128'h6aa66a4669e674a679068526744670e6, /* 1597 */
128'h4481541c808261097ca27c427be26b06, /* 1598 */
128'h082347851af42c23478df93ff0eff3e5, /* 1599 */
128'h7d000513b8eff0ef852202042c2302f4, /* 1600 */
128'h84aa97826b9c679c8522681c43b010ef, /* 1601 */
128'h22231a04282318042e2308842783f945, /* 1602 */
128'h45814601b5eff0ef8522d85c478508f4, /* 1603 */
128'hf14984aacdaff0ef8522f13ff0ef8522, /* 1604 */
128'h00f1102347a1000505a346d000ef8522, /* 1605 */
128'he3991aa007138ff94bdc00ff8737681c, /* 1606 */
128'hc23ec43a8522858a460147d50aa00713, /* 1607 */
128'h15630aa0079300c14703e911be0ff0ef, /* 1608 */
128'h037009933e900913cc1c800207b700f7, /* 1609 */
128'h80020c3700ff8bb74b0502900a934a55, /* 1610 */
128'hc252013110238522858a460140000cb7, /* 1611 */
128'h015110234c18681ce13db9eff0efc402, /* 1612 */
128'he7b301871563c43e0177f7b3c25a4bdc, /* 1613 */
128'hed1db76ff0ef8522858a4601c43e0197, /* 1614 */
128'h3e80051306090863397d0007ca6347b2, /* 1615 */
128'h00e68563800207374c14bf4534b010ef, /* 1616 */
128'hd45c8b8541e7d79bc43ccc1880010737, /* 1617 */
128'hf9200793b55d18f40ca3478506041e23, /* 1618 */
128'hf0ef85224581becff0ef852202f51f63, /* 1619 */
128'h18f40c2347850007d663443ced09c1cf, /* 1620 */
128'h00005517d965c04ff0ef85224585bfd1, /* 1621 */
128'h84aab595fa1004939fcff0efc8450513, /* 1622 */
128'he74eeb4aef26f706f3227161551cb585, /* 1623 */
128'he6eeeaeaeee6f2e2f6defadafed6e352, /* 1624 */
128'h199bc783219010ef45018baae3b54401, /* 1625 */
128'h10234789e7b5180b8ca3198bc783c7b1, /* 1626 */
128'hf0efc482c2be855e008c479d460104f1, /* 1627 */
128'hcf818b851b8ba78312050ae3842aaa2f, /* 1628 */
128'h0de3842aa88ff0ef855e008c46014495, /* 1629 */
128'hf0ef855ea031020ba423f4fd34fd1005, /* 1630 */
128'h695a64fa741a70ba8522d55d842ad99f, /* 1631 */
128'h6d566cf67c167bb67b567af66a1a69ba, /* 1632 */
128'hc163180b8c23048ba7838082615d6db6, /* 1633 */
128'h1493187010ef4501afeff0ef855e0407, /* 1634 */
128'hb1eff0ef855e45853e80091390810205, /* 1635 */
128'h10ef85260007cc63048ba783f155842a, /* 1636 */
128'hbfe91f1010ef0640051308a96fe31630, /* 1637 */
128'h41e7d79b048ba78300fbac23400007b7, /* 1638 */
128'h0737bf0506fb9e23478502fba6238b85, /* 1639 */
128'h4007071b40010737a0292007071b4001, /* 1640 */
128'h0a1300003a178a1d0036571b00ebac23, /* 1641 */
128'h47031086260396529752060a8b3d646a, /* 1642 */
128'h00c7d61b02c7073b018ba88345050f87, /* 1643 */
128'ha42304cba823180bae231a0ba8238a05, /* 1644 */
128'h00e5183b8b3d0107d71b08eba22308eb, /* 1645 */
128'h02cba703090ba8231408dd63090ba623, /* 1646 */
128'hd79b8f7d003f07370107979b14070f63, /* 1647 */
128'h87b300d797b32689078546a18fd90106, /* 1648 */
128'hb8230c0bb4230c0bb0230a0bbc230307, /* 1649 */
128'h07930afbb8230e0bb0230c0bbc230c0b, /* 1650 */
128'h0793090ba70308fba6230107d4632000, /* 1651 */
128'h04cba783c21508fba82300e7f4632000, /* 1652 */
128'h008c46010107979b471100e78e63577d, /* 1653 */
128'h479d8f6ff0efc282c4be04e11023855e, /* 1654 */
128'h0107979b4601495507cbd78304f11023, /* 1655 */
128'h1ce3842a8d8ff0efc4bec2ca855e008c, /* 1656 */
128'h855e08fb80a357fd08fbaa234785e405, /* 1657 */
128'h113000ef855ee40510e3842ac94ff0ef, /* 1658 */
128'he20515e3842aff3fe0ef855e00b54583, /* 1659 */
128'ha0232789100007b754075963018ba703, /* 1660 */
128'h460107cbd78306f110230370079304fb, /* 1661 */
128'h874ff0efd4bed2ca855e0107979b108c, /* 1662 */
128'h1a93033007930bf104934905d2caed05, /* 1663 */
128'h4b210a854991d48206f1102398810209, /* 1664 */
128'h844ff0efd05aec56e826855e108c0810, /* 1665 */
128'h40020737bb75842afe0996e339fdc529, /* 1666 */
128'hd59bbd9140040737bda940030737bd89, /* 1667 */
128'h6705b54508bba82300b515bb89bd0165, /* 1668 */
128'h17828fd901e6d71b8ff90027979b1771, /* 1669 */
128'h00ff05374098bd798a9d938100f6d69b, /* 1670 */
128'h8e698fd50087161b0187179b0187569b, /* 1671 */
128'h8fd58ef1f00706138fd167410087569b, /* 1672 */
128'h0187169b0187559b40d804fbaa232781, /* 1673 */
128'h8f718ecd0087571b8de90087159b8ecd, /* 1674 */
128'h09270d638b3d0187d71b04ebac238f55, /* 1675 */
128'h00ebac238001073708d70e634689c701, /* 1676 */
128'h20000737040ba7830007596302d79713, /* 1677 */
128'h1363800107b7018ba70304fba0238fd9, /* 1678 */
128'h040ba903639c06e787930000579708f7, /* 1679 */
128'h849300003497044ba783f0be0ff10c13, /* 1680 */
128'h02079a93478500f97933fe0c7c9345e4, /* 1681 */
128'h77b300e797bb478540980a8583f97913, /* 1682 */
128'h440787930000379704a1ebc5278100f9, /* 1683 */
128'he15fe0ef8cc5051300005517fef493e3, /* 1684 */
128'hb7bda007071b80011737b949df400413, /* 1685 */
128'h0737b785800207370007456303079713, /* 1686 */
128'h190201000ab70ff104934905bfa98003, /* 1687 */
128'h47990209886339fd09053ac549959881, /* 1688 */
128'h010c040007931030c33e47d508f11023, /* 1689 */
128'h1de3eb7fe0efdc3ef84af426c556855e, /* 1690 */
128'h0713674144dcfbe18b8583a54cdce605, /* 1691 */
128'h97138fd58ff90087d79b0087969bf007, /* 1692 */
128'ha0230087e793040ba783f20750e302e7, /* 1693 */
128'h840b0b1b06010993017d8b37bf0104fb, /* 1694 */
128'h278101a7f7b300f977b30009ad0340dc, /* 1695 */
128'h07b700fd0d6345a1400007b712078e63, /* 1696 */
128'h40bd05b3100005b700fd086345912000, /* 1697 */
128'h0e0519638daa8bfff0ef855e0015b593, /* 1698 */
128'h47912000073700ed0d6347a140000737, /* 1699 */
128'h001d379340fd0d33100007b700ed0863, /* 1700 */
128'h86634705409cd41fe0ef855e02fbaa23, /* 1701 */
128'h0af1102347994d850ae79d63470d00e7, /* 1702 */
128'h00fde7b317c12d81810007b7d33e47d5, /* 1703 */
128'he556e166855e110c040007930110d53e, /* 1704 */
128'h90638bbd010cc783e541dcffe0efc93e, /* 1705 */
128'h17ed088ba583efd91afba823409c09b7, /* 1706 */
128'h855e460118fbae2308bba2230017b793, /* 1707 */
128'h07cbd7830af1102303700793895ff0ef, /* 1708 */
128'he03ad33a855e110c0107979b46014755, /* 1709 */
128'hfe0c7d1347b56702ed05d7ffe0efd53e, /* 1710 */
128'h040007134791d5028dead33a0af11023, /* 1711 */
128'he03ac93ae556e16ae43e855e110c0110, /* 1712 */
128'h4785f3f537fd670267a2c521d51fe0ef, /* 1713 */
128'h180bae23096ba2231afba823017d85b7, /* 1714 */
128'h10bc099181dff0ef855e840585934601, /* 1715 */
128'h9713f6f762e34581472db575def98be3, /* 1716 */
128'h059366c1bf9111872583975283790207, /* 1717 */
128'h0d11000d2783f006869300ff0537040d, /* 1718 */
128'h8e690087961b8f510187971b0187d61b, /* 1719 */
128'h9ee3fefd2e238fd98ff58f510087d79b, /* 1720 */
128'hf8638bbd00c7579b46a5008da703fda5, /* 1721 */
128'h369704d61c63800306b7018ba60300f6, /* 1722 */
128'h171b1487a78397b6078a132686930000, /* 1723 */
128'hd61b17fd67c100cda68308fbae230087, /* 1724 */
128'h77130126d71bc78d27818fd18ff90186, /* 1725 */
128'h0106d69b02e6073b3e800613c30503f7, /* 1726 */
128'ha2230afba02302d606bb02f757bb8a8d, /* 1727 */
128'hc79919cba7831afbaa231b0ba7830adb, /* 1728 */
128'h00ef855e08fba82308fba62320000793, /* 1729 */
128'hb7b708cba70300050623000515234a00, /* 1730 */
128'h8ff9ccc68693aaa78793ccccd6b7aaaa, /* 1731 */
128'h9fb500f037b3068600d036b327818ef9, /* 1732 */
128'h068a00d036b38ef90f068693f0f0f6b7, /* 1733 */
128'h00d036b38ef9f0068693ff0106b79fb5, /* 1734 */
128'h00e037338f750207161376c19fb5068e, /* 1735 */
128'hd7b3ed1092010a8bb783d11c9fb90712, /* 1736 */
128'h84aa06fbc603074bd68307abd70302c7, /* 1737 */
128'hfef53623024505135a85859300004597, /* 1738 */
128'h06cbc603077bc883070ba683a8dfe0ef, /* 1739 */
128'h0ff7f7930ff6f8130106d71b0086d79b, /* 1740 */
128'h58858593000045970186d69b0ff77713, /* 1741 */
128'h00004597074ba603a59fe0ef04d48513, /* 1742 */
128'h0146561b0106569b0624851358458593, /* 1743 */
128'h478500d010ef8526a39fe0ef8a3d8abd, /* 1744 */
128'h04fba0232785100007b7b0cd02fba423, /* 1745 */
128'h400407b700f778631a0bb603400407b7, /* 1746 */
128'h051300004517e611b5f1e225ecf769e3, /* 1747 */
128'h04fba0230016879b700006b7b1294f65, /* 1748 */
128'h0027f5931abba42303f7f5930c464783, /* 1749 */
128'h04dba0230216869bc58900c7f593cd91, /* 1750 */
128'hd7dd8b8504dba0230106e693040ba683, /* 1751 */
128'h400407b704fba02300c7e793040ba783, /* 1752 */
128'h088ba583044ba783040ba983e6f769e3, /* 1753 */
128'h3497daaff0ef2981855e00f9f9b34601, /* 1754 */
128'hfe0b0b1300003b174a85fca484930000, /* 1755 */
128'h00fa97bb409c012c8c9300003c974c2d, /* 1756 */
128'h4517ff6498e304a1eb99278100f9f7b3, /* 1757 */
128'h00003917bd2197bfe0ef432505130000, /* 1758 */
128'h4703409c10000db720000d37fac90913, /* 1759 */
128'h270340dc04f719630017b79317ed0049, /* 1760 */
128'h00894683c3a127818ff900f9f7b30009, /* 1761 */
128'hdbbfe0ef855e0fb6f69345850b700613, /* 1762 */
128'hdabfe0ef855e45850b7006134681c90d, /* 1763 */
128'h08fba223180bae231a0ba823088ba783, /* 1764 */
128'hfb9910e30931941fe0ef855e035baa23, /* 1765 */
128'h00d789634721400006b700092783bfa5, /* 1766 */
128'haa230017b71341b787b301a786634711, /* 1767 */
128'hfeffe0ef855e408c913fe0ef855e02eb, /* 1768 */
128'ha823409ce79d0046f79300892683f14d, /* 1769 */
128'ha2230017b79317ed088ba583ef8d1afb, /* 1770 */
128'h855ec9aff0ef855e460118fbae2308bb, /* 1771 */
128'h0b7006130ff6f693bb35f53d9d9fe0ef, /* 1772 */
128'h65e34581bfa1d171d13fe0ef855e4585, /* 1773 */
128'hbf6d118725839752837902079713fcfc, /* 1774 */
128'h06cb851300ec4641ef2ff06ffa100413, /* 1775 */
128'h460107cbd78304f11023478d6ce000ef, /* 1776 */
128'he0efc2be47d5855ec4be0107979b008c, /* 1777 */
128'h0007d663018ba783ec051163842a943f, /* 1778 */
128'h479d04f1102347a506fb9e2304e15783, /* 1779 */
128'h855e0107979b008c460107cbd783c2be, /* 1780 */
128'h47c64636e8051763842a90ffe0efc4be, /* 1781 */
128'h06fba02304cbae23018ba50345e646d6, /* 1782 */
128'hf0e51c634000073706bba42306dba223, /* 1783 */
128'h6863450d0007081b377d8b3d01a6571b, /* 1784 */
128'h972a8379d3c50513000035171702ef05, /* 1785 */
128'h8082557d80824501c56c8702972a4318, /* 1786 */
128'h879300005797808218b50d238082557d, /* 1787 */
128'h842ae406e02247851141ef9d439cbfa7, /* 1788 */
128'he0ef852212a000efbef7222300005717, /* 1789 */
128'h02c00513fc5ff0ef852200055563ac0f, /* 1790 */
128'h01414501640260a20dc000ef13e000ef, /* 1791 */
128'h631cbb27071300005717808245018082, /* 1792 */
128'h05130000451785aa114102e790636394, /* 1793 */
128'h0141853e478160a2f3cfe0efe4063665, /* 1794 */
128'h853ebfd187b600a604630fc7a6038082, /* 1795 */
128'hc105fbdff0efe42eec06110141488082, /* 1796 */
128'h07930815470302b7006365a210354703, /* 1797 */
128'h5535e97fe06f610560e200f70c630ff0, /* 1798 */
128'hbfcdf8400513bfe545018082610560e2, /* 1799 */
128'hcd09f7dff0ef84aee822ec06e4261101, /* 1800 */
128'h60e2e0800f840413e501ce0ff0ef842a, /* 1801 */
128'h00005797bfd555358082610564a26442, /* 1802 */
128'h05138082c3980015071b438895478793, /* 1803 */
128'h8082438893c787930000579780820f85, /* 1804 */
128'he4266380e822ae678793000057971101, /* 1805 */
128'h610564a2644260e20094176384beec06, /* 1806 */
128'h6000a8cff0ef8522c78119a447838082, /* 1807 */
128'h5797e79ce39cab67879300005797b7d5, /* 1808 */
128'h879300005797e50880828e07a9230000, /* 1809 */
128'h711d8082e308e518e11ce7886798a9e7, /* 1810 */
128'hfc4e6080e8a2a864849300005497e4a6, /* 1811 */
128'hec86e06ae466e862ec5ef05af456f852, /* 1812 */
128'h00004a9724ca0a1300004a1789aae0ca, /* 1813 */
128'h00004b9724cb0b1300004b1724ca8a93, /* 1814 */
128'h830c8c9300004c9700050c1b24cb8b93, /* 1815 */
128'h79e2690664a660e66446029415634d29, /* 1816 */
128'h45176d026ca26c426be27b027aa27a42, /* 1817 */
128'h4901541cdb8fe06f612539a505130000, /* 1818 */
128'h2603681c89560007c36389524c1cc791, /* 1819 */
128'h85ca00090663d9afe0ef638c855a0fc4, /* 1820 */
128'h856685e200978e63601cd8efe0ef855e, /* 1821 */
128'h7b8505130000351701a98863d80fe0ef, /* 1822 */
128'he426ec06e8221101b7716000334010ef, /* 1823 */
128'hcbbd4d5ccfad44014d1cc1414401e04a, /* 1824 */
128'h84aa892ec7ad639cc7bd651ccbad511c, /* 1825 */
128'h57fdcd21842a20a010ef45051c000593, /* 1826 */
128'he90410f502a347850ef52c234799c57c, /* 1827 */
128'hfffff797e65ff0ef0405282303253023, /* 1828 */
128'h2c8787930000179716f43c238fa78793, /* 1829 */
128'h18f434232b8787930000179718f43023, /* 1830 */
128'h10f400230247c78385220ea42e23681c, /* 1831 */
128'h6105690264a2644260e28522e99ff0ef, /* 1832 */
128'h611c6d268693000046971c60106f8082, /* 1833 */
128'he11897360017671302d786b365186294, /* 1834 */
128'h07bb00f7553b93ed836d8f3d0127d713, /* 1835 */
128'h00005517808225018d5d00f717bb40f0, /* 1836 */
128'hf0efe022e4061141fc3ff06f8fc50513, /* 1837 */
128'h60a28d410105151bfe9ff0ef842afeff, /* 1838 */
128'hf0efe022e40611418082014125016402, /* 1839 */
128'h15029001fd1ff0ef14020005041bfdbf, /* 1840 */
128'hc703058587aa80820141640260a28d41, /* 1841 */
128'h8c6347818082fb75fee78fa30785fff5, /* 1842 */
128'h078500f506b30007470300f5873300c7, /* 1843 */
128'h86930007c70387aa8082f76d00e68023, /* 1844 */
128'hfee78fa30785fff5c7030585eb090017, /* 1845 */
128'h87b68082e21987aab7d587b68082fb75, /* 1846 */
128'hc7030585963efb7d001786930007c703, /* 1847 */
128'h8023fec799e3d375fee78fa30785fff5, /* 1848 */
128'h07bbfff5c78300054703058580820007, /* 1849 */
128'hf37d0505e3994187d79b0187979b40f7, /* 1850 */
128'h07b3a015478100e6146347018082853e, /* 1851 */
128'h87bb0007c78300e587b30007c68300e5, /* 1852 */
128'hfee10705e3994187d79b0187979b40f6, /* 1853 */
128'h00b79363000547830ff5f5938082853e, /* 1854 */
128'h0ff5f59380824501bfcd0505c3998082, /* 1855 */
128'hbfcd0505dffd808200b7936300054783, /* 1856 */
128'h0785808240a78533e7010007c70387aa, /* 1857 */
128'hfe5ff0efec06842ae42ee8221101bfcd, /* 1858 */
128'h00b78663000547830ff5f593952265a2, /* 1859 */
128'h80826105644260e24501fe857be3157d, /* 1860 */
128'h8533e7010007c70300b7856387aa95aa, /* 1861 */
128'h468300f507334781b7fd0785808240a7, /* 1862 */
128'h46030705fed60ee38082853eea990007, /* 1863 */
128'h07334781bfd5872eb7d50785fa7d0007, /* 1864 */
128'h00d60863a021872eca890007468300f5, /* 1865 */
128'hb7c507858082853efa7d000746030705, /* 1866 */
128'h0785fee68fe380824501eb1900054703, /* 1867 */
128'h1101bfd587aeb7e50505fafd0007c683, /* 1868 */
128'h00004797e519842a84aeec06e426e822, /* 1869 */
128'hfa1ff0ef85a68522cc1163806fc78793, /* 1870 */
128'h6e07b02300004797ef8100044783942a, /* 1871 */
128'h85a68082610564a2644260e285224401, /* 1872 */
128'h0023c78100054783c519f9fff0ef8522, /* 1873 */
128'h1101bfd96aa7ba230000479705050005, /* 1874 */
128'hf0ef8526842ac891e822ec066104e426, /* 1875 */
128'h644260e2e008050500050023c501f73f, /* 1876 */
128'hcf9900054783c11d8082610564a28526, /* 1877 */
128'h8082e3110017c703ce810007c68387aa, /* 1878 */
128'h80824501b7e5078900d780a300e78023, /* 1879 */
128'h07220ff5f69347a1eb0587aa00757713, /* 1880 */
128'h8833469d00c508b387aaffed8f5537fd, /* 1881 */
128'h02e787335761003657930106ee6340f8, /* 1882 */
128'h07a1808200c79763963e963a97aa078e, /* 1883 */
128'h0463b7f5feb78fa30785bfe9fee7bc23, /* 1884 */
128'h471d4781eb9d872a8b9d00b567b304b5, /* 1885 */
128'h07a100f506b30006b80300f586b3a811, /* 1886 */
128'h00365793fed765e340f606b30106b023, /* 1887 */
128'h00f50733963a95be078e02e787335761, /* 1888 */
128'h0006c80300f586b3808200f613634781, /* 1889 */
128'hf0227179b7e501068023078500f706b3, /* 1890 */
128'hf0efe02ee84af406e432ec26852e842a, /* 1891 */
128'h00c564636582892ace1184aa6622dd3f, /* 1892 */
128'h0023f75ff0ef944a864a8522fff60913, /* 1893 */
128'h8082614564e269428526740270a20004, /* 1894 */
128'hf53ff0ef00a5e963842ae406e0221141, /* 1895 */
128'h461386ae883280820141640260a28522, /* 1896 */
128'h85b300f80733fef605e317fd4781fff6, /* 1897 */
128'h4701b7e500b7002397220005c58300e6, /* 1898 */
128'h00e586b300e507b3a821478100e61463, /* 1899 */
128'h853ed3f59f9507050006c6830007c783, /* 1900 */
128'h8de300054783808200c51363962a8082, /* 1901 */
128'hec26852e842af0227179bfc50505feb7, /* 1902 */
128'h0005049bd19ff0ef892ee44ef406e84a, /* 1903 */
128'h408987bb008509bbd0dff0ef8522c899, /* 1904 */
128'h694264e2740270a2852244010097db63, /* 1905 */
128'hf83ff0ef852285ca86268082614569a2, /* 1906 */
128'h00c514630ff5f593962abfe10405d17d, /* 1907 */
128'hfeb70be3001507930005470380824501, /* 1908 */
128'h260100c7ef630ff5f59347c1b7ed853e, /* 1909 */
128'h1ce30007c7038082853e4781e60187aa, /* 1910 */
128'h4721c39d00757793b7f5367d0785feb7, /* 1911 */
128'hfcb69de30007c68387aa00a7083b9f1d, /* 1912 */
128'h953a93011702fed819e30007869b0785, /* 1913 */
128'h8fd90107179300b7e733008597938e19, /* 1914 */
128'heb1187aa27018edd0036571302079693, /* 1915 */
128'h367d0785f8b71fe30007c703d24d8a1d, /* 1916 */
128'hc70300d80a63008785130007b803bfcd, /* 1917 */
128'h87aabfa5fef51be30785f8b712e30007, /* 1918 */
128'h0300079300054703e7c9419cb7f1377d, /* 1919 */
128'h0f878793000027970015470306f71e63, /* 1920 */
128'h0207071bc6898a850006c68300e786b3, /* 1921 */
128'h0025470304d71763078006930ff77713, /* 1922 */
128'hc19c47c1cf950447f7930007c78397ba, /* 1923 */
128'h0015478302f71f630300079300054703, /* 1924 */
128'h8b0500074703973e0b07071300002717, /* 1925 */
128'h9c63078007130ff7f7930207879bc709, /* 1926 */
128'hbfed47a98082c19c47a1a809050900e7, /* 1927 */
128'h006c842ee82211018082fae78fe34741, /* 1928 */
128'h2817468100c16583f61ff0efc632ec06, /* 1929 */
128'h06330007079b00054703062808130000, /* 1930 */
128'hec0500089863044678930006460300f8, /* 1931 */
128'h8b6300467893808261058536644260e2, /* 1932 */
128'h050502d586b3feb7f4e3fd07879b0008, /* 1933 */
128'h0ff7f793fe07079bc6098a09b7d196be, /* 1934 */
128'hf426f8227139b7e1e008b7cdfc97879b, /* 1935 */
128'hf0ef84b2842ae42e00063023f04afc06, /* 1936 */
128'h790274a2744270e25529e90165a2b03f, /* 1937 */
128'hf5dff0ef8522082c892a862e80826121, /* 1938 */
128'h07858f81cb010007c703fe8782e367e2, /* 1939 */
128'hb7e94501e088fcf718e347a9fd279be3, /* 1940 */
128'hf2dff06f00e6846302d0071300054683, /* 1941 */
128'h40a0053360a2f23ff0efe40605051141, /* 1942 */
128'hf0dff0ef842ee406e022114180820141, /* 1943 */
128'hea6302d704630007c70304b00693601c, /* 1944 */
128'h0141640260a202d70e630470069300e6, /* 1945 */
128'h16e306b0069302d7076304d006938082, /* 1946 */
128'hfce69fe3052a069007130017c683fed7, /* 1947 */
128'he01c078d00e69863042007130027c683, /* 1948 */
128'he8221101bfd50789bff1052a052ab7e9, /* 1949 */
128'h00c16583e0dff0efc632ec06006c842e, /* 1950 */
128'h079b00054703f0e80813000028174681, /* 1951 */
128'h9863044678930006460300f806330007, /* 1952 */
128'h7893808261058536644260e2ec050008, /* 1953 */
128'h86b3feb7f4e3fd07879b00088b630046, /* 1954 */
128'hfe07079bc6098a09b7d196be050502d5, /* 1955 */
128'h1141b7e1e008b7cdfc97879b0ff7f793, /* 1956 */
128'h04b00693601cf87ff0ef842ee406e022, /* 1957 */
128'h0470069300e6ea6302d704630007c703, /* 1958 */
128'h04d0069380820141640260a202d70e63, /* 1959 */
128'h0017c683fed716e306b0069302d70763, /* 1960 */
128'h07130027c683fce69fe3052a06900713, /* 1961 */
128'h052a052ab7e9e01c078d00e698630420, /* 1962 */
128'he589842ae406e0221141bfd50789bff1, /* 1963 */
128'h00002797fff5c70300a405b3951ff0ef, /* 1964 */
128'h8b1100074703973efff58513e3478793, /* 1965 */
128'h7ae3157d80820141557d640260a2e719, /* 1966 */
128'hf77d8b1100074703973e00054703fea4, /* 1967 */
128'hd7dff06f014105054581462960a26402, /* 1968 */
128'h11418d5d05220085579bfa5ff06f4581, /* 1969 */
128'h2c878793000047978082014191411542, /* 1970 */
128'ha93ff06f95be9201160291811582639c, /* 1971 */
128'h8082853ee31900054703462946a54781, /* 1972 */
128'h9fb902f607bb00b6e763fd07059b2701, /* 1973 */
128'h842ee406e0221141b7c50505fd07879b, /* 1974 */
128'h02b455bb45a900b7f86347a500a04563, /* 1975 */
128'h60a2640202a4753b4529fe7ff0ef357d, /* 1976 */
128'h07e2081007935020006f030505130141, /* 1977 */
128'h24f738230000471724f7382300004717, /* 1978 */
128'he4262424041300004417e82211018082, /* 1979 */
128'h600ca05ff0efec06600885aa84ae862e, /* 1980 */
128'h11018082610564a26442e00c95a660e2, /* 1981 */
128'h849300004497e4262187879300004797, /* 1982 */
128'h7d050513000035176380e82260902064, /* 1983 */
128'hc0ef85a26088b5bfd0ef85a29c11ec06, /* 1984 */
128'h7c85051300003517862286aa608ce2df, /* 1985 */
128'hb35fd0ef7d45051300003517b41fd0ef, /* 1986 */
128'h00055e6385bf90efef85051300000517, /* 1987 */
128'h05130000351740a005b364a260e26442, /* 1988 */
128'h610564a260e26442b0dfd06f61057c65, /* 1989 */
128'h874fa0ef8432e406e022114166a0006f, /* 1990 */
128'h80820141640260a28522547d00850363, /* 1991 */
128'h89aae64e01258413f222716980824501, /* 1992 */
128'h0505f76ff0ef892eea4aee26f6068522, /* 1993 */
128'hf0ef95260505f6aff0ef852600a404b3, /* 1994 */
128'h479704e7ee631ff00793fff5071be93f, /* 1995 */
128'h351784aaf48ff0ef852212a7a5230000, /* 1996 */
128'h0ff007939526f3aff0ef53a505130000, /* 1997 */
128'h00003517842af2aff0ef852204a7f263, /* 1998 */
128'h0000351700a405b3f1cff0ef51c50513, /* 1999 */
128'h695264f2741270b2a5dfd0ef73450513, /* 2000 */
128'h272300004717200007938082615569b2, /* 2001 */
128'h855ff0ef850a458110000613b7550cf7, /* 2002 */
128'h4703de0ff0ef850a4d85859300003597, /* 2003 */
128'h85930000359700f7096302f007930129, /* 2004 */
128'hdecff0ef850a85a2df4ff0ef850a7065, /* 2005 */
128'h00003517858a43900887879300004797, /* 2006 */
128'h451107e2081007939edfd0ef6ec50513, /* 2007 */
128'h06f738230000471706f7382300004717, /* 2008 */
128'hf0ef4501e4a7962300004797d87ff0ef, /* 2009 */
128'h000045974611e4a7902300004797d79f, /* 2010 */
128'h000047174785eafff0ef854ee3458593, /* 2011 */
128'he04ae426ec06e8221101b79102f71823, /* 2012 */
128'hf0ef84ae450d892a08c7df638432478d, /* 2013 */
128'h0000451708a7956325010004d783d39f, /* 2014 */
128'h9a6325010024d783d23ff0ef00055503, /* 2015 */
128'h4511da9ff0ef00448513ffc4059b06a7, /* 2016 */
128'h00004517dca7962300004797d07ff0ef, /* 2017 */
128'h9c23000047974611cf3ff0effd055503, /* 2018 */
128'he29ff0ef854adae5859300004597daa7, /* 2019 */
128'h4515fa65d58300004597256000ef4535, /* 2020 */
128'h00004797240000ef02000513d19ff0ef, /* 2021 */
128'h11230000471727850007d783f9078793, /* 2022 */
128'hcf63278d439cf767879300004797f8f7, /* 2023 */
128'h64428d7fd0ef5f650513000035170087, /* 2024 */
128'h644260e2d47ff06f6105690264a260e2, /* 2025 */
128'hc703f022f406717980826105690264a2, /* 2026 */
128'h00e10f230115c70300e10fa346890105, /* 2027 */
128'h740202f70a63478d00d70e6301e15703, /* 2028 */
128'h885fd06f61455d6505130000351770a2, /* 2029 */
128'h875fd0efe42e5ae5051300003517842a, /* 2030 */
128'h7402d8bff06f614570a265a274028522, /* 2031 */
128'hdc010113ebfff06f614505c170a24190, /* 2032 */
128'h84ae842a232130232291342322813823, /* 2033 */
128'hf0ef22113c2300282180061345818932, /* 2034 */
128'hf0efe802c44a08282040061385a6e52f, /* 2035 */
128'h340323813083f63ff0ef8522002ce90f, /* 2036 */
128'h80822401011322013903228134832301, /* 2037 */
128'h000045974611cb81e8c7d78300004797, /* 2038 */
128'h00efe40611418082cf1ff06fc7458593, /* 2039 */
128'h1001a70300e57763878e1041e7035040, /* 2040 */
128'h60a21007e78310a7a22310e1a0232705, /* 2041 */
128'h80824501808201418d5d910117821502, /* 2042 */
128'h842afc1ff0ef84aae426e822ec061101, /* 2043 */
128'h9101150202f407b33e800793440000ef, /* 2044 */
128'h8082610564a28d0502a7d533644260e2, /* 2045 */
128'h414000ef842af95ff0efe022e4061141, /* 2046 */
128'h640260a202f407b324078793000f47b7, /* 2047 */
128'hec061101808202a7d533014191011502, /* 2048 */
128'h00ef892af63ff0ef84aae04ae426e822, /* 2049 */
128'h543324040413000f443702a485333e20, /* 2050 */
128'h60e2fe856ee3f45ff0ef0405944a0285, /* 2051 */
128'h94b7e426110180826105690264a26442, /* 2052 */
128'h892268048493842ae04aec06e8220098, /* 2053 */
128'hfa1ff0ef41240433854a89260084f363, /* 2054 */
128'h002380826105690264a2644260e2f47d, /* 2055 */
128'hc503100007b7808200054503808200b5, /* 2056 */
128'h01474783100007378082020575130147, /* 2057 */
128'h100007b7808200a70023dfe50207f793, /* 2058 */
128'h8023476d00e78623f800071300078223, /* 2059 */
128'hfc70071300e78623470d0007822300e7, /* 2060 */
128'h1141808200e788230200071300e78423, /* 2061 */
128'h640260a2e50900044503842ae406e022, /* 2062 */
128'h00002797b7f50405fa5ff0ef80820141, /* 2063 */
128'h470397aa973e811100f57713d6c78793, /* 2064 */
128'h808200f5802300e580a30007c7830007, /* 2065 */
128'hfd1ff0efec068121842a002ce8221101, /* 2066 */
128'hf5dff0ef00914503f65ff0ef00814503, /* 2067 */
128'hf0ef00814503fb7ff0ef0ff47513002c, /* 2068 */
128'h6105644260e2f43ff0ef00914503f4bf, /* 2069 */
128'h4461892af406e84aec26f02271798082, /* 2070 */
128'hf81ff0ef0ff57513002c0089553b54e1, /* 2071 */
128'hf0ef00914503f13ff0ef346100814503, /* 2072 */
128'h6145694264e2740270a2fe9410e3f0bf, /* 2073 */
128'h0413892af406e84aec26f02271798082, /* 2074 */
128'hf0ef0ff57513002c0089553354e10380, /* 2075 */
128'h00914503ed1ff0ef346100814503f3ff, /* 2076 */
128'h694264e2740270a2fe9410e3ec9ff0ef, /* 2077 */
128'h4503f13ff0efec06002c110180826145, /* 2078 */
128'h60e2e9fff0ef00914503ea7ff0ef0081, /* 2079 */
128'h7139439ce34787930000479780826105, /* 2080 */
128'h84b2842e892aec4efc06f04af426f822, /* 2081 */
128'hf08fb0efbdc505130000451702b78563, /* 2082 */
128'h744270e2e0a7a42300004797c10d2501, /* 2083 */
128'h0000471757fd8082612169e2790274a2, /* 2084 */
128'h05130000451785ca86260074def72623, /* 2085 */
128'ha92300004797c50d2501fe3fa0efba65, /* 2086 */
128'h05130000351785a6049675634632dca7, /* 2087 */
128'hdaf72a23000047174785cdefd0ef24e5, /* 2088 */
128'h0009099b00c4591be05ff0ef4521b775, /* 2089 */
128'h4503993e003979132487879300003797, /* 2090 */
128'h9c25bf5d2f4010ef854ede7ff0ef0009, /* 2091 */
128'h85aae0221141bf95d687ac2300004797, /* 2092 */
128'hc84fd0efe40621e5051300003517842a, /* 2093 */
128'h64028322f14025730ff0000f0000100f, /* 2094 */
128'h114183020141bce585930000259760a2, /* 2095 */
128'h051300004517f0658593000035974605, /* 2096 */
128'h3517c9112501d47fa0efe022e406d365, /* 2097 */
128'hc34fd06f014160a26402202505130000, /* 2098 */
128'h35974605c28fd0ef2105051300003517, /* 2099 */
128'ha0efaba5051300004517222585930000, /* 2100 */
128'hb7e121a5051300003517c5112501d69f, /* 2101 */
128'h00000517bf8fd0ef0985051300003517, /* 2102 */
128'h00004797cc07a42300004797e9850513, /* 2103 */
128'h479700054863842a90ef90efca07ae23, /* 2104 */
128'h6402408005b3cf81439ccae787930000, /* 2105 */
128'hbb4fd06f014106e505130000351760a2, /* 2106 */
128'hc5112501b72fb0efa505051300004517, /* 2107 */
128'h000035974605bfb91c85051300003517, /* 2108 */
128'h3517c5112501c87fa0ef4501e3c58593, /* 2109 */
128'h0023ee1ff0ef8522b7811c2505130000, /* 2110 */
128'ha001d69ff0efe4062501114190020000, /* 2111 */
128'h471780824501808224050513000f4537, /* 2112 */
128'h869300756513157d631cc22707130000, /* 2113 */
128'h8082953e055e10d00513e30895360017, /* 2114 */
128'hf0efe4328532ec06e822110102b50633, /* 2115 */
128'h8522936ff0ef45816622c509842afd1f, /* 2116 */
128'h000035171141808280826105644260e2, /* 2117 */
128'hc0ef20000537afafd0efe40615c50513, /* 2118 */
128'h45018082450180820141450160a2eadf, /* 2119 */
128'h1141808202f5553347a9b00025738082, /* 2120 */
128'h148505130000351785aa862e86b28736, /* 2121 */
128'h1141a001cbbff0ef4505abefd0efe406, /* 2122 */
128'h408007b3f57ff0efe406952e842ae022, /* 2123 */
128'h80824505808201418d7d640260a29522, /* 2124 */
128'hf406ec26f02271798082450580824505, /* 2125 */
128'h64e2740270a20096186300c684bb842e, /* 2126 */
128'hdfffc0efe432852285b2808261454501, /* 2127 */
128'h450980824509bff92605200404136622, /* 2128 */
128'h80824501808280828082808245098082, /* 2129 */
128'he426e822ec061101bbbff06f80824501, /* 2130 */
128'h986300d5043300d584b3003796934781, /* 2131 */
128'h380380826105450164a2644260e200c7, /* 2132 */
128'h000035176090600c02e8036360980004, /* 2133 */
128'h0000351785a286269fcfd0ef0bc50513, /* 2134 */
128'h715dbf5d0785a0019ecfd0ef0d450513, /* 2135 */
128'hf84ae0a20d4505130000351784aafc26, /* 2136 */
128'h4401892ee45ee486e85aec56f052f44e, /* 2137 */
128'h00003a970c498993000039979c0fd0ef, /* 2138 */
128'h854e4a410d4b0b1300003b170cca8a93, /* 2139 */
128'h994fd0ef855685de00040b9b9a0fd0ef, /* 2140 */
128'h85de986fd0ef854e03271863470187a6, /* 2141 */
128'h040503259963458187a697efd0ef855a, /* 2142 */
128'h964fd0ef0fc5051300003517fd4417e3, /* 2143 */
128'hc613c299863e8a85008706b3a0a94501, /* 2144 */
128'h00858733bf6d07a107056394e390fff7, /* 2145 */
128'h02d60b63fff7c693c31986be8b056390, /* 2146 */
128'h3517926fd0ef0665051300003517058e, /* 2147 */
128'h640660a6557d91afd0ef092505130000, /* 2148 */
128'h61616ba26b426ae27a0279a2794274e2, /* 2149 */
128'h6a05fc56e0d27159b75107a105858082, /* 2150 */
128'hf062f45ef85ae4ceeca6020005138aaa, /* 2151 */
128'h8bb28b2ee46ee86aec66e8caf0a2f486, /* 2152 */
128'h00003c179c4a0a134981b53ff0ef4481, /* 2153 */
128'h00fb0cb300fa8db30034979336cc0c13, /* 2154 */
128'h8a4fd0ef064505130000351703749b63, /* 2155 */
128'h6ce27c027ba26a0669a6694670a67406, /* 2156 */
128'h7ae285567b4264e685da86266da26d42, /* 2157 */
128'hbe1fe0ef842abe7fe0efe47ff06f6165, /* 2158 */
128'h0344f7b3bd5fe0ef892abdbfe0ef8d2a, /* 2159 */
128'h01a4643300a96533010d1d1b0105151b, /* 2160 */
128'h00adb02300acb0238d41910114021502, /* 2161 */
128'h97e20039f7930985ac1ff0ef4521ef81, /* 2162 */
128'he42e7139b7ad0485ab1ff0ef0007c503, /* 2163 */
128'he0ef89aaec4ef04af426f822fc06e032, /* 2164 */
128'h84aab73fe0ef892ab79fe0ef842ab7ff, /* 2165 */
128'h8fc18d450109179b0105151bb6dfe0ef, /* 2166 */
128'h971347818d5d9101178265a266021502, /* 2167 */
128'h70e2744200c79c63974e00e588330037, /* 2168 */
128'hd8dff06f6121863e69e2854e790274a2, /* 2169 */
128'h30238f2900083703e3148ea907856314, /* 2170 */
128'hf426f822fc06e032e42e7139b7f100e8, /* 2171 */
128'hb01fe0ef842ab07fe0ef89aaec4ef04a, /* 2172 */
128'h0105151baf5fe0ef84aaafbfe0ef892a, /* 2173 */
128'h178265a2660215028fc18d450109179b, /* 2174 */
128'h974e00e588330037971347818d5d9101, /* 2175 */
128'h69e2854e790274a270e2744200c79c63, /* 2176 */
128'he3148e8907856314d15ff06f6121863e, /* 2177 */
128'he42e7139b7f100e830238f0900083703, /* 2178 */
128'he0ef89aaec4ef04af426f822fc06e032, /* 2179 */
128'h84aaa83fe0ef892aa89fe0ef842aa8ff, /* 2180 */
128'h8fc18d450109179b0105151ba7dfe0ef, /* 2181 */
128'h971347818d5d9101178265a266021502, /* 2182 */
128'h70e2744200c79c63974e00e588330037, /* 2183 */
128'hc9dff06f6121863e69e2854e790274a2, /* 2184 */
128'h073300083703e31402a686b307856314, /* 2185 */
128'hfc06e032e42e7139b7e100e8302302a7, /* 2186 */
128'h842aa13fe0ef89aaec4ef04af426f822, /* 2187 */
128'ha01fe0ef84aaa07fe0ef892aa0dfe0ef, /* 2188 */
128'h660215028fc18d450109179b0105151b, /* 2189 */
128'h88330037971347818d5d9101178265a2, /* 2190 */
128'h790274a270e2744200c79c63974e00e5, /* 2191 */
128'h4505e111c21ff06f6121863e69e2854e, /* 2192 */
128'h573300083703e31402a6d6b307856314, /* 2193 */
128'hfc06e032e42e7139b7d100e8302302a7, /* 2194 */
128'h842a993fe0ef89aaec4ef04af426f822, /* 2195 */
128'h981fe0ef84aa987fe0ef892a98dfe0ef, /* 2196 */
128'h660215028fc18d450109179b0105151b, /* 2197 */
128'h88330037971347818d5d9101178265a2, /* 2198 */
128'h790274a270e2744200c79c63974e00e5, /* 2199 */
128'h07856314ba1ff06f6121863e69e2854e, /* 2200 */
128'hb7f100e830238f4900083703e3148ec9, /* 2201 */
128'hec4ef04af426f822fc06e032e42e7139, /* 2202 */
128'he0ef892a915fe0ef842a91bfe0ef89aa, /* 2203 */
128'h0109179b0105151b909fe0ef84aa90ff, /* 2204 */
128'h8d5d9101178265a2660215028fc18d45, /* 2205 */
128'h00c79c63974e00e58833003797134781, /* 2206 */
128'h6121863e69e2854e790274a270e27442, /* 2207 */
128'h00083703e3148ee907856314b29ff06f, /* 2208 */
128'hfc06e032e42e7139b7f100e830238f69, /* 2209 */
128'h842a8a3fe0ef89aaec4ef04af426f822, /* 2210 */
128'h891fe0ef84aa897fe0ef892a89dfe0ef, /* 2211 */
128'h660214828fc18cc90109179b0105151b, /* 2212 */
128'h88330037169347018fc59081178265a2, /* 2213 */
128'h790274a270e2744200c71c6396ae00d9, /* 2214 */
128'h00f70533ab1ff06f6121863a69e2854e, /* 2215 */
128'h892ae8ca7159bfc9070500a83023e288, /* 2216 */
128'hfc56e0d2e4cef0a2bc85051300003517, /* 2217 */
128'h8b3289aeec66eca6f486f062f45ef85a, /* 2218 */
128'h3b97bb2a0a1300003a17caffc0ef4401, /* 2219 */
128'h0a93bc2c0c1300003c17bbab8b930000, /* 2220 */
128'h855e85a2fff44493c8dfc0ef85520400, /* 2221 */
128'h179314fd460140900cb3c7ffc0ef8885, /* 2222 */
128'he43285520566186397ce00f905b30036, /* 2223 */
128'h85ce6622c59fc0ef856285a2c61fc0ef, /* 2224 */
128'hfb541be32405e12984aaa17ff0ef854a, /* 2225 */
128'h740670a6c39fc0efbd05051300003517, /* 2226 */
128'h7ba27b427ae26a0669a664e669468526, /* 2227 */
128'hc291876600167693808261656ce27c02, /* 2228 */
128'h7159bfc154fdbf590605e198e3988726, /* 2229 */
128'he8caf0a2af4505130000351784aaeca6, /* 2230 */
128'hf486ec66f062f45ef85afc56e0d2e4ce, /* 2231 */
128'h00003997bd9fc0ef44018ab2892ee86a, /* 2232 */
128'h00003b97ddcb0b1300003b17adc98993, /* 2233 */
128'h00003c97ad4c0c1300003c17ddcb8b93, /* 2234 */
128'h7793ba7fc0ef854e04000a13adcc8c93, /* 2235 */
128'hb95fc0ef856285a2000bbd03cba50014, /* 2236 */
128'h97ca00f485b300361793fffd45134601, /* 2237 */
128'h856685a2b79fc0efe432854e05561c63, /* 2238 */
128'h8d2a92fff0ef852685ca6622b71fc0ef, /* 2239 */
128'hae85051300003517fb441ae32405e529, /* 2240 */
128'h69a6694664e6856a740670a6b51fc0ef, /* 2241 */
128'h61656d426ce27c027ba27b427ae26a06, /* 2242 */
128'hc291876a00167693bf49000b3d038082, /* 2243 */
128'h711db7e15d7db7790605e198e398872a, /* 2244 */
128'he0cae4a6a045051300003517842ae8a2, /* 2245 */
128'h84aefc4eec86e862ec5ef05af456f852, /* 2246 */
128'h9f09091300003917aedfc0ef4c018ab2, /* 2247 */
128'ha00b8b9300003b979f8b0b1300003b17, /* 2248 */
128'h85ce000c099bacbfc0ef854a10000a13, /* 2249 */
128'h8fd9008c1793010c1713abffc0ef855a, /* 2250 */
128'h8fd9020c17138fd9018c17130187e7b3, /* 2251 */
128'h038c17138fd9030c17138fd9028c1713, /* 2252 */
128'h1763972600e406b30036171346018fd9, /* 2253 */
128'hc0ef855e85cea7bfc0efe432854a0556, /* 2254 */
128'he91d89aa831ff0ef852285a66622a73f, /* 2255 */
128'hc0ef9ea5051300003517f94c19e30c05, /* 2256 */
128'h7a4279e2690664a6854e644660e6a53f, /* 2257 */
128'he29ce31c808261256c426be27b027aa2, /* 2258 */
128'h351784aaf4a67119bff159fdb74d0605, /* 2259 */
128'he4d6e8d2eccef0caf8a291a505130000, /* 2260 */
128'h892eec6efc86f06af466f862fc5ee0da, /* 2261 */
128'h900a0a1300003a179fdfc0ef44018b32, /* 2262 */
128'h0c13498507f00b93908c8c9300003c97, /* 2263 */
128'h855208000a93906d0d1300003d1703f0, /* 2264 */
128'h408b873b9c9fc0ef856685a29d1fc0ef, /* 2265 */
128'h86b3003617934601008995b300e99733, /* 2266 */
128'h9a5fc0efe432855205661a6397ca00f4, /* 2267 */
128'hf0ef852685ca662299dfc0ef856a85a2, /* 2268 */
128'h00003517fb541be32405e1398daaf5af, /* 2269 */
128'h74a6856e744670e697dfc0ef91450513, /* 2270 */
128'h7ca27c427be26b066aa66a4669e67906, /* 2271 */
128'he28ce38c008c6663808261096de27d02, /* 2272 */
128'h7119b7f15dfdbfe5e298e398bf610605, /* 2273 */
128'hf0caf8a2834505130000351784aaf4a6, /* 2274 */
128'hf06af466f862fc5ee0dae4d6e8d2ecce, /* 2275 */
128'h3a17917fc0ef44018b32892eec6efc86, /* 2276 */
128'h0b93822c8c9300003c9781aa0a130000, /* 2277 */
128'h820d0d1300003d1703f00c13498507f0, /* 2278 */
128'hc0ef856685a28ebfc0ef855208000a93, /* 2279 */
128'hc793008996b300f997b3408b87bb8e3f, /* 2280 */
128'h00e485b3003617134601fff6c693fff7, /* 2281 */
128'h85a28b7fc0efe432855205661a63974a, /* 2282 */
128'he6cff0ef852685ca66228affc0ef856a, /* 2283 */
128'h051300003517fb5417e32405e1398daa, /* 2284 */
128'h790674a6856e744670e688ffc0ef8265, /* 2285 */
128'h7d027ca27c427be26b066aa66a4669e6, /* 2286 */
128'h0605e194e314008c6663808261096de2, /* 2287 */
128'hf4a67119b7f15dfdbfe5e19ce31cbf61, /* 2288 */
128'heccef0caf8a2746505130000251784aa, /* 2289 */
128'hfc86f06af466f862fc5ee0dae4d6e8d2, /* 2290 */
128'h00002997829fc0ef44018a32892eec6e, /* 2291 */
128'h07f00a93734c0c1300002c1772c98993, /* 2292 */
128'h8c9300002c9703f00b9308100b134d05, /* 2293 */
128'hff4fc0ef856285a2ffcfc0ef854e72ec, /* 2294 */
128'h00ed173300fd17b3408b07bb408a873b, /* 2295 */
128'h8fd5008d16b300fd17b30024079b8f5d, /* 2296 */
128'h8533003616934601fff7c893fff74313, /* 2297 */
128'hfb4fc0efe432854e05461c6396ca00d4, /* 2298 */
128'hf0ef852685ca6622facfc0ef856685a2, /* 2299 */
128'hf8f41be3080007932405ed298daad6af, /* 2300 */
128'h744670e6f88fc0ef7205051300002517, /* 2301 */
128'h7be26b066aa66a4669e6790674a6856e, /* 2302 */
128'h00167813808261096de27d027ca27c42, /* 2303 */
128'he10ce28c85c60008036385be008bea63, /* 2304 */
128'h5dfdbfc5859afe080be385bab7610605, /* 2305 */
128'h6305051300002517892af0ca7119bf75, /* 2306 */
128'hf8a2fc86ec6ef06af466fc5ee8d2ecce, /* 2307 */
128'hc0ef4b81e03289aef862e0dae4d6f4a6, /* 2308 */
128'h8c9300002c97616a0a1300002a17f12f, /* 2309 */
128'h9c3347854da1626d0d1300002d1761ec, /* 2310 */
128'h8b3bee6fc0ef85524401003b949b0177, /* 2311 */
128'h4601fffc4a93edafc0ef856685da0084, /* 2312 */
128'h06f61063974e00e90833003617136782, /* 2313 */
128'heb4fc0ef856a85daebcfc0efe4328552, /* 2314 */
128'h2405e9318b2ac72ff0ef854a85ce6622, /* 2315 */
128'hfafb90e3040007932b85fbb41be38c56, /* 2316 */
128'h744670e6e88fc0ef6205051300002517, /* 2317 */
128'h7be26b066aa66a4669e6790674a6855a, /* 2318 */
128'h00167513808261096de27d027ca27c42, /* 2319 */
128'hb749060500b83023e30c85d6e11185e2, /* 2320 */
128'h84ae892af4cef8cafca67175b7e95b7d, /* 2321 */
128'he0e2e4dee8daecd6f0d2698502000513, /* 2322 */
128'hf0ef8acae032f46ee122e506f86afc66, /* 2323 */
128'h148c0c1300003c174b014a098ba68a6f, /* 2324 */
128'h4d818b2d0d1300003d179c4989934ca1, /* 2325 */
128'h85a6866e04fd966396d6003d96936782, /* 2326 */
128'h8aa68bca4785ed4d842abb6ff0ef854a, /* 2327 */
128'hdd4fc0ef594505130000251702fa1863, /* 2328 */
128'h6ae67a0679a6794674e6640a60aa8522, /* 2329 */
128'h808261497da27d427ce26c066ba66b46, /* 2330 */
128'h910fe0ef842a916fe0efec36b7754a05, /* 2331 */
128'h664267a2904fe0efe42a90afe0efe82a, /* 2332 */
128'h140215028c510106161b8d5d0105151b, /* 2333 */
128'he2880aa7b523000037978d4166e29101, /* 2334 */
128'h078500fb86330006c683018786b34781, /* 2335 */
128'h033df7b3ff9795e300d600230ff6f693, /* 2336 */
128'h8b1b001b079bfcffe0ef4521ef910ba1, /* 2337 */
128'h0d85fbbfe0ef0007c50397ea8b8d0007, /* 2338 */
128'h892af4cef8cafca67175bfb1547dbf05, /* 2339 */
128'he4dee8daecd6f0d269850200051384ae, /* 2340 */
128'h8acae032f46ee122e506f86afc66e0e2, /* 2341 */
128'h0c1300003c174b014a098ba6f85fe0ef, /* 2342 */
128'h790d0d1300002d179c4989934ca102ec, /* 2343 */
128'h866e04fd966396d6003d969367824d81, /* 2344 */
128'h8bca4785ed4d842aa94ff0ef854a85a6, /* 2345 */
128'hc0ef472505130000251702fa18638aa6, /* 2346 */
128'h7a0679a6794674e6640a60aa8522cb2f, /* 2347 */
128'h61497da27d427ce26c066ba66b466ae6, /* 2348 */
128'hd0ef842aff5fd0efec36b7754a058082, /* 2349 */
128'h67a2fe3fd0efe42afe9fd0efe82afeff, /* 2350 */
128'h15028c510106161b8d5d0105151b6642, /* 2351 */
128'hf8a7b823000037978d4166e291011402, /* 2352 */
128'h00fb86330006d683018786b34781e288, /* 2353 */
128'hf7b3ff9795e300d6102392c116c20789, /* 2354 */
128'h001b079beadfe0ef4521ef910ba1033d, /* 2355 */
128'he99fe0ef0007c50397ea8b8d00078b1b, /* 2356 */
128'hecce711980826505bfb1547dbf050d85, /* 2357 */
128'h842a892e962af0caf8a2fff5861389b2, /* 2358 */
128'he4d6e8d2f4a63ae505130000251785aa, /* 2359 */
128'he436fc86ec6ef06af466f862fc5ee0da, /* 2360 */
128'h2b1744854a81e03e00395793bd0fc0ef, /* 2361 */
128'h2c173a2b8b9300002b973a2b0b130000, /* 2362 */
128'h2d173a2c8c9300002c973a2c0c130000, /* 2363 */
128'h3a173aad8d9300002d973aad0d130000, /* 2364 */
128'h0513000025170299f863eaaa0a130000, /* 2365 */
128'h790674a68556744670e6b7efc0ef39e5, /* 2366 */
128'h7d027ca27c427be26b066aa66a4669e6, /* 2367 */
128'h8663b56fc0ef855a85a6808261096de2, /* 2368 */
128'hb44fc0ef8562b4afc0ef855e85ce0009, /* 2369 */
128'h952ff0ef85226582b3cfc0ef856a85e6, /* 2370 */
128'h4c636722010a2783b2cfc0ef856ee129, /* 2371 */
128'h3205051300002517c985000a358302f7, /* 2372 */
128'h0049561300195593008a3783b10fc0ef, /* 2373 */
128'hc0ef30a50513000025179782852295a2, /* 2374 */
128'hc0ef0c25051300002517b7d14a89af2f, /* 2375 */
128'h2f850513000025177179bf890485ae2f, /* 2376 */
128'h0593c45fe0efe44ee84aec26f022f406, /* 2377 */
128'h2517ab6fc0ef2f650513000025170400, /* 2378 */
128'h051300002517aaafc0ef312505130000, /* 2379 */
128'h44850725051300002517a9efc0ef3365, /* 2380 */
128'h008495b3497901f499934441a90fc0ef, /* 2381 */
128'h17e3e73ff0ef24050135853346054685, /* 2382 */
128'h8082614569a2694264e2740270a2ff24, /* 2383 */
128'h1e1346814881470100c5131b46058082, /* 2384 */
128'h97aa000780234000081387f245a901f6, /* 2385 */
128'h0007802397aa0007802397aa00078023, /* 2386 */
128'h267302b71d632705fe0813e397aa387d, /* 2387 */
128'h411686b33e800513c00026f38e15c020, /* 2388 */
128'h02b345bb02c747334000059302a68733, /* 2389 */
128'h2d0505130000251702a7473302a767b3, /* 2390 */
128'hc00028f3c02026f3fac710e39f0fc06f, /* 2391 */
128'hf0ef4505f7bff0ef4501e4061141bf51, /* 2392 */
128'h4521f69ff0ef4511f6fff0ef4509f75f, /* 2393 */
128'h91011502bff1f5dff0ef4541f63ff0ef, /* 2394 */
128'h25016388400007b78082e388400007b7, /* 2395 */
128'h808225016b880007b823400007b78082, /* 2396 */
128'h8d5d0085979b808225017b88400007b7, /* 2397 */
128'h47812581f788400007b78d510106161b, /* 2398 */
128'h3e80079300b76f630007871b40000637, /* 2399 */
128'h07b7ffe537fdc3198b097a98400006b7, /* 2400 */
128'h00076703973600279713808273884000, /* 2401 */
128'h842a4785e406e0221141bfc1f6180785, /* 2402 */
128'h883dfedff0ef0045551b35fd00b7d763, /* 2403 */
128'h640200044503943e2407879300002797, /* 2404 */
128'h579b9d3d00b007b7a45fe06f014160a2, /* 2405 */
128'h65133007071311010085151b67050185, /* 2406 */
128'h458946010034842ec62ae8228fd90585, /* 2407 */
128'h460100344589f55ff0efec06c43e454d, /* 2408 */
128'h56b357610380079385a2f49ff0ef454d, /* 2409 */
128'h60e2fee79ae3058537e100d5802300f5, /* 2410 */
128'hf456f852e0cae4a6711d808261056442, /* 2411 */
128'h84b28aae8b2afc4ee8a2ec86ec5ef05a, /* 2412 */
128'h09b30009041b40000bb7ff860a1b4901, /* 2413 */
128'hf6dff0ef002c03446863008a853b012b, /* 2414 */
128'hed3fd0ef9201854e002c16024084863b, /* 2415 */
128'h7b027aa27a4279e2690664a6644660e6, /* 2416 */
128'hf0ef00c4541b85ce2421808261256be2, /* 2417 */
128'h000025171141bf4d008bb0230921f3bf, /* 2418 */
128'h05130000051782afc0efe406ccc50513, /* 2419 */
128'h40a005b360a200055c63d51f70eff7c5, /* 2420 */
128'h60a2806fc06f0141cc05051300002517, /* 2421 */
128'he06f1d25051300002517b69fe06f0141, /* 2422 */
128'he852ec4ef04af426f822fc067139971f, /* 2423 */
128'h1105051300002517929fe0efe05ae456, /* 2424 */
128'h091300002917400009b7440194ffe0ef, /* 2425 */
128'h0004059b639097ce00341793449510e9, /* 2426 */
128'hdb4f80effe9416e3fadfb0ef0405854a, /* 2427 */
128'h2a97400004b720eb0b1300002b174901, /* 2428 */
128'h49910faa0a1300002a170eaa8a930000, /* 2429 */
128'h608ce09c090585560007c783016907b3, /* 2430 */
128'h0004b823f69fb0ef8622240125816080, /* 2431 */
128'h7413fd391be3f5bfb0ef25818552688c, /* 2432 */
128'h0000071702f7646347190054579b0ff4, /* 2433 */
128'h2517878297ba439c97ba078a68470713, /* 2434 */
128'hac3fe0ef8522f2bfb0ef0ba505130000, /* 2435 */
128'h8522f17fb0ef0b65051300002517a001, /* 2436 */
128'hb0ef0b25051300002517b7f5edbff0ef, /* 2437 */
128'h0b05051300002517bfe9c25ff0eff03f, /* 2438 */
128'h051300002517b7e1de2f80efef1fb0ef, /* 2439 */
128'h00000000bf5dcfdff0efedffb0ef0ae5, /* 2440 */
128'h00000000000000000000000000000000, /* 2441 */
128'h00000000000000000000000000000000, /* 2442 */
128'h00000000000000000000000000000000, /* 2443 */
128'h00000000000000000000000000000000, /* 2444 */
128'h00000000000000000000000000000000, /* 2445 */
128'h00000000000000000000000000000000, /* 2446 */
128'h00000000000000000000000000000000, /* 2447 */
128'h08082828282828080808080808080808, /* 2448 */
128'h08080808080808080808080808080808, /* 2449 */
128'h101010101010101010101010101010a0, /* 2450 */
128'h10101010101004040404040404040404, /* 2451 */
128'h01010101010101010141414141414110, /* 2452 */
128'h10101010100101010101010101010101, /* 2453 */
128'h02020202020202020242424242424210, /* 2454 */
128'h08101010100202020202020202020202, /* 2455 */
128'h00000000000000000000000000000000, /* 2456 */
128'h00000000000000000000000000000000, /* 2457 */
128'h101010101010101010101010101010a0, /* 2458 */
128'h10101010101010101010101010101010, /* 2459 */
128'h01010101010101010101010101010101, /* 2460 */
128'h02010101010101011001010101010101, /* 2461 */
128'h02020202020202020202020202020202, /* 2462 */
128'h02020202020202021002020202020202, /* 2463 */
128'hc1bdceee242070dbe8c7b756d76aa478, /* 2464 */
128'hfd469501a83046134787c62af57c0faf, /* 2465 */
128'h895cd7beffff5bb18b44f7af698098d8, /* 2466 */
128'h49b40821a679438efd9871936b901122, /* 2467 */
128'he9b6c7aa265e5a51c040b340f61e2562, /* 2468 */
128'he7d3fbc8d8a1e68102441453d62f105d, /* 2469 */
128'h455a14edf4d50d87c33707d621e1cde6, /* 2470 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /* 2471 */
128'hfde5380c6d9d61228771f681fffa3942, /* 2472 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /* 2473 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /* 2474 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /* 2475 */
128'hfc93a039ab9423a7432aff97f4292244, /* 2476 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /* 2477 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /* 2478 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /* 2479 */
128'h0c07020d08030e09040f0a05000b0601, /* 2480 */
128'h020f0c090603000d0a0704010e0b0805, /* 2481 */
128'h09020b040d060f08010a030c050e0700, /* 2482 */
128'h6c5f7465735f64735f63736972776f6c, /* 2483 */
128'h6e67696c615f64730000000000006465, /* 2484 */
128'h645f6b6c635f64730000000000000000, /* 2485 */
128'h69747465735f64730000000000007669, /* 2486 */
128'h735f646d635f6473000000000000676e, /* 2487 */
128'h74657365725f64730000000074726174, /* 2488 */
128'h6e636b6c625f64730000000000000000, /* 2489 */
128'h69736b6c625f64730000000000000074, /* 2490 */
128'h6f656d69745f6473000000000000657a, /* 2491 */
128'h655f7172695f64730000000000007475, /* 2492 */
128'h5f63736972776f6c000000000000006e, /* 2493 */
128'h00000000646d635f74726174735f6473, /* 2494 */
128'h746e695f746961775f63736972776f6c, /* 2495 */
128'h000000000067616c665f747075727265, /* 2496 */
128'h00007172695f64735f63736972776f6c, /* 2497 */
128'h695f646d635f64735f63736972776f6c, /* 2498 */
128'h5f63736972776f6c0000000000007172, /* 2499 */
128'h007172695f646e655f617461645f6473, /* 2500 */
128'h00000000bffe9c8800000000bffeaf60, /* 2501 */
128'h004c4b40004c4b400030000020000000, /* 2502 */
128'h6d6d5f6472616f62000000020000ffff, /* 2503 */
128'h00000000bffe4e580064637465675f63, /* 2504 */
128'h00000000bffe4cc600000000bffe4a68, /* 2505 */
128'h00000000000000000000000000000000, /* 2506 */
128'hffffbb42ffffbb3effffbb3effffbb1a, /* 2507 */
128'hffffbb46ffffbb46ffffbb46ffffbb46, /* 2508 */
128'hffffcb68ffffcb62ffffcb5cffffc9b8, /* 2509 */
128'h00000000bffeb28800000000bffeb278, /* 2510 */
128'h00000000bffeb2b000000000bffeb298, /* 2511 */
128'h00000000bffeb2e000000000bffeb2c8, /* 2512 */
128'h00000000bffeb31000000000bffeb2f8, /* 2513 */
128'h00000000bffeb34000000000bffeb328, /* 2514 */
128'h00000000bffeb37000000000bffeb358, /* 2515 */
128'h40040300400402004004010040040000, /* 2516 */
128'h40050000400405004004040140040400, /* 2517 */
128'h30000000000000030000000040050100, /* 2518 */
128'h60000000000000053000000000000001, /* 2519 */
128'h70000000000000027000000000000004, /* 2520 */
128'h00000001400000007000000000000000, /* 2521 */
128'h00000005000000012000000000000006, /* 2522 */
128'h20000000000000020000000040000000, /* 2523 */
128'h00000000100000000000000100000000, /* 2524 */
128'h1e19140f0d0c0a000000000000000000, /* 2525 */
128'h000186a00000271050463c37322d2823, /* 2526 */
128'h017d7840017d784000989680000f4240, /* 2527 */
128'h031975000319750002faf080018cba80, /* 2528 */
128'h02faf08005f5e10002faf080017d7840, /* 2529 */
128'h00000020000000000bebc2000c65d400, /* 2530 */
128'h00000200000001000000008000000040, /* 2531 */
128'h00002000000010000000080000000400, /* 2532 */
128'h0000c000000080000000600000004000, /* 2533 */
128'h37363534333231300002000000010000, /* 2534 */
128'h2043534952776f4c4645444342413938, /* 2535 */
128'h746f6f622d7520646573696d696e696d, /* 2536 */
128'h00000000647261432d445320726f6620, /* 2537 */
128'hfffff9a0fffff9b6fffff9a2fffff98e, /* 2538 */
128'h00000000fffff9dafffff9a0fffff9c8, /* 2539 */
128'he00600003800000039080000edfe0dd0, /* 2540 */
128'h00000000100000001100000028000000, /* 2541 */
128'h0000000000000000a806000059010000, /* 2542 */
128'h00000000010000000000000000000000, /* 2543 */
128'h02000000000000000400000003000000, /* 2544 */
128'h020000000f0000000400000003000000, /* 2545 */
128'h2c6874651b0000001400000003000000, /* 2546 */
128'h007665642d657261622d656e61697261, /* 2547 */
128'h2c687465260000001000000003000000, /* 2548 */
128'h0100000000657261622d656e61697261, /* 2549 */
128'h1a0000000300000000006e65736f6863, /* 2550 */
128'h303140747261752f636f732f2c000000, /* 2551 */
128'h0000003030323531313a303030303030, /* 2552 */
128'h00000000737570630100000002000000, /* 2553 */
128'h01000000000000000400000003000000, /* 2554 */
128'h000000000f0000000400000003000000, /* 2555 */
128'h40787d01380000000400000003000000, /* 2556 */
128'h03000000000000304075706301000000, /* 2557 */
128'h0300000080f0fa024b00000004000000, /* 2558 */
128'h03000000007570635b00000004000000, /* 2559 */
128'h03000000000000006700000004000000, /* 2560 */
128'h0000000079616b6f6b00000005000000, /* 2561 */
128'h7a6874651b0000001300000003000000, /* 2562 */
128'h0000766373697200656e61697261202c, /* 2563 */
128'h34367672720000000b00000003000000, /* 2564 */
128'h0b000000030000000000636466616d69, /* 2565 */
128'h0000393376732c76637369727c000000, /* 2566 */
128'h01000000850000000000000003000000, /* 2567 */
128'h6f72746e6f632d747075727265746e69, /* 2568 */
128'h04000000030000000000000072656c6c, /* 2569 */
128'h0000000003000000010000008f000000, /* 2570 */
128'h1b0000000f00000003000000a0000000, /* 2571 */
128'h000063746e692d7570632c7663736972, /* 2572 */
128'h01000000b50000000400000003000000, /* 2573 */
128'h01000000bb0000000400000003000000, /* 2574 */
128'h01000000020000000200000002000000, /* 2575 */
128'h0030303030303030384079726f6d656d, /* 2576 */
128'h6f6d656d5b0000000700000003000000, /* 2577 */
128'h67000000100000000300000000007972, /* 2578 */
128'h00000040000000000000008000000000, /* 2579 */
128'h0300000000636f730100000002000000, /* 2580 */
128'h03000000020000000000000004000000, /* 2581 */
128'h03000000020000000f00000004000000, /* 2582 */
128'h616972612c6874651b0000001f000000, /* 2583 */
128'h706d697300636f732d657261622d656e, /* 2584 */
128'h000000000300000000007375622d656c, /* 2585 */
128'h303240746e696c6301000000c3000000, /* 2586 */
128'h0d000000030000000000003030303030, /* 2587 */
128'h30746e696c632c76637369721b000000, /* 2588 */
128'hca000000100000000300000000000000, /* 2589 */
128'h07000000010000000300000001000000, /* 2590 */
128'h00000000670000001000000003000000, /* 2591 */
128'h0300000000000c000000000000000002, /* 2592 */
128'h006c6f72746e6f63de00000008000000, /* 2593 */
128'h7075727265746e690100000002000000, /* 2594 */
128'h3030634072656c6c6f72746e6f632d74, /* 2595 */
128'h04000000030000000000000030303030, /* 2596 */
128'h04000000030000000000000000000000, /* 2597 */
128'h0c00000003000000010000008f000000, /* 2598 */
128'h003063696c702c76637369721b000000, /* 2599 */
128'h03000000a00000000000000003000000, /* 2600 */
128'h0b00000001000000ca00000010000000, /* 2601 */
128'h10000000030000000900000001000000, /* 2602 */
128'h000000000000000c0000000067000000, /* 2603 */
128'he8000000040000000300000000000004, /* 2604 */
128'hfb000000040000000300000007000000, /* 2605 */
128'hb5000000040000000300000003000000, /* 2606 */
128'hbb000000040000000300000002000000, /* 2607 */
128'h75626564010000000200000002000000, /* 2608 */
128'h0000304072656c6c6f72746e6f632d67, /* 2609 */
128'h637369721b0000001000000003000000, /* 2610 */
128'h03000000003331302d67756265642c76, /* 2611 */
128'hffff000001000000ca00000008000000, /* 2612 */
128'h00000000670000001000000003000000, /* 2613 */
128'h03000000001000000000000000000000, /* 2614 */
128'h006c6f72746e6f63de00000008000000, /* 2615 */
128'h30303140747261750100000002000000, /* 2616 */
128'h08000000030000000000003030303030, /* 2617 */
128'h03000000003035373631736e1b000000, /* 2618 */
128'h00000010000000006700000010000000, /* 2619 */
128'h04000000030000000010000000000000, /* 2620 */
128'h040000000300000080f0fa024b000000, /* 2621 */
128'h040000000300000000c2010006010000, /* 2622 */
128'h04000000030000000200000014010000, /* 2623 */
128'h04000000030000000100000025010000, /* 2624 */
128'h04000000030000000200000030010000, /* 2625 */
128'h0100000002000000040000003a010000, /* 2626 */
128'h3030303240636d6d2d63736972776f6c, /* 2627 */
128'h10000000030000000000000030303030, /* 2628 */
128'h00000000000000200000000067000000, /* 2629 */
128'h14010000040000000300000000000100, /* 2630 */
128'h25010000040000000300000002000000, /* 2631 */
128'h1b0000000c0000000300000002000000, /* 2632 */
128'h0200000000636d6d2d63736972776f6c, /* 2633 */
128'h406874652d63736972776f6c01000000, /* 2634 */
128'h03000000000000003030303030303033, /* 2635 */
128'h2d63736972776f6c1b0000000c000000, /* 2636 */
128'h5b000000080000000300000000687465, /* 2637 */
128'h0400000003000000006b726f7774656e, /* 2638 */
128'h04000000030000000200000014010000, /* 2639 */
128'h06000000030000000300000025010000, /* 2640 */
128'h0300000000007fe3023e180047010000, /* 2641 */
128'h00000030000000006700000010000000, /* 2642 */
128'h01000000020000000080000000000000, /* 2643 */
128'h303440646e7277682d63736972776f6c, /* 2644 */
128'h0e000000030000000000303030303030, /* 2645 */
128'h6e7277682d63736972776f6c1b000000, /* 2646 */
128'h67000000100000000300000000000064, /* 2647 */
128'h00100000000000000000004000000000, /* 2648 */
128'h09000000020000000200000002000000, /* 2649 */
128'h2300736c6c65632d7373657264646123, /* 2650 */
128'h61706d6f6300736c6c65632d657a6973, /* 2651 */
128'h6f647473006c65646f6d00656c626974, /* 2652 */
128'h65736162656d697400687461702d7475, /* 2653 */
128'h6b636f6c630079636e6575716572662d, /* 2654 */
128'h63697665640079636e6575716572662d, /* 2655 */
128'h75746174730067657200657079745f65, /* 2656 */
128'h2d756d6d006173692c76637369720073, /* 2657 */
128'h230074696c70732d626c740065707974, /* 2658 */
128'h00736c6c65632d747075727265746e69, /* 2659 */
128'h6f72746e6f632d747075727265746e69, /* 2660 */
128'h646e6168702c78756e696c0072656c6c, /* 2661 */
128'h727265746e69007365676e617200656c, /* 2662 */
128'h6572006465646e657478652d73747075, /* 2663 */
128'h616d2c76637369720073656d616e2d67, /* 2664 */
128'h766373697200797469726f6972702d78, /* 2665 */
128'h70732d746e6572727563007665646e2c, /* 2666 */
128'h61702d747075727265746e6900646565, /* 2667 */
128'h0073747075727265746e6900746e6572, /* 2668 */
128'h6f692d6765720074666968732d676572, /* 2669 */
128'h63616d2d6c61636f6c0068746469772d, /* 2670 */
128'h0000000000000000737365726464612d, /* 2671 */
128'h0000000000203a642520656369766544, /* 2672 */
128'h00203a6425206563697665642073250a, /* 2673 */
128'h00000000203a6425206563697665440a, /* 2674 */
128'h000a656369766564206e776f6e6b6e75, /* 2675 */
128'h00000a2973252c73252870756b6f6f6c, /* 2676 */
128'h7265206c616e7265746e692070636864, /* 2677 */
128'h00000000000000000a7025202c726f72, /* 2678 */
128'h5145525f5043484420676e69646e6553, /* 2679 */
128'h4b434120504348440000000a54534555, /* 2680 */
128'h696c432050434844000000000000000a, /* 2681 */
128'h203a7373657264644120504920746e65, /* 2682 */
128'h0000000a64252e64252e64252e642520, /* 2683 */
128'h73657264644120504920726576726553, /* 2684 */
128'h0a64252e64252e64252e642520203a73, /* 2685 */
128'h6120726574756f520000000000000000, /* 2686 */
128'h252e64252e642520203a737365726464, /* 2687 */
128'h6b73616d2074654e0000000a64252e64, /* 2688 */
128'h64252e642520203a7373657264646120, /* 2689 */
128'h697420657361654c000a64252e64252e, /* 2690 */
128'h7364253a6d64253a686425203d20656d, /* 2691 */
128'h3d206e69616d6f44000000000000000a, /* 2692 */
128'h4820746e65696c4300000a2273252220, /* 2693 */
128'h000a22732522203d20656d616e74736f, /* 2694 */
128'h000000000a44455050494b53204b4341, /* 2695 */
128'h000000000000000a4b414e2050434844, /* 2696 */
128'h73657264646120646574736575716552, /* 2697 */
128'h0000000000000a646573756665722073, /* 2698 */
128'h000000000000000a732520726f727245, /* 2699 */
128'h6e6f6974706f2064656c646e61686e75, /* 2700 */
128'h656c646e61686e55000000000a642520, /* 2701 */
128'h64252065646f63706f20504348442064, /* 2702 */
128'h20676e69646e6553000000000000000a, /* 2703 */
128'h000a595245564f435349445f50434844, /* 2704 */
128'h00000000000a29732528726f72726570, /* 2705 */
128'h3a2043414d2073250000000030687465, /* 2706 */
128'h3a583230253a583230253a5832302520, /* 2707 */
128'h000a583230253a583230253a58323025, /* 2708 */
128'h484420646e65732074276e646c756f43, /* 2709 */
128'h206e6f20595245564f43534944205043, /* 2710 */
128'h00000a7325203a732520656369766564, /* 2711 */
128'h5043484420726f6620676e6974696157, /* 2712 */
128'h2020202020202020000a524546464f5f, /* 2713 */
128'h00000000000063250000000000000020, /* 2714 */
128'h0000005832302520000000000000002e, /* 2715 */
128'h00000000732573250000000000000a0a, /* 2716 */
128'h00000000007325203a646c697542202c, /* 2717 */
128'h73257a4820756c250000000000007325, /* 2718 */
128'h0000000000756c250000000000000000, /* 2719 */
128'h0073257a4863252000000000646c252e, /* 2720 */
128'h00000000007325736574794220756c25, /* 2721 */
128'h00003a786c3830250073254269632520, /* 2722 */
128'h000a73252020202000786c6c2a302520, /* 2723 */
128'h000000203a5d64255b6e6f6974636553, /* 2724 */
128'h727265207974696e6173207264646170, /* 2725 */
128'h2c7825286e666c6500000a702520726f, /* 2726 */
128'h000000000a3b29782578302c78257830, /* 2727 */
128'h782578302c302c7825287465736d656d, /* 2728 */
128'h464f5f4f4c43414d00000000000a3b29, /* 2729 */
128'h464f5f494843414d0000000054455346, /* 2730 */
128'h46464f5f524c50540000000054455346, /* 2731 */
128'h46464f5f534346540000000000544553, /* 2732 */
128'h4c5254434f49444d0000000000544553, /* 2733 */
128'h46464f5f534346520054455346464f5f, /* 2734 */
128'h5346464f5f5253520000000000544553, /* 2735 */
128'h46464f5f444142520000000000005445, /* 2736 */
128'h46464f5f524c50520000000000544553, /* 2737 */
128'h000000003f3f3f3f0000000000544553, /* 2738 */
128'h000064252b54455346464f5f524c5052, /* 2739 */
128'h6f746f72502050490000000000000047, /* 2740 */
128'h00000000000000000a50495049203d20, /* 2741 */
128'h6f746f72502050490000000000000054, /* 2742 */
128'h6f746f7250205049000a504745203d20, /* 2743 */
128'h6165682074736574000a505550203d20, /* 2744 */
128'h6e6f6320747365740000000a3a726564, /* 2745 */
128'h6f746f7250205049000a3a73746e6574, /* 2746 */
128'h6f746f7250205049000a504449203d20, /* 2747 */
128'h6f746f725020504900000a5054203d20, /* 2748 */
128'h00000000000000000a50434344203d20, /* 2749 */
128'h6f746f72502050490000000000000036, /* 2750 */
128'h00000000000000000a50565352203d20, /* 2751 */
128'h000a455247203d206f746f7250205049, /* 2752 */
128'h000a505345203d206f746f7250205049, /* 2753 */
128'h00000a4841203d206f746f7250205049, /* 2754 */
128'h000a50544d203d206f746f7250205049, /* 2755 */
128'h5054454542203d206f746f7250205049, /* 2756 */
128'h6f746f72502050490000000000000a48, /* 2757 */
128'h000000000000000a5041434e45203d20, /* 2758 */
128'h6f746f7250205049000000000000004d, /* 2759 */
128'h00000000000000000a504d4f43203d20, /* 2760 */
128'h0a50544353203d206f746f7250205049, /* 2761 */
128'h6f746f72502050490000000000000000, /* 2762 */
128'h00000000000a4554494c504455203d20, /* 2763 */
128'h0a534c504d203d206f746f7250205049, /* 2764 */
128'h6f746f72502050490000000000000000, /* 2765 */
128'h6f746f7270205049000a574152203d20, /* 2766 */
128'h2820646574726f707075736e75203d20, /* 2767 */
128'h79745f6f746f7270000000000a297825, /* 2768 */
128'h0000000000000a78257830203d206570, /* 2769 */
128'h727265746e692064656c646e61686e75, /* 2770 */
128'h414d2070757465530000000a21747075, /* 2771 */
128'h4d454f2049505351000a726464612043, /* 2772 */
128'h0000000000000a7825203d205d64255b, /* 2773 */
128'h00000a786c253a786c25203d2043414d, /* 2774 */
128'h3025203d20737365726464612043414d, /* 2775 */
128'h3230253a783230253a783230253a7832, /* 2776 */
128'h0000000a2e783230253a783230253a78, /* 2777 */
128'h00007f7c5d5b3f3e3d3c3b3a2c2b2a22, /* 2778 */
128'h007f7c5d5b3f3e3d3c3b3a2e2c2b2a22, /* 2779 */
128'h66656463626139383736353433323130, /* 2780 */
128'h72776f6c2f6372730000000000000000, /* 2781 */
128'h00000000000000632e636d6d5f637369, /* 2782 */
128'h61625f6473203d3d20657361625f6473, /* 2783 */
128'h5f63736972776f6c00726464615f6573, /* 2784 */
128'h000a74756f656d6974207325203a6473, /* 2785 */
128'h616d202c6465766f6d65722064726143, /* 2786 */
128'h6425206f74206465676e616863206b73, /* 2787 */
128'h736e692064726143000000000000000a, /* 2788 */
128'h6e616863206b73616d202c6465747265, /* 2789 */
128'h0000000000000a6425206f7420646567, /* 2790 */
128'h25207461206465746165726320636d6d, /* 2791 */
128'h0000000a7825203d2074736f68202c78, /* 2792 */
128'h0000000000006f4e0000000000736559, /* 2793 */
128'h002020203a434d4d0000000052444420, /* 2794 */
128'h00000000000a7325203a656369766544, /* 2795 */
128'h3a4449207265727574636166756e614d, /* 2796 */
128'h0a7825203a4d454f000000000a782520, /* 2797 */
128'h6325203a656d614e0000000000000000, /* 2798 */
128'h0000000000000a206325632563256325, /* 2799 */
128'h00000a6425203a646565705320737542, /* 2800 */
128'h25203a79746963617061432068676948, /* 2801 */
128'h79746963617061430000000000000a73, /* 2802 */
128'h7464695720737542000000000000203a, /* 2803 */
128'h000000000a73257469622d6425203a68, /* 2804 */
128'h0000007825782520000000203a78250a, /* 2805 */
128'h00000000000064735f63736972776f6c, /* 2806 */
128'h0000000065646f6d206e776f6e6b6e55, /* 2807 */
128'h7830203a726f72724520737574617453, /* 2808 */
128'h2074756f656d69540000000a58383025, /* 2809 */
128'h616572206472616320676e6974696177, /* 2810 */
128'h6c69616620636d6d00000000000a7964, /* 2811 */
128'h6d6320706f747320646e6573206f7420, /* 2812 */
128'h6f6c62203a434d4d0000000000000a64, /* 2813 */
128'h20786c257830207265626d756e206b63, /* 2814 */
128'h6c2578302878616d2073646565637865, /* 2815 */
128'h203d3e20434d4d6500000000000a2978, /* 2816 */
128'h726f6620646572697571657220342e34, /* 2817 */
128'h642072657375206465636e61686e6520, /* 2818 */
128'h000000000000000a6165726120617461, /* 2819 */
128'h757320746f6e2073656f642064726143, /* 2820 */
128'h696e6f697469747261702074726f7070, /* 2821 */
128'h656f64206472614300000000000a676e, /* 2822 */
128'h20434820656e6966656420746f6e2073, /* 2823 */
128'h00000a657a69732070756f7267205057, /* 2824 */
128'h636e61686e6520617461642072657355, /* 2825 */
128'h5720434820746f6e2061657261206465, /* 2826 */
128'h696c6120657a69732070756f72672050, /* 2827 */
128'h72617020692550470000000a64656e67, /* 2828 */
128'h505720434820746f6e206e6f69746974, /* 2829 */
128'h67696c6120657a69732070756f726720, /* 2830 */
128'h656f642064726143000000000a64656e, /* 2831 */
128'h6e652074726f7070757320746f6e2073, /* 2832 */
128'h657475626972747461206465636e6168, /* 2833 */
128'h6e65206c61746f54000000000000000a, /* 2834 */
128'h6563786520657a6973206465636e6168, /* 2835 */
128'h20752528206d756d6978616d20736465, /* 2836 */
128'h656f64206472614300000a297525203e, /* 2837 */
128'h6f682074726f7070757320746f6e2073, /* 2838 */
128'h61702064656c6c6f72746e6f63207473, /* 2839 */
128'h6572206574697277206e6f6974697472, /* 2840 */
128'h6e6974746573207974696c696261696c, /* 2841 */
128'h726c61206472614300000000000a7367, /* 2842 */
128'h64656e6f697469747261702079646165, /* 2843 */
128'h206f6e203a434d4d000000000000000a, /* 2844 */
128'h0000000a746e65736572702064726163, /* 2845 */
128'h73657220746f6e206469642064726143, /* 2846 */
128'h20656761746c6f76206f7420646e6f70, /* 2847 */
128'h00000000000000000a217463656c6573, /* 2848 */
128'h7463656c6573206f7420656c62616e75, /* 2849 */
128'h00000000000000000a65646f6d206120, /* 2850 */
128'h646e756f66206473635f747865206f4e, /* 2851 */
128'h78363025206e614d0000000000000a21, /* 2852 */
128'h000000783430257834302520726e5320, /* 2853 */
128'h00000000632563256325632563256325, /* 2854 */
128'h6167656c20434d4d00000064252e6425, /* 2855 */
128'h636167654c2044530000000000007963, /* 2856 */
128'h6867694820434d4d0000000000000079, /* 2857 */
128'h0000297a484d36322820646565705320, /* 2858 */
128'h35282064656570532068676948204453, /* 2859 */
128'h6867694820434d4d000000297a484d30, /* 2860 */
128'h0000297a484d32352820646565705320, /* 2861 */
128'h7a484d32352820323552444420434d4d, /* 2862 */
128'h31524453205348550000000000000029, /* 2863 */
128'h00000000000000297a484d3532282032, /* 2864 */
128'h7a484d30352820353252445320534855, /* 2865 */
128'h35524453205348550000000000000029, /* 2866 */
128'h000000000000297a484d303031282030, /* 2867 */
128'h7a484d30352820303552444420534855, /* 2868 */
128'h31524453205348550000000000000029, /* 2869 */
128'h0000000000297a484d38303228203430, /* 2870 */
128'h0000297a484d30303228203030325348, /* 2871 */
128'h6f6e2064252065636976654420434d4d, /* 2872 */
128'h00000000000000000a646e756f662074, /* 2873 */
128'h00000000434d4d650000000000004453, /* 2874 */
128'h000000297325282000006425203a7325, /* 2875 */
128'h6e656c20656c69460000000000636d6d, /* 2876 */
128'h000000000000000a6425203d20687467, /* 2877 */
128'h0a7325203d202964252c70252835646d, /* 2878 */
128'h666c652064616f6c0000000000000000, /* 2879 */
128'h000a79726f6d656d20524444206f7420, /* 2880 */
128'h2064656c696166206461657220666c65, /* 2881 */
128'h000000646c252065646f632068746977, /* 2882 */
128'h6f6f7420687461702074736575716552, /* 2883 */
128'h00000000000a646c25202e676e6f6c20, /* 2884 */
128'h732522203a717277000000000000002f, /* 2885 */
128'h0a64253d657a69736b636f6c62202c22, /* 2886 */
128'h20657669656365520000000000000000, /* 2887 */
128'h0000000000000a2e646e6520656c6966, /* 2888 */
128'h656c6c6163207172775f656c646e6168, /* 2889 */
128'h206c6167656c6c4900000000000a2e64, /* 2890 */
128'h0a2e6e6f6974617265706f2050544654, /* 2891 */
128'h75716572206e656c0000000000000000, /* 2892 */
128'h6175746361202c5825203d2064657269, /* 2893 */
128'h000000005c2d2f7c000a7825203d206c, /* 2894 */
128'h20646564616f6c2065687420746f6f42, /* 2895 */
128'h6572646461207461206d6172676f7270, /* 2896 */
128'h000000000000000a2e2e2e7025207373, /* 2897 */
128'h445320746e756f6d206f74206c696146, /* 2898 */
128'h000000000000000a2172657669726420, /* 2899 */
128'h6e69206e69622e746f6f622064616f4c, /* 2900 */
128'h0000000000000a79726f6d656d206f74, /* 2901 */
128'h00000000000000006e69622e746f6f62, /* 2902 */
128'h62206e65706f206f742064656c696146, /* 2903 */
128'h206f74206c6961660000000a21746f6f, /* 2904 */
128'h000000000021656c69662065736f6c63, /* 2905 */
128'h6420746e756f6d75206f74206c696166, /* 2906 */
128'h20746f6f622d750a00000000216b7369, /* 2907 */
128'h67617473207473726966206465736162, /* 2908 */
128'h00000a726564616f6c20746f6f622065, /* 2909 */
128'h696166207325206e6f69747265737361, /* 2910 */
128'h696c202c732520656c6966202c64656c, /* 2911 */
128'h206e6f6974636e7566202c642520656e, /* 2912 */
128'h3a4552554c49414600000000000a7325, /* 2913 */
128'h74612078257830203d21207825783020, /* 2914 */
128'h00000a2e782578302074657366666f20, /* 2915 */
128'h7025203d203270202c7025203d203170, /* 2916 */
128'h2020202020202020000000000000000a, /* 2917 */
128'h08080808080808080000000000202020, /* 2918 */
128'h20676e69747465730000000000080808, /* 2919 */
128'h20676e69747365740000000000007525, /* 2920 */
128'h3a4552554c4941460000000000007525, /* 2921 */
128'h64612064616220656c626973736f7020, /* 2922 */
128'h666f20746120656e696c207373657264, /* 2923 */
128'h00000000000a2e782578302074657366, /* 2924 */
128'h7478656e206f7420676e697070696b53, /* 2925 */
128'h000000000000000a2e2e2e7473657420, /* 2926 */
128'h20202020200808080808080808080808, /* 2927 */
128'h08080808080808080808202020202020, /* 2928 */
128'h00000000000820080000000000000008, /* 2929 */
128'h78302073692065676e61722074736574, /* 2930 */
128'h00000000000a70257830206f74207025, /* 2931 */
128'h000000000075252f00752520706f6f4c, /* 2932 */
128'h6441206b637574530000000000000a3a, /* 2933 */
128'h0000203a732520200000007373657264, /* 2934 */
128'h00000a2e656e6f4400000000000a6b6f, /* 2935 */
128'h4d415244206c6174656d20657261420a, /* 2936 */
128'h65747365746d656d00000a7473657420, /* 2937 */
128'h20302e332e34206e6f69737265762072, /* 2938 */
128'h000000000000000a297469622d642528, /* 2939 */
128'h30322029432820746867697279706f43, /* 2940 */
128'h2073656c7261684320323130322d3130, /* 2941 */
128'h000000000000000a2e6e6f62617a6143, /* 2942 */
128'h74207265646e75206465736e6563694c, /* 2943 */
128'h50206c6172656e654720554e47206568, /* 2944 */
128'h65762065736e6563694c2063696c6275, /* 2945 */
128'h0a2e29796c6e6f282032206e6f697372, /* 2946 */
128'h5f676e696b726f770000000000000000, /* 2947 */
128'h20646c25202c424b6425203d20746573, /* 2948 */
128'h6c25202c736e6f697463757274736e69, /* 2949 */
128'h203d20495043202c73656c6379632064, /* 2950 */
128'h00000000000000000a646c252e646c25, /* 2951 */
128'h46454443424139383736353433323130, /* 2952 */
128'h6f57206f6c6c65480000000000000000, /* 2953 */
128'h205d64255b70777300000a0d21646c72, /* 2954 */
128'h73206863746977530000000a5825203d, /* 2955 */
128'h000a58252c5825203d20676e69747465, /* 2956 */
128'h5825203d2064656573206d6f646e6152, /* 2957 */
128'h0a746f6f62204453000000000000000a, /* 2958 */
128'h6f6f6220495053510000000000000000, /* 2959 */
128'h736574204d4152440000000000000a74, /* 2960 */
128'h6f6f6220505446540000000000000a74, /* 2961 */
128'h65742065686361430000000000000a74, /* 2962 */
128'h00000a0d7061727400000000000a7473, /* 2963 */
128'h00000002464c457fcccccccccccccccd, /* 2964 */
128'h1032547698badcfeefcdab8967452301, /* 2965 */
128'h5851f42d4c957f2d1000000020000000, /* 2966 */
128'haaaaaaaaaaaaaaaa5555555555555555, /* 2967 */
128'h00004b4d47545045000000030f060301, /* 2968 */
128'h000000003000000000000000004b4d47, /* 2969 */
128'h00000000ffffffff0000000000000000, /* 2970 */
128'h0000646d635f6473000000000c000000, /* 2971 */
128'h00000000bffeb20800006772615f6473, /* 2972 */
128'h000000000000000000000000cc33aa55, /* 2973 */
128'h00000000000000000000000000000000, /* 2974 */
128'h00000000000000000000000000000000, /* 2975 */
128'h000000002f7c5c2d00000000ffffffff, /* 2976 */
128'hffffffff0000000600000000bffeb3c0, /* 2977 */
128'h00000000bffe70800000000000000000, /* 2978 */
128'h00000000000000000000000000000042, /* 2979 */
128'h00000000000000000000000000000000, /* 2980 */
128'h00000000000000000000000000000000, /* 2981 */
128'h00000000000000000000000000000000, /* 2982 */
128'h00000000000000000000000000000000, /* 2983 */
128'h00000000000000000000000000000000, /* 2984 */
128'h00000000000000000000000000000000, /* 2985 */
128'h00000000000000000000000000000000, /* 2986 */
128'h00000000000000000000000000000000, /* 2987 */
128'h00000000000000000000000000000000, /* 2988 */
128'h00000000000000000000000000000000, /* 2989 */
128'h00000000000000000000000000000000, /* 2990 */
128'h00000000000000000000000000000000, /* 2991 */
128'h00000000000000000000000000000000, /* 2992 */
128'h00000000000000000000000000000000, /* 2993 */
128'h00000000000000000000000000000000, /* 2994 */
128'h00000000000000000000000000000000, /* 2995 */
128'h00000000000000000000000000000000, /* 2996 */
128'h00000000000000000000000000000000, /* 2997 */
128'h00000000000000000000000000000000, /* 2998 */
128'h00000000000000000000000000000000, /* 2999 */
128'h00000000000000000000000000000000, /* 3000 */
128'h00000000000000000000000000000000, /* 3001 */
128'h00000000000000000000000000000000, /* 3002 */
128'h00000000000000000000000000000000, /* 3003 */
128'h00000000000000000000000000000000, /* 3004 */
128'h00000000000000000000000000000000, /* 3005 */
128'h00000000000000000000000000000000, /* 3006 */
128'h00000000000000000000000000000000, /* 3007 */
128'h00000000000000000000000000000000, /* 3008 */
128'h00000000000000000000000000000000, /* 3009 */
128'h00000000000000000000000000000000, /* 3010 */
128'h00000000000000000000000000000000, /* 3011 */
128'h00000000000000000000000000000000, /* 3012 */
128'h00000000000000000000000000000000, /* 3013 */
128'h00000000000000000000000000000000, /* 3014 */
128'h00000000000000000000000000000000, /* 3015 */
128'h00000000000000000000000000000000, /* 3016 */
128'h00000000000000000000000000000000, /* 3017 */
128'h00000000000000000000000000000000, /* 3018 */
128'h00000000000000000000000000000000, /* 3019 */
128'h00000000000000000000000000000000, /* 3020 */
128'h00000000000000000000000000000000, /* 3021 */
128'h00000000000000000000000000000000, /* 3022 */
128'h00000000000000000000000000000000, /* 3023 */
128'h00000000000000000000000000000000, /* 3024 */
128'h00000000000000000000000000000000, /* 3025 */
128'h00000000000000000000000000000000, /* 3026 */
128'h00000000000000000000000000000000, /* 3027 */
128'h00000000000000000000000000000000, /* 3028 */
128'h00000000000000000000000000000000, /* 3029 */
128'h00000000000000000000000000000000, /* 3030 */
128'h00000000000000000000000000000000, /* 3031 */
128'h00000000000000000000000000000000, /* 3032 */
128'h00000000000000000000000000000000, /* 3033 */
128'h00000000000000000000000000000000, /* 3034 */
128'h00000000000000000000000000000000, /* 3035 */
128'h00000000000000000000000000000000, /* 3036 */
128'h00000000000000000000000000000000, /* 3037 */
128'h00000000000000000000000000000000, /* 3038 */
128'h00000000000000000000000000000000, /* 3039 */
128'h00000000000000000000000000000000, /* 3040 */
128'h00000000000000000000000000000000, /* 3041 */
128'h00000000000000000000000000000000, /* 3042 */
128'h00000000000000000000000000000000, /* 3043 */
128'h00000000000000000000000000000000, /* 3044 */
128'h00000000000000000000000000000000, /* 3045 */
128'h00000000000000000000000000000000, /* 3046 */
128'h00000000000000000000000000000000, /* 3047 */
128'h00000000000000000000000000000000, /* 3048 */
128'h00000000000000000000000000000000, /* 3049 */
128'h00000000000000000000000000000000, /* 3050 */
128'h00000000000000000000000000000000, /* 3051 */
128'h00000000000000000000000000000000, /* 3052 */
128'h00000000000000000000000000000000, /* 3053 */
128'h00000000000000000000000000000000, /* 3054 */
128'h00000000000000000000000000000000, /* 3055 */
128'h00000000000000000000000000000000, /* 3056 */
128'h00000000000000000000000000000000, /* 3057 */
128'h00000000000000000000000000000000, /* 3058 */
128'h00000000000000000000000000000000, /* 3059 */
128'h00000000000000000000000000000000, /* 3060 */
128'h00000000000000000000000000000000, /* 3061 */
128'h00000000000000000000000000000000, /* 3062 */
128'h00000000000000000000000000000000, /* 3063 */
128'h00000000000000000000000000000000, /* 3064 */
128'h00000000000000000000000000000000, /* 3065 */
128'h00000000000000000000000000000000, /* 3066 */
128'h00000000000000000000000000000000, /* 3067 */
128'h00000000000000000000000000000000, /* 3068 */
128'h00000000000000000000000000000000, /* 3069 */
128'h00000000000000000000000000000000, /* 3070 */
128'h00000000000000000000000000000000, /* 3071 */
128'h00000000000000000000000000000000, /* 3072 */
128'h00000000000000000000000000000000, /* 3073 */
128'h00000000000000000000000000000000, /* 3074 */
128'h00000000000000000000000000000000, /* 3075 */
128'h00000000000000000000000000000000, /* 3076 */
128'h00000000000000000000000000000000, /* 3077 */
128'h00000000000000000000000000000000, /* 3078 */
128'h00000000000000000000000000000000, /* 3079 */
128'h00000000000000000000000000000000, /* 3080 */
128'h00000000000000000000000000000000, /* 3081 */
128'h00000000000000000000000000000000, /* 3082 */
128'h00000000000000000000000000000000, /* 3083 */
128'h00000000000000000000000000000000, /* 3084 */
128'h00000000000000000000000000000000, /* 3085 */
128'h00000000000000000000000000000000, /* 3086 */
128'h00000000000000000000000000000000, /* 3087 */
128'h00000000000000000000000000000000, /* 3088 */
128'h00000000000000000000000000000000, /* 3089 */
128'h00000000000000000000000000000000, /* 3090 */
128'h00000000000000000000000000000000, /* 3091 */
128'h00000000000000000000000000000000, /* 3092 */
128'h00000000000000000000000000000000, /* 3093 */
128'h00000000000000000000000000000000, /* 3094 */
128'h00000000000000000000000000000000, /* 3095 */
128'h00000000000000000000000000000000, /* 3096 */
128'h00000000000000000000000000000000, /* 3097 */
128'h00000000000000000000000000000000, /* 3098 */
128'h00000000000000000000000000000000, /* 3099 */
128'h00000000000000000000000000000000, /* 3100 */
128'h00000000000000000000000000000000, /* 3101 */
128'h00000000000000000000000000000000, /* 3102 */
128'h00000000000000000000000000000000, /* 3103 */
128'h00000000000000000000000000000000, /* 3104 */
128'h00000000000000000000000000000000, /* 3105 */
128'h00000000000000000000000000000000, /* 3106 */
128'h00000000000000000000000000000000, /* 3107 */
128'h00000000000000000000000000000000, /* 3108 */
128'h00000000000000000000000000000000, /* 3109 */
128'h00000000000000000000000000000000, /* 3110 */
128'h00000000000000000000000000000000, /* 3111 */
128'h00000000000000000000000000000000, /* 3112 */
128'h00000000000000000000000000000000, /* 3113 */
128'h00000000000000000000000000000000, /* 3114 */
128'h00000000000000000000000000000000, /* 3115 */
128'h00000000000000000000000000000000, /* 3116 */
128'h00000000000000000000000000000000, /* 3117 */
128'h00000000000000000000000000000000, /* 3118 */
128'h00000000000000000000000000000000, /* 3119 */
128'h00000000000000000000000000000000, /* 3120 */
128'h00000000000000000000000000000000, /* 3121 */
128'h00000000000000000000000000000000, /* 3122 */
128'h00000000000000000000000000000000, /* 3123 */
128'h00000000000000000000000000000000, /* 3124 */
128'h00000000000000000000000000000000, /* 3125 */
128'h00000000000000000000000000000000, /* 3126 */
128'h00000000000000000000000000000000, /* 3127 */
128'h00000000000000000000000000000000, /* 3128 */
128'h00000000000000000000000000000000, /* 3129 */
128'h00000000000000000000000000000000, /* 3130 */
128'h00000000000000000000000000000000, /* 3131 */
128'h00000000000000000000000000000000, /* 3132 */
128'h00000000000000000000000000000000, /* 3133 */
128'h00000000000000000000000000000000, /* 3134 */
128'h00000000000000000000000000000000, /* 3135 */
128'h00000000000000000000000000000000, /* 3136 */
128'h00000000000000000000000000000000, /* 3137 */
128'h00000000000000000000000000000000, /* 3138 */
128'h00000000000000000000000000000000, /* 3139 */
128'h00000000000000000000000000000000, /* 3140 */
128'h00000000000000000000000000000000, /* 3141 */
128'h00000000000000000000000000000000, /* 3142 */
128'h00000000000000000000000000000000, /* 3143 */
128'h00000000000000000000000000000000, /* 3144 */
128'h00000000000000000000000000000000, /* 3145 */
128'h00000000000000000000000000000000, /* 3146 */
128'h00000000000000000000000000000000, /* 3147 */
128'h00000000000000000000000000000000, /* 3148 */
128'h00000000000000000000000000000000, /* 3149 */
128'h00000000000000000000000000000000, /* 3150 */
128'h00000000000000000000000000000000, /* 3151 */
128'h00000000000000000000000000000000, /* 3152 */
128'h00000000000000000000000000000000, /* 3153 */
128'h00000000000000000000000000000000, /* 3154 */
128'h00000000000000000000000000000000, /* 3155 */
128'h00000000000000000000000000000000, /* 3156 */
128'h00000000000000000000000000000000, /* 3157 */
128'h00000000000000000000000000000000, /* 3158 */
128'h00000000000000000000000000000000, /* 3159 */
128'h00000000000000000000000000000000, /* 3160 */
128'h00000000000000000000000000000000, /* 3161 */
128'h00000000000000000000000000000000, /* 3162 */
128'h00000000000000000000000000000000, /* 3163 */
128'h00000000000000000000000000000000, /* 3164 */
128'h00000000000000000000000000000000, /* 3165 */
128'h00000000000000000000000000000000, /* 3166 */
128'h00000000000000000000000000000000, /* 3167 */
128'h00000000000000000000000000000000, /* 3168 */
128'h00000000000000000000000000000000, /* 3169 */
128'h00000000000000000000000000000000, /* 3170 */
128'h00000000000000000000000000000000, /* 3171 */
128'h00000000000000000000000000000000, /* 3172 */
128'h00000000000000000000000000000000, /* 3173 */
128'h00000000000000000000000000000000, /* 3174 */
128'h00000000000000000000000000000000, /* 3175 */
128'h00000000000000000000000000000000, /* 3176 */
128'h00000000000000000000000000000000, /* 3177 */
128'h00000000000000000000000000000000, /* 3178 */
128'h00000000000000000000000000000000, /* 3179 */
128'h00000000000000000000000000000000, /* 3180 */
128'h00000000000000000000000000000000, /* 3181 */
128'h00000000000000000000000000000000, /* 3182 */
128'h00000000000000000000000000000000, /* 3183 */
128'h00000000000000000000000000000000, /* 3184 */
128'h00000000000000000000000000000000, /* 3185 */
128'h00000000000000000000000000000000, /* 3186 */
128'h00000000000000000000000000000000, /* 3187 */
128'h00000000000000000000000000000000, /* 3188 */
128'h00000000000000000000000000000000, /* 3189 */
128'h00000000000000000000000000000000, /* 3190 */
128'h00000000000000000000000000000000, /* 3191 */
128'h00000000000000000000000000000000, /* 3192 */
128'h00000000000000000000000000000000, /* 3193 */
128'h00000000000000000000000000000000, /* 3194 */
128'h00000000000000000000000000000000, /* 3195 */
128'h00000000000000000000000000000000, /* 3196 */
128'h00000000000000000000000000000000, /* 3197 */
128'h00000000000000000000000000000000, /* 3198 */
128'h00000000000000000000000000000000, /* 3199 */
128'h00000000000000000000000000000000, /* 3200 */
128'h00000000000000000000000000000000, /* 3201 */
128'h00000000000000000000000000000000, /* 3202 */
128'h00000000000000000000000000000000, /* 3203 */
128'h00000000000000000000000000000000, /* 3204 */
128'h00000000000000000000000000000000, /* 3205 */
128'h00000000000000000000000000000000, /* 3206 */
128'h00000000000000000000000000000000, /* 3207 */
128'h00000000000000000000000000000000, /* 3208 */
128'h00000000000000000000000000000000, /* 3209 */
128'h00000000000000000000000000000000, /* 3210 */
128'h00000000000000000000000000000000, /* 3211 */
128'h00000000000000000000000000000000, /* 3212 */
128'h00000000000000000000000000000000, /* 3213 */
128'h00000000000000000000000000000000, /* 3214 */
128'h00000000000000000000000000000000, /* 3215 */
128'h00000000000000000000000000000000, /* 3216 */
128'h00000000000000000000000000000000, /* 3217 */
128'h00000000000000000000000000000000, /* 3218 */
128'h00000000000000000000000000000000, /* 3219 */
128'h00000000000000000000000000000000, /* 3220 */
128'h00000000000000000000000000000000, /* 3221 */
128'h00000000000000000000000000000000, /* 3222 */
128'h00000000000000000000000000000000, /* 3223 */
128'h00000000000000000000000000000000, /* 3224 */
128'h00000000000000000000000000000000, /* 3225 */
128'h00000000000000000000000000000000, /* 3226 */
128'h00000000000000000000000000000000, /* 3227 */
128'h00000000000000000000000000000000, /* 3228 */
128'h00000000000000000000000000000000, /* 3229 */
128'h00000000000000000000000000000000, /* 3230 */
128'h00000000000000000000000000000000, /* 3231 */
128'h00000000000000000000000000000000, /* 3232 */
128'h00000000000000000000000000000000, /* 3233 */
128'h00000000000000000000000000000000, /* 3234 */
128'h00000000000000000000000000000000, /* 3235 */
128'h00000000000000000000000000000000, /* 3236 */
128'h00000000000000000000000000000000, /* 3237 */
128'h00000000000000000000000000000000, /* 3238 */
128'h00000000000000000000000000000000, /* 3239 */
128'h00000000000000000000000000000000, /* 3240 */
128'h00000000000000000000000000000000, /* 3241 */
128'h00000000000000000000000000000000, /* 3242 */
128'h00000000000000000000000000000000, /* 3243 */
128'h00000000000000000000000000000000, /* 3244 */
128'h00000000000000000000000000000000, /* 3245 */
128'h00000000000000000000000000000000, /* 3246 */
128'h00000000000000000000000000000000, /* 3247 */
128'h00000000000000000000000000000000, /* 3248 */
128'h00000000000000000000000000000000, /* 3249 */
128'h00000000000000000000000000000000, /* 3250 */
128'h00000000000000000000000000000000, /* 3251 */
128'h00000000000000000000000000000000, /* 3252 */
128'h00000000000000000000000000000000, /* 3253 */
128'h00000000000000000000000000000000, /* 3254 */
128'h00000000000000000000000000000000, /* 3255 */
128'h00000000000000000000000000000000, /* 3256 */
128'h00000000000000000000000000000000, /* 3257 */
128'h00000000000000000000000000000000, /* 3258 */
128'h00000000000000000000000000000000, /* 3259 */
128'h00000000000000000000000000000000, /* 3260 */
128'h00000000000000000000000000000000, /* 3261 */
128'h00000000000000000000000000000000, /* 3262 */
128'h00000000000000000000000000000000, /* 3263 */
128'h00000000000000000000000000000000, /* 3264 */
128'h00000000000000000000000000000000, /* 3265 */
128'h00000000000000000000000000000000, /* 3266 */
128'h00000000000000000000000000000000, /* 3267 */
128'h00000000000000000000000000000000, /* 3268 */
128'h00000000000000000000000000000000, /* 3269 */
128'h00000000000000000000000000000000, /* 3270 */
128'h00000000000000000000000000000000, /* 3271 */
128'h00000000000000000000000000000000, /* 3272 */
128'h00000000000000000000000000000000, /* 3273 */
128'h00000000000000000000000000000000, /* 3274 */
128'h00000000000000000000000000000000, /* 3275 */
128'h00000000000000000000000000000000, /* 3276 */
128'h00000000000000000000000000000000, /* 3277 */
128'h00000000000000000000000000000000, /* 3278 */
128'h00000000000000000000000000000000, /* 3279 */
128'h00000000000000000000000000000000, /* 3280 */
128'h00000000000000000000000000000000, /* 3281 */
128'h00000000000000000000000000000000, /* 3282 */
128'h00000000000000000000000000000000, /* 3283 */
128'h00000000000000000000000000000000, /* 3284 */
128'h00000000000000000000000000000000, /* 3285 */
128'h00000000000000000000000000000000, /* 3286 */
128'h00000000000000000000000000000000, /* 3287 */
128'h00000000000000000000000000000000, /* 3288 */
128'h00000000000000000000000000000000, /* 3289 */
128'h00000000000000000000000000000000, /* 3290 */
128'h00000000000000000000000000000000, /* 3291 */
128'h00000000000000000000000000000000, /* 3292 */
128'h00000000000000000000000000000000, /* 3293 */
128'h00000000000000000000000000000000, /* 3294 */
128'h00000000000000000000000000000000, /* 3295 */
128'h00000000000000000000000000000000, /* 3296 */
128'h00000000000000000000000000000000, /* 3297 */
128'h00000000000000000000000000000000, /* 3298 */
128'h00000000000000000000000000000000, /* 3299 */
128'h00000000000000000000000000000000, /* 3300 */
128'h00000000000000000000000000000000, /* 3301 */
128'h00000000000000000000000000000000, /* 3302 */
128'h00000000000000000000000000000000, /* 3303 */
128'h00000000000000000000000000000000, /* 3304 */
128'h00000000000000000000000000000000, /* 3305 */
128'h00000000000000000000000000000000, /* 3306 */
128'h00000000000000000000000000000000, /* 3307 */
128'h00000000000000000000000000000000, /* 3308 */
128'h00000000000000000000000000000000, /* 3309 */
128'h00000000000000000000000000000000, /* 3310 */
128'h00000000000000000000000000000000, /* 3311 */
128'h00000000000000000000000000000000, /* 3312 */
128'h00000000000000000000000000000000, /* 3313 */
128'h00000000000000000000000000000000, /* 3314 */
128'h00000000000000000000000000000000, /* 3315 */
128'h00000000000000000000000000000000, /* 3316 */
128'h00000000000000000000000000000000, /* 3317 */
128'h00000000000000000000000000000000, /* 3318 */
128'h00000000000000000000000000000000, /* 3319 */
128'h00000000000000000000000000000000, /* 3320 */
128'h00000000000000000000000000000000, /* 3321 */
128'h00000000000000000000000000000000, /* 3322 */
128'h00000000000000000000000000000000, /* 3323 */
128'h00000000000000000000000000000000, /* 3324 */
128'h00000000000000000000000000000000, /* 3325 */
128'h00000000000000000000000000000000, /* 3326 */
128'h00000000000000000000000000000000, /* 3327 */
128'h00000000000000000000000000000000, /* 3328 */
128'h00000000000000000000000000000000, /* 3329 */
128'h00000000000000000000000000000000, /* 3330 */
128'h00000000000000000000000000000000, /* 3331 */
128'h00000000000000000000000000000000, /* 3332 */
128'h00000000000000000000000000000000, /* 3333 */
128'h00000000000000000000000000000000, /* 3334 */
128'h00000000000000000000000000000000, /* 3335 */
128'h00000000000000000000000000000000, /* 3336 */
128'h00000000000000000000000000000000, /* 3337 */
128'h00000000000000000000000000000000, /* 3338 */
128'h00000000000000000000000000000000, /* 3339 */
128'h00000000000000000000000000000000, /* 3340 */
128'h00000000000000000000000000000000, /* 3341 */
128'h00000000000000000000000000000000, /* 3342 */
128'h00000000000000000000000000000000, /* 3343 */
128'h00000000000000000000000000000000, /* 3344 */
128'h00000000000000000000000000000000, /* 3345 */
128'h00000000000000000000000000000000, /* 3346 */
128'h00000000000000000000000000000000, /* 3347 */
128'h00000000000000000000000000000000, /* 3348 */
128'h00000000000000000000000000000000, /* 3349 */
128'h00000000000000000000000000000000, /* 3350 */
128'h00000000000000000000000000000000, /* 3351 */
128'h00000000000000000000000000000000, /* 3352 */
128'h00000000000000000000000000000000, /* 3353 */
128'h00000000000000000000000000000000, /* 3354 */
128'h00000000000000000000000000000000, /* 3355 */
128'h00000000000000000000000000000000, /* 3356 */
128'h00000000000000000000000000000000, /* 3357 */
128'h00000000000000000000000000000000, /* 3358 */
128'h00000000000000000000000000000000, /* 3359 */
128'h00000000000000000000000000000000, /* 3360 */
128'h00000000000000000000000000000000, /* 3361 */
128'h00000000000000000000000000000000, /* 3362 */
128'h00000000000000000000000000000000, /* 3363 */
128'h00000000000000000000000000000000, /* 3364 */
128'h00000000000000000000000000000000, /* 3365 */
128'h00000000000000000000000000000000, /* 3366 */
128'h00000000000000000000000000000000, /* 3367 */
128'h00000000000000000000000000000000, /* 3368 */
128'h00000000000000000000000000000000, /* 3369 */
128'h00000000000000000000000000000000, /* 3370 */
128'h00000000000000000000000000000000, /* 3371 */
128'h00000000000000000000000000000000, /* 3372 */
128'h00000000000000000000000000000000, /* 3373 */
128'h00000000000000000000000000000000, /* 3374 */
128'h00000000000000000000000000000000, /* 3375 */
128'h00000000000000000000000000000000, /* 3376 */
128'h00000000000000000000000000000000, /* 3377 */
128'h00000000000000000000000000000000, /* 3378 */
128'h00000000000000000000000000000000, /* 3379 */
128'h00000000000000000000000000000000, /* 3380 */
128'h00000000000000000000000000000000, /* 3381 */
128'h00000000000000000000000000000000, /* 3382 */
128'h00000000000000000000000000000000, /* 3383 */
128'h00000000000000000000000000000000, /* 3384 */
128'h00000000000000000000000000000000, /* 3385 */
128'h00000000000000000000000000000000, /* 3386 */
128'h00000000000000000000000000000000, /* 3387 */
128'h00000000000000000000000000000000, /* 3388 */
128'h00000000000000000000000000000000, /* 3389 */
128'h00000000000000000000000000000000, /* 3390 */
128'h00000000000000000000000000000000, /* 3391 */
128'h00000000000000000000000000000000, /* 3392 */
128'h00000000000000000000000000000000, /* 3393 */
128'h00000000000000000000000000000000, /* 3394 */
128'h00000000000000000000000000000000, /* 3395 */
128'h00000000000000000000000000000000, /* 3396 */
128'h00000000000000000000000000000000, /* 3397 */
128'h00000000000000000000000000000000, /* 3398 */
128'h00000000000000000000000000000000, /* 3399 */
128'h00000000000000000000000000000000, /* 3400 */
128'h00000000000000000000000000000000, /* 3401 */
128'h00000000000000000000000000000000, /* 3402 */
128'h00000000000000000000000000000000, /* 3403 */
128'h00000000000000000000000000000000, /* 3404 */
128'h00000000000000000000000000000000, /* 3405 */
128'h00000000000000000000000000000000, /* 3406 */
128'h00000000000000000000000000000000, /* 3407 */
128'h00000000000000000000000000000000, /* 3408 */
128'h00000000000000000000000000000000, /* 3409 */
128'h00000000000000000000000000000000, /* 3410 */
128'h00000000000000000000000000000000, /* 3411 */
128'h00000000000000000000000000000000, /* 3412 */
128'h00000000000000000000000000000000, /* 3413 */
128'h00000000000000000000000000000000, /* 3414 */
128'h00000000000000000000000000000000, /* 3415 */
128'h00000000000000000000000000000000, /* 3416 */
128'h00000000000000000000000000000000, /* 3417 */
128'h00000000000000000000000000000000, /* 3418 */
128'h00000000000000000000000000000000, /* 3419 */
128'h00000000000000000000000000000000, /* 3420 */
128'h00000000000000000000000000000000, /* 3421 */
128'h00000000000000000000000000000000, /* 3422 */
128'h00000000000000000000000000000000, /* 3423 */
128'h00000000000000000000000000000000, /* 3424 */
128'h00000000000000000000000000000000, /* 3425 */
128'h00000000000000000000000000000000, /* 3426 */
128'h00000000000000000000000000000000, /* 3427 */
128'h00000000000000000000000000000000, /* 3428 */
128'h00000000000000000000000000000000, /* 3429 */
128'h00000000000000000000000000000000, /* 3430 */
128'h00000000000000000000000000000000, /* 3431 */
128'h00000000000000000000000000000000, /* 3432 */
128'h00000000000000000000000000000000, /* 3433 */
128'h00000000000000000000000000000000, /* 3434 */
128'h00000000000000000000000000000000, /* 3435 */
128'h00000000000000000000000000000000, /* 3436 */
128'h00000000000000000000000000000000, /* 3437 */
128'h00000000000000000000000000000000, /* 3438 */
128'h00000000000000000000000000000000, /* 3439 */
128'h00000000000000000000000000000000, /* 3440 */
128'h00000000000000000000000000000000, /* 3441 */
128'h00000000000000000000000000000000, /* 3442 */
128'h00000000000000000000000000000000, /* 3443 */
128'h00000000000000000000000000000000, /* 3444 */
128'h00000000000000000000000000000000, /* 3445 */
128'h00000000000000000000000000000000, /* 3446 */
128'h00000000000000000000000000000000, /* 3447 */
128'h00000000000000000000000000000000, /* 3448 */
128'h00000000000000000000000000000000, /* 3449 */
128'h00000000000000000000000000000000, /* 3450 */
128'h00000000000000000000000000000000, /* 3451 */
128'h00000000000000000000000000000000, /* 3452 */
128'h00000000000000000000000000000000, /* 3453 */
128'h00000000000000000000000000000000, /* 3454 */
128'h00000000000000000000000000000000, /* 3455 */
128'h00000000000000000000000000000000, /* 3456 */
128'h00000000000000000000000000000000, /* 3457 */
128'h00000000000000000000000000000000, /* 3458 */
128'h00000000000000000000000000000000, /* 3459 */
128'h00000000000000000000000000000000, /* 3460 */
128'h00000000000000000000000000000000, /* 3461 */
128'h00000000000000000000000000000000, /* 3462 */
128'h00000000000000000000000000000000, /* 3463 */
128'h00000000000000000000000000000000, /* 3464 */
128'h00000000000000000000000000000000, /* 3465 */
128'h00000000000000000000000000000000, /* 3466 */
128'h00000000000000000000000000000000, /* 3467 */
128'h00000000000000000000000000000000, /* 3468 */
128'h00000000000000000000000000000000, /* 3469 */
128'h00000000000000000000000000000000, /* 3470 */
128'h00000000000000000000000000000000, /* 3471 */
128'h00000000000000000000000000000000, /* 3472 */
128'h00000000000000000000000000000000, /* 3473 */
128'h00000000000000000000000000000000, /* 3474 */
128'h00000000000000000000000000000000, /* 3475 */
128'h00000000000000000000000000000000, /* 3476 */
128'h00000000000000000000000000000000, /* 3477 */
128'h00000000000000000000000000000000, /* 3478 */
128'h00000000000000000000000000000000, /* 3479 */
128'h00000000000000000000000000000000, /* 3480 */
128'h00000000000000000000000000000000, /* 3481 */
128'h00000000000000000000000000000000, /* 3482 */
128'h00000000000000000000000000000000, /* 3483 */
128'h00000000000000000000000000000000, /* 3484 */
128'h00000000000000000000000000000000, /* 3485 */
128'h00000000000000000000000000000000, /* 3486 */
128'h00000000000000000000000000000000, /* 3487 */
128'h00000000000000000000000000000000, /* 3488 */
128'h00000000000000000000000000000000, /* 3489 */
128'h00000000000000000000000000000000, /* 3490 */
128'h00000000000000000000000000000000, /* 3491 */
128'h00000000000000000000000000000000, /* 3492 */
128'h00000000000000000000000000000000, /* 3493 */
128'h00000000000000000000000000000000, /* 3494 */
128'h00000000000000000000000000000000, /* 3495 */
128'h00000000000000000000000000000000, /* 3496 */
128'h00000000000000000000000000000000, /* 3497 */
128'h00000000000000000000000000000000, /* 3498 */
128'h00000000000000000000000000000000, /* 3499 */
128'h00000000000000000000000000000000, /* 3500 */
128'h00000000000000000000000000000000, /* 3501 */
128'h00000000000000000000000000000000, /* 3502 */
128'h00000000000000000000000000000000, /* 3503 */
128'h00000000000000000000000000000000, /* 3504 */
128'h00000000000000000000000000000000, /* 3505 */
128'h00000000000000000000000000000000, /* 3506 */
128'h00000000000000000000000000000000, /* 3507 */
128'h00000000000000000000000000000000, /* 3508 */
128'h00000000000000000000000000000000, /* 3509 */
128'h00000000000000000000000000000000, /* 3510 */
128'h00000000000000000000000000000000, /* 3511 */
128'h00000000000000000000000000000000, /* 3512 */
128'h00000000000000000000000000000000, /* 3513 */
128'h00000000000000000000000000000000, /* 3514 */
128'h00000000000000000000000000000000, /* 3515 */
128'h00000000000000000000000000000000, /* 3516 */
128'h00000000000000000000000000000000, /* 3517 */
128'h00000000000000000000000000000000, /* 3518 */
128'h00000000000000000000000000000000, /* 3519 */
128'h00000000000000000000000000000000, /* 3520 */
128'h00000000000000000000000000000000, /* 3521 */
128'h00000000000000000000000000000000, /* 3522 */
128'h00000000000000000000000000000000, /* 3523 */
128'h00000000000000000000000000000000, /* 3524 */
128'h00000000000000000000000000000000, /* 3525 */
128'h00000000000000000000000000000000, /* 3526 */
128'h00000000000000000000000000000000, /* 3527 */
128'h00000000000000000000000000000000, /* 3528 */
128'h00000000000000000000000000000000, /* 3529 */
128'h00000000000000000000000000000000, /* 3530 */
128'h00000000000000000000000000000000, /* 3531 */
128'h00000000000000000000000000000000, /* 3532 */
128'h00000000000000000000000000000000, /* 3533 */
128'h00000000000000000000000000000000, /* 3534 */
128'h00000000000000000000000000000000, /* 3535 */
128'h00000000000000000000000000000000, /* 3536 */
128'h00000000000000000000000000000000, /* 3537 */
128'h00000000000000000000000000000000, /* 3538 */
128'h00000000000000000000000000000000, /* 3539 */
128'h00000000000000000000000000000000, /* 3540 */
128'h00000000000000000000000000000000, /* 3541 */
128'h00000000000000000000000000000000, /* 3542 */
128'h00000000000000000000000000000000, /* 3543 */
128'h00000000000000000000000000000000, /* 3544 */
128'h00000000000000000000000000000000, /* 3545 */
128'h00000000000000000000000000000000, /* 3546 */
128'h00000000000000000000000000000000, /* 3547 */
128'h00000000000000000000000000000000, /* 3548 */
128'h00000000000000000000000000000000, /* 3549 */
128'h00000000000000000000000000000000, /* 3550 */
128'h00000000000000000000000000000000, /* 3551 */
128'h00000000000000000000000000000000, /* 3552 */
128'h00000000000000000000000000000000, /* 3553 */
128'h00000000000000000000000000000000, /* 3554 */
128'h00000000000000000000000000000000, /* 3555 */
128'h00000000000000000000000000000000, /* 3556 */
128'h00000000000000000000000000000000, /* 3557 */
128'h00000000000000000000000000000000, /* 3558 */
128'h00000000000000000000000000000000, /* 3559 */
128'h00000000000000000000000000000000, /* 3560 */
128'h00000000000000000000000000000000, /* 3561 */
128'h00000000000000000000000000000000, /* 3562 */
128'h00000000000000000000000000000000, /* 3563 */
128'h00000000000000000000000000000000, /* 3564 */
128'h00000000000000000000000000000000, /* 3565 */
128'h00000000000000000000000000000000, /* 3566 */
128'h00000000000000000000000000000000, /* 3567 */
128'h00000000000000000000000000000000, /* 3568 */
128'h00000000000000000000000000000000, /* 3569 */
128'h00000000000000000000000000000000, /* 3570 */
128'h00000000000000000000000000000000, /* 3571 */
128'h00000000000000000000000000000000, /* 3572 */
128'h00000000000000000000000000000000, /* 3573 */
128'h00000000000000000000000000000000, /* 3574 */
128'h00000000000000000000000000000000, /* 3575 */
128'h00000000000000000000000000000000, /* 3576 */
128'h00000000000000000000000000000000, /* 3577 */
128'h00000000000000000000000000000000, /* 3578 */
128'h00000000000000000000000000000000, /* 3579 */
128'h00000000000000000000000000000000, /* 3580 */
128'h00000000000000000000000000000000, /* 3581 */
128'h00000000000000000000000000000000, /* 3582 */
128'h00000000000000000000000000000000, /* 3583 */
128'h00000000000000000000000000000000, /* 3584 */
128'h00000000000000000000000000000000, /* 3585 */
128'h00000000000000000000000000000000, /* 3586 */
128'h00000000000000000000000000000000, /* 3587 */
128'h00000000000000000000000000000000, /* 3588 */
128'h00000000000000000000000000000000, /* 3589 */
128'h00000000000000000000000000000000, /* 3590 */
128'h00000000000000000000000000000000, /* 3591 */
128'h00000000000000000000000000000000, /* 3592 */
128'h00000000000000000000000000000000, /* 3593 */
128'h00000000000000000000000000000000, /* 3594 */
128'h00000000000000000000000000000000, /* 3595 */
128'h00000000000000000000000000000000, /* 3596 */
128'h00000000000000000000000000000000, /* 3597 */
128'h00000000000000000000000000000000, /* 3598 */
128'h00000000000000000000000000000000, /* 3599 */
128'h00000000000000000000000000000000, /* 3600 */
128'h00000000000000000000000000000000, /* 3601 */
128'h00000000000000000000000000000000, /* 3602 */
128'h00000000000000000000000000000000, /* 3603 */
128'h00000000000000000000000000000000, /* 3604 */
128'h00000000000000000000000000000000, /* 3605 */
128'h00000000000000000000000000000000, /* 3606 */
128'h00000000000000000000000000000000, /* 3607 */
128'h00000000000000000000000000000000, /* 3608 */
128'h00000000000000000000000000000000, /* 3609 */
128'h00000000000000000000000000000000, /* 3610 */
128'h00000000000000000000000000000000, /* 3611 */
128'h00000000000000000000000000000000, /* 3612 */
128'h00000000000000000000000000000000, /* 3613 */
128'h00000000000000000000000000000000, /* 3614 */
128'h00000000000000000000000000000000, /* 3615 */
128'h00000000000000000000000000000000, /* 3616 */
128'h00000000000000000000000000000000, /* 3617 */
128'h00000000000000000000000000000000, /* 3618 */
128'h00000000000000000000000000000000, /* 3619 */
128'h00000000000000000000000000000000, /* 3620 */
128'h00000000000000000000000000000000, /* 3621 */
128'h00000000000000000000000000000000, /* 3622 */
128'h00000000000000000000000000000000, /* 3623 */
128'h00000000000000000000000000000000, /* 3624 */
128'h00000000000000000000000000000000, /* 3625 */
128'h00000000000000000000000000000000, /* 3626 */
128'h00000000000000000000000000000000, /* 3627 */
128'h00000000000000000000000000000000, /* 3628 */
128'h00000000000000000000000000000000, /* 3629 */
128'h00000000000000000000000000000000, /* 3630 */
128'h00000000000000000000000000000000, /* 3631 */
128'h00000000000000000000000000000000, /* 3632 */
128'h00000000000000000000000000000000, /* 3633 */
128'h00000000000000000000000000000000, /* 3634 */
128'h00000000000000000000000000000000, /* 3635 */
128'h00000000000000000000000000000000, /* 3636 */
128'h00000000000000000000000000000000, /* 3637 */
128'h00000000000000000000000000000000, /* 3638 */
128'h00000000000000000000000000000000, /* 3639 */
128'h00000000000000000000000000000000, /* 3640 */
128'h00000000000000000000000000000000, /* 3641 */
128'h00000000000000000000000000000000, /* 3642 */
128'h00000000000000000000000000000000, /* 3643 */
128'h00000000000000000000000000000000, /* 3644 */
128'h00000000000000000000000000000000, /* 3645 */
128'h00000000000000000000000000000000, /* 3646 */
128'h00000000000000000000000000000000, /* 3647 */
128'h00000000000000000000000000000000, /* 3648 */
128'h00000000000000000000000000000000, /* 3649 */
128'h00000000000000000000000000000000, /* 3650 */
128'h00000000000000000000000000000000, /* 3651 */
128'h00000000000000000000000000000000, /* 3652 */
128'h00000000000000000000000000000000, /* 3653 */
128'h00000000000000000000000000000000, /* 3654 */
128'h00000000000000000000000000000000, /* 3655 */
128'h00000000000000000000000000000000, /* 3656 */
128'h00000000000000000000000000000000, /* 3657 */
128'h00000000000000000000000000000000, /* 3658 */
128'h00000000000000000000000000000000, /* 3659 */
128'h00000000000000000000000000000000, /* 3660 */
128'h00000000000000000000000000000000, /* 3661 */
128'h00000000000000000000000000000000, /* 3662 */
128'h00000000000000000000000000000000, /* 3663 */
128'h00000000000000000000000000000000, /* 3664 */
128'h00000000000000000000000000000000, /* 3665 */
128'h00000000000000000000000000000000, /* 3666 */
128'h00000000000000000000000000000000, /* 3667 */
128'h00000000000000000000000000000000, /* 3668 */
128'h00000000000000000000000000000000, /* 3669 */
128'h00000000000000000000000000000000, /* 3670 */
128'h00000000000000000000000000000000, /* 3671 */
128'h00000000000000000000000000000000, /* 3672 */
128'h00000000000000000000000000000000, /* 3673 */
128'h00000000000000000000000000000000, /* 3674 */
128'h00000000000000000000000000000000, /* 3675 */
128'h00000000000000000000000000000000, /* 3676 */
128'h00000000000000000000000000000000, /* 3677 */
128'h00000000000000000000000000000000, /* 3678 */
128'h00000000000000000000000000000000, /* 3679 */
128'h00000000000000000000000000000000, /* 3680 */
128'h00000000000000000000000000000000, /* 3681 */
128'h00000000000000000000000000000000, /* 3682 */
128'h00000000000000000000000000000000, /* 3683 */
128'h00000000000000000000000000000000, /* 3684 */
128'h00000000000000000000000000000000, /* 3685 */
128'h00000000000000000000000000000000, /* 3686 */
128'h00000000000000000000000000000000, /* 3687 */
128'h00000000000000000000000000000000, /* 3688 */
128'h00000000000000000000000000000000, /* 3689 */
128'h00000000000000000000000000000000, /* 3690 */
128'h00000000000000000000000000000000, /* 3691 */
128'h00000000000000000000000000000000, /* 3692 */
128'h00000000000000000000000000000000, /* 3693 */
128'h00000000000000000000000000000000, /* 3694 */
128'h00000000000000000000000000000000, /* 3695 */
128'h00000000000000000000000000000000, /* 3696 */
128'h00000000000000000000000000000000, /* 3697 */
128'h00000000000000000000000000000000, /* 3698 */
128'h00000000000000000000000000000000, /* 3699 */
128'h00000000000000000000000000000000, /* 3700 */
128'h00000000000000000000000000000000, /* 3701 */
128'h00000000000000000000000000000000, /* 3702 */
128'h00000000000000000000000000000000, /* 3703 */
128'h00000000000000000000000000000000, /* 3704 */
128'h00000000000000000000000000000000, /* 3705 */
128'h00000000000000000000000000000000, /* 3706 */
128'h00000000000000000000000000000000, /* 3707 */
128'h00000000000000000000000000000000, /* 3708 */
128'h00000000000000000000000000000000, /* 3709 */
128'h00000000000000000000000000000000, /* 3710 */
128'h00000000000000000000000000000000, /* 3711 */
128'h00000000000000000000000000000000, /* 3712 */
128'h00000000000000000000000000000000, /* 3713 */
128'h00000000000000000000000000000000, /* 3714 */
128'h00000000000000000000000000000000, /* 3715 */
128'h00000000000000000000000000000000, /* 3716 */
128'h00000000000000000000000000000000, /* 3717 */
128'h00000000000000000000000000000000, /* 3718 */
128'h00000000000000000000000000000000, /* 3719 */
128'h00000000000000000000000000000000, /* 3720 */
128'h00000000000000000000000000000000, /* 3721 */
128'h00000000000000000000000000000000, /* 3722 */
128'h00000000000000000000000000000000, /* 3723 */
128'h00000000000000000000000000000000, /* 3724 */
128'h00000000000000000000000000000000, /* 3725 */
128'h00000000000000000000000000000000, /* 3726 */
128'h00000000000000000000000000000000, /* 3727 */
128'h00000000000000000000000000000000, /* 3728 */
128'h00000000000000000000000000000000, /* 3729 */
128'h00000000000000000000000000000000, /* 3730 */
128'h00000000000000000000000000000000, /* 3731 */
128'h00000000000000000000000000000000, /* 3732 */
128'h00000000000000000000000000000000, /* 3733 */
128'h00000000000000000000000000000000, /* 3734 */
128'h00000000000000000000000000000000, /* 3735 */
128'h00000000000000000000000000000000, /* 3736 */
128'h00000000000000000000000000000000, /* 3737 */
128'h00000000000000000000000000000000, /* 3738 */
128'h00000000000000000000000000000000, /* 3739 */
128'h00000000000000000000000000000000, /* 3740 */
128'h00000000000000000000000000000000, /* 3741 */
128'h00000000000000000000000000000000, /* 3742 */
128'h00000000000000000000000000000000, /* 3743 */
128'h00000000000000000000000000000000, /* 3744 */
128'h00000000000000000000000000000000, /* 3745 */
128'h00000000000000000000000000000000, /* 3746 */
128'h00000000000000000000000000000000, /* 3747 */
128'h00000000000000000000000000000000, /* 3748 */
128'h00000000000000000000000000000000, /* 3749 */
128'h00000000000000000000000000000000, /* 3750 */
128'h00000000000000000000000000000000, /* 3751 */
128'h00000000000000000000000000000000, /* 3752 */
128'h00000000000000000000000000000000, /* 3753 */
128'h00000000000000000000000000000000, /* 3754 */
128'h00000000000000000000000000000000, /* 3755 */
128'h00000000000000000000000000000000, /* 3756 */
128'h00000000000000000000000000000000, /* 3757 */
128'h00000000000000000000000000000000, /* 3758 */
128'h00000000000000000000000000000000, /* 3759 */
128'h00000000000000000000000000000000, /* 3760 */
128'h00000000000000000000000000000000, /* 3761 */
128'h00000000000000000000000000000000, /* 3762 */
128'h00000000000000000000000000000000, /* 3763 */
128'h00000000000000000000000000000000, /* 3764 */
128'h00000000000000000000000000000000, /* 3765 */
128'h00000000000000000000000000000000, /* 3766 */
128'h00000000000000000000000000000000, /* 3767 */
128'h00000000000000000000000000000000, /* 3768 */
128'h00000000000000000000000000000000, /* 3769 */
128'h00000000000000000000000000000000, /* 3770 */
128'h00000000000000000000000000000000, /* 3771 */
128'h00000000000000000000000000000000, /* 3772 */
128'h00000000000000000000000000000000, /* 3773 */
128'h00000000000000000000000000000000, /* 3774 */
128'h00000000000000000000000000000000, /* 3775 */
128'h00000000000000000000000000000000, /* 3776 */
128'h00000000000000000000000000000000, /* 3777 */
128'h00000000000000000000000000000000, /* 3778 */
128'h00000000000000000000000000000000, /* 3779 */
128'h00000000000000000000000000000000, /* 3780 */
128'h00000000000000000000000000000000, /* 3781 */
128'h00000000000000000000000000000000, /* 3782 */
128'h00000000000000000000000000000000, /* 3783 */
128'h00000000000000000000000000000000, /* 3784 */
128'h00000000000000000000000000000000, /* 3785 */
128'h00000000000000000000000000000000, /* 3786 */
128'h00000000000000000000000000000000, /* 3787 */
128'h00000000000000000000000000000000, /* 3788 */
128'h00000000000000000000000000000000, /* 3789 */
128'h00000000000000000000000000000000, /* 3790 */
128'h00000000000000000000000000000000, /* 3791 */
128'h00000000000000000000000000000000, /* 3792 */
128'h00000000000000000000000000000000, /* 3793 */
128'h00000000000000000000000000000000, /* 3794 */
128'h00000000000000000000000000000000, /* 3795 */
128'h00000000000000000000000000000000, /* 3796 */
128'h00000000000000000000000000000000, /* 3797 */
128'h00000000000000000000000000000000, /* 3798 */
128'h00000000000000000000000000000000, /* 3799 */
128'h00000000000000000000000000000000, /* 3800 */
128'h00000000000000000000000000000000, /* 3801 */
128'h00000000000000000000000000000000, /* 3802 */
128'h00000000000000000000000000000000, /* 3803 */
128'h00000000000000000000000000000000, /* 3804 */
128'h00000000000000000000000000000000, /* 3805 */
128'h00000000000000000000000000000000, /* 3806 */
128'h00000000000000000000000000000000, /* 3807 */
128'h00000000000000000000000000000000, /* 3808 */
128'h00000000000000000000000000000000, /* 3809 */
128'h00000000000000000000000000000000, /* 3810 */
128'h00000000000000000000000000000000, /* 3811 */
128'h00000000000000000000000000000000, /* 3812 */
128'h00000000000000000000000000000000, /* 3813 */
128'h00000000000000000000000000000000, /* 3814 */
128'h00000000000000000000000000000000, /* 3815 */
128'h00000000000000000000000000000000, /* 3816 */
128'h00000000000000000000000000000000, /* 3817 */
128'h00000000000000000000000000000000, /* 3818 */
128'h00000000000000000000000000000000, /* 3819 */
128'h00000000000000000000000000000000, /* 3820 */
128'h00000000000000000000000000000000, /* 3821 */
128'h00000000000000000000000000000000, /* 3822 */
128'h00000000000000000000000000000000, /* 3823 */
128'h00000000000000000000000000000000, /* 3824 */
128'h00000000000000000000000000000000, /* 3825 */
128'h00000000000000000000000000000000, /* 3826 */
128'h00000000000000000000000000000000, /* 3827 */
128'h00000000000000000000000000000000, /* 3828 */
128'h00000000000000000000000000000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00000000000000000000000000000000, /* 3840 */
128'h00000000000000000000000000000000, /* 3841 */
128'h00000000000000000000000000000000, /* 3842 */
128'h00000000000000000000000000000000, /* 3843 */
128'h00000000000000000000000000000000, /* 3844 */
128'h00000000000000000000000000000000, /* 3845 */
128'h00000000000000000000000000000000, /* 3846 */
128'h00000000000000000000000000000000, /* 3847 */
128'h00000000000000000000000000000000, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule

