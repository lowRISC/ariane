/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'h01111113fff1011b0000613711249463, /*    1 */
128'h00008297000280e706e2829300008297, /*    2 */
128'h000280e7130505130000051709428293, /*    3 */
128'h81c606130000c617fc05859300000597, /*    4 */
128'h000f4eb701169693fff6869b000066b7, /*    5 */
128'h0085b703fffe8e930005b703240e8e9b, /*    6 */
128'hff81011301b111130110011bfe0e9ae3, /*    7 */
128'h0085b70300e6b0230005b7030006b703, /*    8 */
128'h0185b70300e6b8230105b70300e6b423, /*    9 */
128'hfcc5cce3020686930205859300e6bc23, /*   10 */
128'h40b787b300d787b30147879300000797, /*   11 */
128'h30579073090787930000079700078067, /*   12 */
128'hd90606130000c617830585930000c597, /*   13 */
128'h0005bc230005b8230005b4230005b023, /*   14 */
128'h020004b74ce090effec5c6e302058593, /*   15 */
128'h02000937004484930124a02300100913, /*   16 */
128'h3440297310500073ff24c6e34009091b, /*   17 */
128'hf1402973020004b7fe090ae300897913, /*   18 */
128'h0004a903000920230099093300291913, /*   19 */
128'h4009091b0200093700448493fe091ee3, /*   20 */
128'h1050007334102373342022f3ff24c6e3, /*   21 */
128'h41206d6f7266206f6c6c6548ffdff06f, /*   22 */
128'h617720657361656c502021656e616972, /*   23 */
128'h000a2e2e2e746e656d6f6d2061207469, /*   24 */
128'h00000000000000000000000000000000, /*   25 */
128'h00000000000000000000000000000000, /*   26 */
128'h00000000000000000000000000000000, /*   27 */
128'h00000000000000000000000000000000, /*   28 */
128'h00000000000000000000000000000000, /*   29 */
128'h00000000000000000000000000000000, /*   30 */
128'h00000000000000000000000000000000, /*   31 */
128'hd963454c0005cc635735c28587ae6914, /*   32 */
128'he21c97b6470102a787b30a00051300b7, /*   33 */
128'h853e85b200030563018533038082853a, /*   34 */
128'h510686930000b697b7edfda007138302, /*   35 */
128'h87930000b7976294624707130000b717, /*   36 */
128'h87b30280069302d787bb878d8f9961a7, /*   37 */
128'h47148082853a470100e7956397ba02d7, /*   38 */
128'hf0efe4061141b7f502870713fea68de3, /*   39 */
128'hbfe545018082014160a26108c509fbbf, /*   40 */
128'hf0efe852ec4ef04af426f822fc067139, /*   41 */
128'h0000ba17440144814985892acd31f9bf, /*   42 */
128'hc091553500f44d6300c9278301ca0a13, /*   43 */
128'h61216a4269e2790274a2744270e24501, /*   44 */
128'h67a2ed19f29ff0ef854a85a200308082, /*   45 */
128'h50ef8552000995632485cb990087c783, /*   46 */
128'h0513bf652405192080ef498165224b40, /*   47 */
128'hf2dff0efe42ef406f0227179b7c1fda0, /*   48 */
128'h842aee7ff0ef083065a2c105fda00413, /*   49 */
128'h00f7096300c547030ff007936562e911, /*   50 */
128'h547980826145740270a28522158080ef, /*   51 */
128'hf0efec4ef04af426f822fc067139bfd5, /*   52 */
128'h0000a9970ff00913440184aacd01eebf, /*   53 */
128'h74a2744270e200f4496344dc17498993, /*   54 */
128'hf0ef852685a200308082612169e27902, /*   55 */
128'h85a20127896300c7c78367a2ed09e83f, /*   56 */
128'hb7d924050f2080ef6522410050ef854e, /*   57 */
128'he8dff0ef892eec26f406e84af0227179, /*   58 */
128'he45ff0ef84aa85ca0030c11dfda00413, /*   59 */
128'h118505130000a517864a608ced01842a, /*   60 */
128'h740270a285220b4080ef65223d2050ef, /*   61 */
128'hf406ec26f022717980826145694264e2, /*   62 */
128'h85a6842ac11dfda00413e47ff0ef84ae, /*   63 */
128'hcf63445c39a050ef0f0505130000a517, /*   64 */
128'h543507a080ef0ee505130000a51700f4, /*   65 */
128'h003085228082614564e2740270a28522, /*   66 */
128'h04e080ef6522f565842adcfff0ef85a6, /*   67 */
128'h5479fcf71be30ff0079300c7c70367a2, /*   68 */
128'he50965a2de1ff0eff406e42e7179bfc1, /*   69 */
128'hf96dd97ff0ef08308082614570a24501, /*   70 */
128'he42eec064108842ae8221101bfc56562, /*   71 */
128'h852200030e6302053303c919db9ff0ef, /*   72 */
128'h60e2fda005138302610560e265a26442, /*   73 */
128'h0000b7977139bfdd4501808261056442, /*   74 */
128'h04130000b417f426f822639c29c78793, /*   75 */
128'h043b840d8c053a2484930000b4973aa4, /*   76 */
128'h892afc06e852ec4ef04a0280079302f4, /*   77 */
128'h942602f4043302ea0a130000aa1789ae, /*   78 */
128'h69e2790274a2744270e2450100849b63, /*   79 */
128'h296050ef855285ca6090808261216a42, /*   80 */
128'hbfc902848493c5016a3060ef854a608c, /*   81 */
128'hb7e16522f569cdbff0ef852685ce0030, /*   82 */
128'h84b68432e42efc06f04af426f8227139, /*   83 */
128'hcb5ff0ef083065a2c115cf7ff0ef893a, /*   84 */
128'h70e2978285a2615c862686ca6562e519, /*   85 */
128'hbfc5fda0051380826121790274a27442, /*   86 */
128'h84b68432e42efc06f04af426f8227139, /*   87 */
128'hc75ff0ef083065a2c115cb7ff0ef893a, /*   88 */
128'h70e2978285a2655c862686ca6562e519, /*   89 */
128'hbfc5fda0051380826121790274a27442, /*   90 */
128'hc7dff0ef84b2e42ef822fc06f4267139, /*   91 */
128'h701ce509c39ff0ef842a083065a2c105, /*   92 */
128'h8082612174a2744270e2978285a66562, /*   93 */
128'h2785c3190017f713419cbfcdfda00513, /*   94 */
128'hd71b8e5927a106220086571b419cc19c, /*   95 */
128'h0ff77713c19c0087d7138ed906a20086, /*   96 */
128'h122300d5112300c510238fd90087979b, /*   97 */
128'hf022f4067179419c80820005132300f5, /*   98 */
128'h419c00f510230457879b6785c19c27d1, /*   99 */
128'h0087979b0ff777130087d713c632842a, /*  100 */
128'hc4360509084c57fd460900f11a238fd9, /*  101 */
128'h0513016105934609791060ef00f11b23, /*  102 */
128'h00041323082c462147c1783060ef0044, /*  103 */
128'h00f404a347c576f060efec3e00840513, /*  104 */
128'h759060ef00c4051300041523006c4611, /*  105 */
128'h0144069374d060ef01040513002c4611, /*  106 */
128'hfed79ce39f31ffe7d6030789470187a2, /*  107 */
128'h9fb94107d71b9fb9934117424107579b, /*  108 */
128'h80826145740270a200f41523fff7c793, /*  109 */
128'h97ba46a167856398138787930000b797, /*  110 */
128'hc7bb27850077e793fff6079b8007bc23, /*  111 */
128'h3823973e678500f547636805450102d7, /*  112 */
128'h010686bb0035169b0005b883808280c7, /*  113 */
128'he0221141bff105a125050116b02396ba, /*  114 */
128'hfa5ff0efe406450185aa86220005841b, /*  115 */
128'hec26f022717980820141640260a28522, /*  116 */
128'h699060efe436f4064619051984b2842a, /*  117 */
128'h162347a168d060ef85b64619852266a2, /*  118 */
128'h614564e200e4859b70a27402852200f4, /*  119 */
128'h3a8130236785737dc5010113fadff06f, /*  120 */
128'h3931342338913c233a11342339213823, /*  121 */
128'h377134233761382337513c2339413023, /*  122 */
128'h3507879335a1382335913c2337813023, /*  123 */
128'hce042023d00007b7943e747d978a911a, /*  124 */
128'hd0040023f0040023e0040023ca040b23, /*  125 */
128'ha51785aa00e7ea63892a5800073797aa, /*  126 */
128'h00054703a0017ad040efd32505130000, /*  127 */
128'h970a3507871374fd678526f711634789, /*  128 */
128'hcb848b13970a350787139abacd848a93, /*  129 */
128'h9c3a9b3a49818a368cb28baed0048c13, /*  130 */
128'hc7830015cd03013907b395ca0f098593, /*  131 */
128'h869b01a989bb058902a0071329890f07, /*  132 */
128'h24e78163471904f76b6326e78d630007, /*  133 */
128'hcc848513470d2ae78963470502f76263, /*  134 */
128'h40efe32505130000a51785b622e78963, /*  135 */
128'hfee794e3473d22e785634731b77d7250, /*  136 */
128'h953e866ae0048513978a350787936785, /*  137 */
128'h03600713b759e00d0023553060ef9d22, /*  138 */
128'h22e780630330071300f76e6322e78363, /*  139 */
128'haad94605cb648513fae798e303500713, /*  140 */
128'hf8e79ce30ff0071324e7856303800713, /*  141 */
128'h24e781630007859b747d471500614783, /*  142 */
128'h000ca7833ae79d63470938e781634719, /*  143 */
128'h05134985978a350a87936a8516079263, /*  144 */
128'h60ef013ca023953e461101090593ce44, /*  145 */
128'h01490593ce840513978a350a87934d70, /*  146 */
128'hc08505130000a5174c1060ef953e4611, /*  147 */
128'h978a350a879365d040efde0254e25a52, /*  148 */
128'h447060ef854a55fd4619993ecf840913, /*  149 */
128'h879346f115231350079300f103a3478d, /*  150 */
128'h85a6460594becb740493c2a6978a350a, /*  151 */
128'h06a30320079346f060efc0d246c10513, /*  152 */
128'h4a1195becf040593978a350a879346f1, /*  153 */
128'h079344b060ef4741072346f105134611, /*  154 */
128'hcf440593978a350a879346f109a30360, /*  155 */
128'h429060ef47410a2347510513461195be, /*  156 */
128'h03a346f10ca347b1051385a6460557fd, /*  157 */
128'h06131020079340f060ef47310d230001, /*  158 */
128'h07933a9060efde3e37a1051345810f00, /*  159 */
128'h3961051385de4799464136f11d231010, /*  160 */
128'h13232637879377e13e1060ef36f10e23, /*  161 */
128'h350a879346f1142335378793679946f1, /*  162 */
128'h0440061304300693943ecec40413978a, /*  163 */
128'h85a2460156fdba1ff0ef3721051385a2, /*  164 */
128'h0e8885de86ca5672bd5ff0ef35e10513, /*  165 */
128'h3a0134033a813083911a6305cebff0ef, /*  166 */
128'h38013a03388139833901390339813483, /*  167 */
128'h36013c0336813b8337013b0337813a83, /*  168 */
128'h851380823b01011335013d0335813c83, /*  169 */
128'ha00d953e978a3507879367854611cd04, /*  170 */
128'h953e866af0048513978a350787936785, /*  171 */
128'h85564611b39df00d0023333060ef9d22, /*  172 */
128'h87936785bfdd855a4611bbb1325060ef, /*  173 */
128'h309060ef4611953ece048513978a3507, /*  174 */
128'h00f40123ce14478300f401a3ce044783, /*  175 */
128'h00f40023ce34478300f400a3ce244783, /*  176 */
128'h866ab759cc048513bb29cef42023401c, /*  177 */
128'h2783b311d00d00232d1060ef9d228562, /*  178 */
128'h0000a51700fa2023478512079a63000a, /*  179 */
128'h0e8801090593461145f040efa1c50513, /*  180 */
128'hcb840513978a3504879364852a5060ef, /*  181 */
128'h3531470328d060ef014905934611953e, /*  182 */
128'h0000a517350145833511460335214683, /*  183 */
128'h00a146833501578341f040ef9ec50513, /*  184 */
128'h35215783dcf71e230000b71700914603, /*  185 */
128'h0000b7179ec505130000a51700814583, /*  186 */
128'h01b147033eb040ef00b14703dcf71323, /*  187 */
128'h0000a517018145830191460301a14683, /*  188 */
128'h01214683013147033cf040ef9ec50513, /*  189 */
128'h9f0505130000a5170101458301114603, /*  190 */
128'h05130000a51755c2010157833b3040ef, /*  191 */
128'hb71701215783d6f713230000b7179fe5, /*  192 */
128'hf6bb02f5d63b03c00793d4f71e230000, /*  193 */
128'h02f5d5bbe107879b678502f6763b02f5, /*  194 */
128'h95bee0040593978a35048793373040ef, /*  195 */
128'h3504879335b040ef9d8505130000a517, /*  196 */
128'h9d0505130000a51795be978af0040593, /*  197 */
128'h40ef9da505130000a517b501343040ef, /*  198 */
128'h20234785de0796e3000a2783bbcd3350, /*  199 */
128'ha517319040ef9ce505130000a51700fa, /*  200 */
128'h35078793678530d040ef9d2505130000, /*  201 */
128'h9d8505130000a51795be978ad0040593, /*  202 */
128'hb35d2e9040ef9de505130000a517bf45, /*  203 */
128'hf852fc4ee0cae4a6e8a2ec86711d737d, /*  204 */
128'h6a859f2505130000a517911a89aaf456, /*  205 */
128'h0493978a020a8793747d2c1040efca02, /*  206 */
128'hb7970a9060ef852655fd461994beff84, /*  207 */
128'hc83e4a05fef40913439cb02787930000, /*  208 */
128'h993e978a020a879312f11d2313500793, /*  209 */
128'h07930cb060ef014107a31a68460585ca, /*  210 */
128'h020a879312f10f23479112f10ea30370, /*  211 */
128'h60ef13f10513461195beff040593978a, /*  212 */
128'h14f101a314510513460585ca57fd0a70, /*  213 */
128'h0fc0079308d060ef000107a315410223, /*  214 */
128'h027060efca3e04a1051345810f000613, /*  215 */
128'h05134641479985ce04f1152310100793, /*  216 */
128'h2637879377e105f060ef04f106230661, /*  217 */
128'h879312f11c2335378793679912f11b23, /*  218 */
128'h06930421051385a2943e1451978a020a, /*  219 */
128'h02e1051385a2821ff0ef044006130430, /*  220 */
128'h85ce86a610084652855ff0ef460156fd, /*  221 */
128'h64a66446450160e6911a630596bff0ef, /*  222 */
128'ha51785aa808261257aa27a4279e26906, /*  223 */
128'h34238101011319d0406f8e2505130000, /*  224 */
128'h34237d2138237c913c237e8130237e11, /*  225 */
128'h893689b2e04605a1051384aa71597d31, /*  226 */
128'h101867857bc060efd602e83eec3ae442, /*  227 */
128'h943e7fc404136762747d97ba81078793, /*  228 */
128'hf8aff0efd64e0521051385a2864a86ba, /*  229 */
128'hf0ef03e10513863e86c285a267c26822, /*  230 */
128'h8cfff0ef86c685a6180856326882fbaf, /*  231 */
128'h7d8134837e01340345017e8130836165, /*  232 */
128'h716d80827f0101137c8139837d013903, /*  233 */
128'h003547830045480300554883e222e606, /*  234 */
128'ha597842a000546030015468300254703, /*  235 */
128'h40ef832505130000a517832585930000, /*  236 */
128'ha597860ac10d842adedff0ef85220d50, /*  237 */
128'h40ef83a505130000a517812585930000, /*  238 */
128'h0000a51780826151641260b285220b50, /*  239 */
128'h097040ef9e07ae230000b79785450513, /*  240 */
128'hf85afc56e0d2e4ceeca6f0a27159b7cd, /*  241 */
128'h8a2ae46ee8caf486e86aec66f062f45e, /*  242 */
128'h540a8a930000aa974401ff05049389ae, /*  243 */
128'h0000ac1706000b93828b0b130000ab17, /*  244 */
128'hfff58d1b824c8c930000ac97834c0c13, /*  245 */
128'h6a0669a6694664e6740670a603344163, /*  246 */
128'h61656da26d426ce27c027ba27b427ae2, /*  247 */
128'h017040ef855ae7a9c42900f477938082, /*  248 */
128'hfe05879b0007c583012487b34dc14901, /*  249 */
128'h09057f8040ef856602fbe2630ff7f793, /*  250 */
128'h7e6040ef314505130000a517ffb912e3, /*  251 */
128'hb7c57d8040ef8562a0317e0040ef8556, /*  252 */
128'h40ef7b250513000095170104c583dbe5, /*  253 */
128'h00f979134d81fffd4913028d1d637c40, /*  254 */
128'h855aff2dcce32d857ae040ef8556a029, /*  255 */
128'h00f45b630009079bff0479137a2040ef, /*  256 */
128'h0485240578a040ef2b8505130000a517, /*  257 */
128'hf793fe05879b0007c583012a07b3b781, /*  258 */
128'hb7e9090576a040ef856600fbe7630ff7, /*  259 */
128'he44ee84aec267179bfdd760040ef8562, /*  260 */
128'h86930000a697893289ae84b6f022f406, /*  261 */
128'h0000971772c6869300009697c509fce6, /*  262 */
128'h854a85a67246061300009617bfc70713, /*  263 */
128'h85bb00955d6300098f63842a6e2040ef, /*  264 */
128'h40ef954a70c606130000961786ce40a4, /*  265 */
128'hffd4841b00f44463ffe4879b9c296c40, /*  266 */
128'h27c060ef6dc585930000959700890533, /*  267 */
128'h8082614569a2694264e2854a740270a2, /*  268 */
128'h0613002c7115f73ff06f4581862e86b2, /*  269 */
128'h00009517002cfebff0efed8645050c80, /*  270 */
128'h8082612d450160ee6ae040ef6c450513, /*  271 */
128'h47b704a76963862e9ff787133b9ad7b7, /*  272 */
128'hf7633e70079304a7676323f78713000f, /*  273 */
128'h6e8707130000a7173e80079346890ca7, /*  274 */
128'he426e822ec0600074903e04a97361101, /*  275 */
128'h951785aa690264a260e2644202091663, /*  276 */
128'h8793468164a0406f610566a505130000, /*  277 */
128'h02f57433bf7d240787934685b7d9a007, /*  278 */
128'h0287e66347293e800793c02102f555b3, /*  279 */
128'h0287746306300713c70502f4773347a9, /*  280 */
128'h0324341302e4743302f457b306400713, /*  281 */
128'h5433bfc102e45433a039943e00144413, /*  282 */
128'h40ef84b26145051300009517f86102f4, /*  283 */
128'h40ef60a505130000951785a2c8015e40, /*  284 */
128'h9517690264a285ca862660e264425d40, /*  285 */
128'h951785aa5ba0406f61055fa505130000, /*  286 */
128'h481958d94781862eb78d5ca505130000, /*  287 */
128'h1782cd8500e555b303c6871b02f886bb, /*  288 */
128'he42697c211015f6808130000a8179381, /*  289 */
128'h60e26442e495e04ae822ec060007c483, /*  290 */
128'h61055aa505130000951785aa690264a2, /*  291 */
128'h0000951785aafb079de327855620406f, /*  292 */
128'hfff7c79300e797b357fdb7f559450513, /*  293 */
128'h03b6869b02f5053347a9c10d44018d7d, /*  294 */
128'hf46300e45433942a47a500d414334405, /*  295 */
128'h89325425051300009517058514590087, /*  296 */
128'h538505130000951785a2c801512040ef, /*  297 */
128'h64a2690285a6864a60e26442502040ef, /*  298 */
128'h71514e80406f61055405051300009517, /*  299 */
128'he96ae5cee9caf1a202c7073b8cbaed66, /*  300 */
128'he56ef162f55ef95afd56e1d2eda6f586, /*  301 */
128'h00e7f66384368d3289ae892a04000793, /*  302 */
128'hdcbb4cc1000c956302ccdcbb04000c93, /*  303 */
128'h0017849be03e020d1a13001d179b03ac, /*  304 */
128'h4e8b0b1300009b1703810a93020a5a13, /*  305 */
128'h3d8c0c1300008c17450b8b9300009b97, /*  306 */
128'h6a0e69ae694e64ee740e70ae4501e00d, /*  307 */
128'h616d6daa6d4a6cea7c0a7baa7b4a7aea, /*  308 */
128'h446040ef4a4505130000951785ca8082, /*  309 */
128'h470186ce000c8d9b008cf46300040d9b, /*  310 */
128'h971305b66c630007061b430948a14811, /*  311 */
128'h06bb0d9de66399ba034707339301020d, /*  312 */
128'h415705bb0006861b02e00813875603bd, /*  313 */
128'h05130000951785d6963e011c0ac5ed63, /*  314 */
128'h043b66a23ea040effa060c23e43645e5, /*  315 */
128'h557dd135022070ef99369281168241b4, /*  316 */
128'h260195d6002715934290030d1b63b795, /*  317 */
128'hec42f046f41a855a658292011602c190, /*  318 */
128'h96d27322674266a23ae040efe436e83a, /*  319 */
128'h15936290011d1863bf85686278820705, /*  320 */
128'h0006d603006d1c63bfc1e19095d60037, /*  321 */
128'hbf6500c590239241164295d600171593, /*  322 */
128'h00c580230ff6761300ea85b30006c603, /*  323 */
128'h6ae32705672204e070efe43a855eb75d, /*  324 */
128'h053300074583bfdd4701bf1d3cfdfe97, /*  325 */
128'h0185959bc519097575130005450300bc, /*  326 */
128'hbf390705010700230005d4634185d59b, /*  327 */
128'h8082e21c00b7f4634501918187aa1582, /*  328 */
128'h668312b7f46304000793bfd58f8d2505, /*  329 */
128'h10e69c63478957f70713464c47370005, /*  330 */
128'h07930385570310e69763470900454683, /*  331 */
128'h9a93fc567100f0a202f7073371590380, /*  332 */
128'hf45ef85ae0d2e4cee8caeca6f4860205, /*  333 */
128'h478d9722020ada93e46ee86aec66f062, /*  334 */
128'h9b974b054a01942a84aa892e06eae663, /*  335 */
128'h9c97352c0c1300009c17312b8b930000, /*  336 */
128'h478100fa64630384d783332c8c930000, /*  337 */
128'h855e85d2cbc1741c09679b63401ca835, /*  338 */
128'h3d03640c04098d6302043983272040ef, /*  339 */
128'h9517864a02bafa6395ce00b48db30184, /*  340 */
128'h740670a6478d24c040ef2d2505130000, /*  341 */
128'h7c027ba27b427ae26a0669a6694664e6, /*  342 */
128'h85ea866e80826165853e6da26d426ce2, /*  343 */
128'h60ef856a85ee864e21e040ef856686ce, /*  344 */
128'h01843d030337f163701c028439830660, /*  345 */
128'h1f6040ef856285ea9d3e864e40f989b3, /*  346 */
128'h038404132a057ed050ef856a4581864e, /*  347 */
128'h05378082057e45058082853e4785bf99, /*  348 */
128'h157d631c354707130000a71780824000, /*  349 */
128'h20000537e30895360017869300756513, /*  350 */
128'h8207871367858082953e057e450597aa, /*  351 */
128'h95178087871308a74463862a0ce50763, /*  352 */
128'h079b04c7496306e60b63272505130000, /*  353 */
128'h87936785c3ad24e50513000095178006, /*  354 */
128'h77fd04c7c9632ce505130000951787f7, /*  355 */
128'h2c058593000095979e3d11417c07879b, /*  356 */
128'h60a2124040efe4062b8505130000a517, /*  357 */
128'h81078713808201412a8505130000a517, /*  358 */
128'h8187879300e60a632205051300009517, /*  359 */
128'h87138082faf612e32205051300009517, /*  360 */
128'h4963fee609e323e50513000095178307, /*  361 */
128'hbfe921a50513000095178287879300c7, /*  362 */
128'hfce608e322c505130000951783878713, /*  363 */
128'h9517bf7522c505130000951784078793, /*  364 */
128'he84aec26f022717980821e2505130000, /*  365 */
128'h0104551302904463440184ae892af406, /*  366 */
128'h740270a2952201045513942a90411442, /*  367 */
128'h808261459141694264e21542fff54513, /*  368 */
128'h090900c147836df050ef0068460985ca, /*  369 */
128'h578300f1072300d1478300f107a334f9, /*  370 */
128'hfc26e486e0a26785715dbf55943e00e1, /*  371 */
128'h67a13cf50563842e80678793f44ef84a, /*  372 */
128'h44079a638005079b0af50e636dd78793, /*  373 */
128'h0064091368d050ef4611082884b205e9, /*  374 */
128'h679050ef1ac505130000a517461985ca, /*  375 */
128'h08b7e76332f5896302e0079301744583, /*  376 */
128'h1af58363479104b7e5631cf5826347b1, /*  377 */
128'h00009517478910f58463478502b7e363, /*  378 */
128'h308505130000951702f5836316c50513, /*  379 */
128'h951747a118f582634799a41d7e3030ef, /*  380 */
128'ha4317c9030effef591e3172505130000, /*  381 */
128'h16f58a6347c500b7ed632cf5826347f5, /*  382 */
128'hbf6dfef580e318e505130000951747d9, /*  383 */
128'hfaf596e3029007932af5866302100793, /*  384 */
128'h826306200793b7c91a85051300009517, /*  385 */
128'hef632af582630330079304b7e2632cf5, /*  386 */
128'h95170320079328f5876302f0079300b7, /*  387 */
128'h05c00793b7bdf8f58ae31aa505130000, /*  388 */
128'h1c0505130000951705e0079328f58463, /*  389 */
128'hef6328f5866308400793bf91f6f58de3, /*  390 */
128'h951706c0079326f58b630670079300b7, /*  391 */
128'h08900793b73df4f58ae31d2505130000, /*  392 */
128'h0880079326f589630ff0079326f58863, /*  393 */
128'h5703b73d1dc5051300009517f0f59ce3, /*  394 */
128'h89930000a9970be7d7830000a79701e4, /*  395 */
128'hd7830000a7970204570312f714630b69, /*  396 */
128'h519050ef852285ca461910f71c630a87, /*  397 */
128'h509050ef854a076585930000a5974619, /*  398 */
128'h00f41f23020412230204012301a45783, /*  399 */
128'h02f4102302240513fde4859b01c45783, /*  400 */
128'h00f41e230029d78300f41d230009d783, /*  401 */
128'h578300a10e23812100a10ea3db9ff0ef, /*  402 */
128'hda5fe0ef450185a202f41223862601c1, /*  403 */
128'h00009517bd41fde5051300009517a06d, /*  404 */
128'hbdb5ffa5051300009517b559fec50513, /*  405 */
128'h0254478300f10ea30264470302444783, /*  406 */
128'h0274470300e10ea301c1178300f10e23, /*  407 */
128'h0ea301c119030224470300e10e232781, /*  408 */
128'h56830450071300e10e230234470300e1, /*  409 */
128'h47e2f8d79b230000a79704e79b6301c1, /*  410 */
128'h05130000a517f6e585930000a5974619, /*  411 */
128'h429050efe436f6f72b230000a717f765, /*  412 */
128'hff89061bf4c787930000a79766a24762, /*  413 */
128'h74e2640660a6508060ef450102a40593, /*  414 */
128'h04e69463043007138082616179a27942, /*  415 */
128'h87930000a797f2f72b230000a71747e2, /*  416 */
128'h439cf2a787930000a797c799439cf3a7, /*  417 */
128'h06130000a617f1e686930000a697f7e9, /*  418 */
128'he0ef02a40513f1e585930000a597f1a6, /*  419 */
128'h0000951702e798634d200713b765d47f, /*  420 */
128'hcb6ff0ef852285a654f030eff1450513, /*  421 */
128'h051385ca53b030eff105051300009517, /*  422 */
128'hf6e787e35fe00713bf95ca0ff0ef02a4, /*  423 */
128'h02045703f6f701e317fd67c101e45703, /*  424 */
128'h0868eda585930000a5974611f4f70de3, /*  425 */
128'hb335eea5051300009517b799355050ef, /*  426 */
128'h051300009517b30def05051300009517, /*  427 */
128'h9517b339f145051300009517bb21f065, /*  428 */
128'hf305051300009517b311f2a505130000, /*  429 */
128'h00009517b9c5f4e5051300009517b9ed, /*  430 */
128'hb9f1f725051300009517b1ddf5c50513, /*  431 */
128'h051300009517b9c9f985051300009517, /*  432 */
128'he587d7830000a7970265d703b1e1fa65, /*  433 */
128'h0285d703ecf711e3e50484930000a497, /*  434 */
128'h20000793eaf719e3e427d7830000a797, /*  435 */
128'h85ce461900f59a230165899302058913, /*  436 */
128'he00585930000a59746192a3050ef854a, /*  437 */
128'hdf0585930000a5974619293050ef854e, /*  438 */
128'h50ef852285ca4619281050ef00640513, /*  439 */
128'h578302f4132302a0061301c457832770, /*  440 */
128'hd78300f41e230004d78302f4142301e4, /*  441 */
128'hb36900f416236080079300f41f230024, /*  442 */
128'h46013e9030eff2e505130000951785aa, /*  443 */
128'h30239f0101138307b603300017b7bba5, /*  444 */
128'h759366850034171b00f6741326016081, /*  445 */
128'hb783972a300005379f2d8406871b0387, /*  446 */
128'h849b2581601134235e913c23630c8387, /*  447 */
128'h05938a1d08b8696335b95f200813ffc5, /*  448 */
128'hcfb527818ff1fff7c79300c5963b1010, /*  449 */
128'h0084179bea254390d28787930000a797, /*  450 */
128'h46d496aa068e9ebd8006869b7007f793, /*  451 */
128'hd69b0106d69b0106969b00d100a38726, /*  452 */
128'hc6918005069b0001550300d100230086, /*  453 */
128'h8005859b658502d51a63806686936685, /*  454 */
128'h473b1782270546a1007767139fad377d, /*  455 */
128'h97c285b6300008378f95868a83f502d7, /*  456 */
128'h300017b70405aa1ff0ef862602e64463, /*  457 */
128'h3483852660013403608130838287b823, /*  458 */
128'h0008380300d788338082610101135f81, /*  459 */
128'h0c2007b71101b7e1ff06bc2306a12605, /*  460 */
128'h300014b747812401ec06e42643c0e822, /*  461 */
128'h9517e7990206c163033716938304b703, /*  462 */
128'hc3c00c2007b72ad030efe0a505130000, /*  463 */
128'h4785eb9ff0ef8082610564a2644260e2, /*  464 */
128'ha597461184ae8432ec26f0227179bfc1, /*  465 */
128'ha7970cb050eff4060068c52585930000, /*  466 */
128'h85a6862247b20007a803c0a787930000, /*  467 */
128'hbf4757030000a717bf0888930000a897, /*  468 */
128'h8aeff0efbfc505130000a51704500693, /*  469 */
128'h0085579b8082614564e2740270a28522, /*  470 */
128'h579b0185171b8082914115428d5d0522, /*  471 */
128'h8f750085571bf00686938fd966c10185, /*  472 */
128'h25018d5d8d7900ff07370085151b8fd9, /*  473 */
128'he0a2e486d6c5051300009517715d8082, /*  474 */
128'h1e7030efe85aec56f052f44ef84afc26, /*  475 */
128'h03a30000a71747e1b80788230000a797, /*  476 */
128'h4789b6f70e230000a71703e00793b8f7, /*  477 */
128'h05230000a717578db6f709a30000a717, /*  478 */
128'hb5a585930000a59707f007934611b6f7, /*  479 */
128'h05a30000a717b4e404130000a4170028, /*  480 */
128'h7d8050ef006885a246097e2050efb4f7, /*  481 */
128'hf4fff0efb14989930000a99744814522, /*  482 */
128'h82a10086971bf00606130100063746b2, /*  483 */
128'h9101300017b715028f558f710ff6f693, /*  484 */
128'h8007b70380e7b423934180a7b0231742, /*  485 */
128'hb4234721cbc50513000095178087b703, /*  486 */
128'haa17008007378087b5838007b60382e7, /*  487 */
128'h80e7b4238f4d91c115c2ac2a0a130000, /*  488 */
128'h0000a797abf747030000a717113030ef, /*  489 */
128'h0000a697ab1848030000a817ab87c783, /*  490 */
128'h0000a597a9d646030000a617aa66c683, /*  491 */
128'h0d7030efc6c5051300009517a945c583, /*  492 */
128'h0f230000a71700262b376a8900044783, /*  493 */
128'h07a30000a7173000193700144783a6f7, /*  494 */
128'h4783a6f702230000a71700244783a6f7, /*  495 */
128'ha71700444783a4f70ca30000a7170034, /*  496 */
128'h01a30000a71700544783a4f707230000, /*  497 */
128'ha7230000a797a0079d230000a797a4f7, /*  498 */
128'ha5230000a797a007ab230000a797a007, /*  499 */
128'h0009a783e4a99e07af230000a797a007, /*  500 */
128'h830937835a0b0493f4bfe0ef8522e78d, /*  501 */
128'h03379713830937830207456303379713, /*  502 */
128'h54fd000a2783bfc5c4fff0effc075de3, /*  503 */
128'hf0efbfc1710a84937bf050ef4501dff1, /*  504 */
128'h8087b703300017b7b7d914fdb7e9c35f, /*  505 */
128'h80e7b4238f75e40616fd1141ff8006b7, /*  506 */
128'h95178307b58382e7b823f00707136705, /*  507 */
128'h0513000095177dc030efba2505130000, /*  508 */
128'h880707136709300027f37d0030efbbe5, /*  509 */
128'h95173417907307fe4785300790738fd9, /*  510 */
128'h000f0000100f7ac030efbba505130000, /*  511 */
128'h001547838082014160a2302000730ff0, /*  512 */
128'h00354503002547838f5d07a200054703, /*  513 */
128'h367d57fd808225018d5d05628fd907c2, /*  514 */
128'h0fa3058505050005c703808200f61363, /*  515 */
128'h0023808200f61363367d57fdb7f5fee5, /*  516 */
128'he426ec06e8221101495cbfcd050500b5, /*  517 */
128'h0513478101853903cfa500958413e04a, /*  518 */
128'hc703462d02e0031348a5481586ca0200, /*  519 */
128'h0e5007130107146300a70e6327850006, /*  520 */
128'h040500e4002304050064002301179563, /*  521 */
128'h84ae01c9051300b94783fcc79ee30685, /*  522 */
128'h470301994783c088f59ff0ef00f58423, /*  523 */
128'h0179478300f492238fd90087979b0189, /*  524 */
128'h002300f493238fd90087979b01694703, /*  525 */
128'h611c80826105690264a2644260e20004, /*  526 */
128'h0007468303a0061302000593cf99873e, /*  527 */
128'h00d706630017869300c6986302d5fc63, /*  528 */
128'h577d46050007c683b7dd0705a00d577d, /*  529 */
128'h871b078900b666630ff6f593fd06869b, /*  530 */
128'h850747030000a7178082853ae11c0006, /*  531 */
128'hd683c70d0007c703cb85611cc915bfd5, /*  532 */
128'hc503e406114102e69063008557030067, /*  533 */
128'h4525c391450100157793320060ef0017, /*  534 */
128'hc70301b5c783808245258082014160a2, /*  535 */
128'h1d630007079b8f5d0087979b468d01a5, /*  536 */
128'h8fd50087979b0145c6830155c78300d5, /*  537 */
128'hf02271798082853e27818fd90107979b, /*  538 */
128'h03450993e052e84af4065904e44eec26, /*  539 */
128'h2ae060ef85ce8626468500154503842a, /*  540 */
128'h40f487bb000402234c58505ce1312501, /*  541 */
128'h69a2694264e2740270a2450100e7eb63, /*  542 */
128'hff2a74e34a0500344903808261456a02, /*  543 */
128'h60ef85ce86269cbd4685001445034c5c, /*  544 */
128'hc39900454783b7f94505b7e5397d26c0, /*  545 */
128'hec06e8221101591c80824501f8dff06f, /*  546 */
128'hf0ef892e84aa02b787634401e04ae426, /*  547 */
128'h864a46850014c503ec190005041bfddf, /*  548 */
128'h597d4405c11925011f4060ef03448593, /*  549 */
128'h6105690264a2644260e285220324a823, /*  550 */
128'h022357fde04ae426ec06e82211018082, /*  551 */
128'h4783e52d2501fa3ff0ef842ad91c0005, /*  552 */
128'h979b8fd90087979b4509232447032334, /*  553 */
128'h02f71f63a55707134107d79b776d0107, /*  554 */
128'h010005370005079bd59ff0ef06a40513, /*  555 */
128'h0127f7b31465049300544537fff50913, /*  556 */
128'h2501d33ff0ef0864051300978c634501, /*  557 */
128'h64a2644260e200a035338d0501257533, /*  558 */
128'hf44ef84a715dbfcd450d808261056902, /*  559 */
128'h00053023e85aec56f052fc26e0a2e486, /*  560 */
128'h02054e6347addd9ff0ef8932852e89aa, /*  561 */
128'h638097ba654787930000979700351713, /*  562 */
128'hcb85000447830089b023c01547b184aa, /*  563 */
128'h0563e38d0015779313e060ef00144503, /*  564 */
128'h794274e2640660a647a9c11189110009, /*  565 */
128'hf51380826161853e6b426ae27a0279a2, /*  566 */
128'h7713050060ef00a400a3000400230ff4, /*  567 */
128'h4581f569891100090463fb71478d0015, /*  568 */
128'h0913848a04f51a634785ee1ff0ef8522, /*  569 */
128'hc7894501ffc9478389a623a40a131fa4, /*  570 */
128'h0991094100a9a0232501c5bff0ef854a, /*  571 */
128'h876345090004aa8301048913ff2a14e3, /*  572 */
128'h15e30491c10de9dff0ef852285d6000a, /*  573 */
128'h4785470db7bd00e519634785470dfe99, /*  574 */
128'h04044783bfb947b5c1194a81f6e504e3, /*  575 */
128'hd79b0107979b8fd90087979b03f44703, /*  576 */
128'h478304b44983fef711e3200007134107, /*  577 */
128'h29811a09866300f9e9b30089999b04a4, /*  578 */
128'h01a3fff9079b470501342e2304444903, /*  579 */
128'h012304144b03faf769e30ff7f7930124, /*  580 */
128'hffc900fb77b3fffb079bfa0b03e30164, /*  581 */
128'h00fa6a33008a1a1b0454478304644a03, /*  582 */
128'h448304844503f3c100fa779301441423, /*  583 */
128'h0434478314050e638d450085151b0474, /*  584 */
128'h06bbdfb18fd90087979b250104244703, /*  585 */
128'h873200d7063b9f3d004a571b27810339, /*  586 */
128'hdd8d84ae0364d5bb40c504bbf4c564e3, /*  587 */
128'h73630905165500b93933664119556905, /*  588 */
128'hd458015787bb248900ea873b490d00b6, /*  589 */
128'h15e310e91263470dd05c03542023cc04, /*  590 */
128'h0024949bd408b17ff0ef06040513f00a, /*  591 */
128'h57fdee99e7e324810094d49b1ff4849b, /*  592 */
128'h1963478d00f402a3f8000793c45cc81c, /*  593 */
128'h8fd90087979b064447030654478308f9, /*  594 */
128'h859b06f71b6347054107d79b0107979b, /*  595 */
128'h23344783e13d2501ce5ff0ef8522001a, /*  596 */
128'h979b8fd90087979b000402a323244703, /*  597 */
128'h04f71263a55707134107d79b776d0107, /*  598 */
128'h87932501416157b7a99ff0ef03440513, /*  599 */
128'h77b7a83ff0ef2184051302f517632527, /*  600 */
128'h21c4051300f51c632727879325016141, /*  601 */
128'hc448a63ff0ef22040513c808a6dff0ef, /*  602 */
128'h971793c117c227853da7d78300009797, /*  603 */
128'h2a230124002300f413233cf716230000, /*  604 */
128'h099ba33ff0ef05840513b35147810004, /*  605 */
128'h05e3b545a25ff0ef05440513b5b90005, /*  606 */
128'h0014949b00f915634789d41c9fb5e00a, /*  607 */
128'h9cbd0017d79b8885029787bb478db701, /*  608 */
128'hbffff0ef842ae426ec06e8221101bdc5, /*  609 */
128'h47030cf71063478d00044703ed692501, /*  610 */
128'h20000613034404930af71b6347850054, /*  611 */
128'h22f4092305500793a01ff0ef85264581, /*  612 */
128'h02f40a230520079322f409a3faa00793, /*  613 */
128'h20f40da302f40b230610079302f40aa3, /*  614 */
128'h971b20e40d2302e40ba304100713481c, /*  615 */
128'h0ea320f40e230087571b0107571b0107, /*  616 */
128'h445c20f40fa30187d79b0107d71b20e4, /*  617 */
128'h571b0107571b0107971b501020e40f23, /*  618 */
128'h00a322f4002307200693001445030087, /*  619 */
128'h20d40c230187d79b0107d71b260522e4, /*  620 */
128'h4685d81022f401a322e4012320d40ca3, /*  621 */
128'h460100144503000402a3599050ef85a6, /*  622 */
128'h644260e200a03533250158d050ef4581, /*  623 */
128'hf96337f9ffe5869b4d1c8082610564a2, /*  624 */
128'h80829d2d02d585bb55480025458300f6, /*  625 */
128'he84a71794d180eb7f763478580824501, /*  626 */
128'h470302e5f963892ae44eec26f022f406, /*  627 */
128'h08d70e63468d06d70c63842e46890005, /*  628 */
128'h0094d59b9cad515c0015d49b00f71e63, /*  629 */
128'h740270a257fdc9112501ac7ff0ef9dbd, /*  630 */
128'h0249278380826145853e69a2694264e2, /*  631 */
128'h9dbd94ca1ff4f4930099d59b0014899b, /*  632 */
128'hf993f5792501a93ff0ef0344c483854a, /*  633 */
128'h8fc50087979b880503494783994e1ff9, /*  634 */
128'h515cbf458fe9157d6505bf658391c019, /*  635 */
128'h141bfd592501a63ff0ef9dbd0085d59b, /*  636 */
128'h034945030359478399221fe474130014, /*  637 */
128'h9dbd0075d59b515cb7598fc90087979b, /*  638 */
128'h1fc575130024151bf9352501a39ff0ef, /*  639 */
128'h2501100007b7807ff0ef954a03450513, /*  640 */
128'h4540f82271398082853e4785b76517fd, /*  641 */
128'h00b51523e456e852ec4ef426fc06f04a, /*  642 */
128'h74a2744270e2450900f41c63892a4785, /*  643 */
128'h4f98611c808261216aa26a4269e27902, /*  644 */
128'h9463470d0007c683e02184aefee474e3, /*  645 */
128'h5788fce4f7e30087d703eb15579800e6, /*  646 */
128'h000937839d3d0044d79bd17100892823, /*  647 */
128'h3c2300a92a2394be03478793049688bd, /*  648 */
128'h5a7d843a0027c9838722b75d45010099, /*  649 */
128'hf0ef0134f66385a2000935034a850992, /*  650 */
128'h0c630005041be6fff0efbf752501e59f, /*  651 */
128'hf6f476e34f9c00093783f68afbe30144, /*  652 */
128'h110100a55583b78d4505bfc1413484bb, /*  653 */
128'h0005049bf33ff0ef842aec06e426e822, /*  654 */
128'hec990005049b933ff0ef6008484ce495, /*  655 */
128'h57156c1cf3cff0ef4581020006136c08, /*  656 */
128'h644260e200e782234705601c00e78023, /*  657 */
128'hf822fc06e85271398082610564a28526, /*  658 */
128'h4d1c16ba75634a05e456ec4ef04af426, /*  659 */
128'h89324709000547830af5f063498984aa, /*  660 */
128'h154794630ee78863470d0ae78f63842e, /*  661 */
128'h9dbd009a559b00ba0a3b515c0015da1b, /*  662 */
128'h0a9b8805060996630005099b8b9ff0ef, /*  663 */
128'h014487b3cc191ffa7a130ff97793001a, /*  664 */
128'h0049179b00f7f71316c166850347c783, /*  665 */
128'h478502fa0a239a260ff7f7938fd98ff5, /*  666 */
128'hf0ef9dbd8526009ad59b50dc00f48223, /*  667 */
128'hc40d1ffafa9300099f630005099b86bf, /*  668 */
128'h4785032a8a239aa60ff979130049591b, /*  669 */
128'h69e2790274a2854e744270e200f48223, /*  670 */
128'h0347c783015487b3808261216aa26a42, /*  671 */
128'hb7e90127e9339bc100f979130089591b, /*  672 */
128'h0005099b811ff0ef9dbd0085d59b515c, /*  673 */
128'h0a2394261fe474130014141bfc0992e3, /*  674 */
128'h0aa30089591b0109591b0109191b0324, /*  675 */
128'h9dbd0075d59b515cbf79014482230324, /*  676 */
128'h0024141bf80996e30005099bfd8ff0ef, /*  677 */
128'hda0ff0ef85569aa603440a931fc47413, /*  678 */
128'h0109179b012569338d71f00006372501, /*  679 */
128'h80a30087d79b03240a230107d79b9426, /*  680 */
128'h81a300fa81230189591b0109579b00fa, /*  681 */
128'hfc06ec4ef4267139bf3d4989b745012a, /*  682 */
128'h2903e19d89ae84aae456e852f04af822, /*  683 */
128'h4a05844a04f977634d1c04090a6300c5, /*  684 */
128'h4401052a606304f4636324054c9c5afd, /*  685 */
128'h0887f86347850005041bc43ff0efa821, /*  686 */
128'h74a2744270e28522547d00f41d6357fd, /*  687 */
128'h894e4c9c808261216aa26a4269e27902, /*  688 */
128'h852685a24409bf554905b7d5faf47ee3, /*  689 */
128'h05450863fd5507e3c9012501c05ff0ef, /*  690 */
128'h852685a2167d10000637b76dfb2411e3, /*  691 */
128'hc4c0489c02099063e9052501de9ff0ef, /*  692 */
128'he7930054c783c89c37fdfae783e3577d, /*  693 */
128'hf0ef852685ce8622bf4900f482a30017, /*  694 */
128'hbfad4405f6f50fe34785dd612501dbbf, /*  695 */
128'h17932905f822fc0600a55903f04a7139, /*  696 */
128'h4511eb9993c1e456e852ec4ef4260309, /*  697 */
128'h61216aa26a4269e2790274a2744270e2, /*  698 */
128'h9d63842a8a2e00f97993d7ed495c8082, /*  699 */
128'h00855783e18dc85c61082785480c0009, /*  700 */
128'h012415230996601cfcf775e30009071b, /*  701 */
128'h00254783bf5d4501ec1c97ce03478793, /*  702 */
128'hf0effc0a9fe30157fab337fd00495a9b, /*  703 */
128'hbf4945090097e46347850005049bb27f, /*  704 */
128'he0634d1c6008b761450500f4946357fd, /*  705 */
128'h0005049be81ff0ef480cf60a0ee306f4, /*  706 */
128'hfcf48de357fdfcf48be34785d4bd451d, /*  707 */
128'h200006136008f5792501dd8ff0ef6008, /*  708 */
128'h85a600043a03beeff0ef034505134581, /*  709 */
128'h478360084a0502aa2823aa5ff0ef8552, /*  710 */
128'h6008d91c415787bb591c00faed630025, /*  711 */
128'h01450223b7b9c848a83ff0ef85a6c804, /*  712 */
128'h27855b1c2a856018f1412501d1cff0ef, /*  713 */
128'hec4ef04afc06f426f8227139b7e9db1c, /*  714 */
128'h84aa02f007130005c783e05ae456e852, /*  715 */
128'h04050ce7906305c0071300e78663842e, /*  716 */
128'h0a130ae7fc6347fd000447030004a623, /*  717 */
128'h000447834b2102e0099305c00a9302f0, /*  718 */
128'h0593462d0204b9030d5780630d478263, /*  719 */
128'h0d37926300044783b40ff0ef854a0200, /*  720 */
128'h02e007930b3790630014478301390023, /*  721 */
128'h9763470d1b378e630024478300f900a3, /*  722 */
128'h8526458100f905a302000793943a0947, /*  723 */
128'hf0ef608848cc100510632501adbff0ef, /*  724 */
128'h4783c7e5000747836c98e96d2501cdaf, /*  725 */
128'h0cb78d6300b78593709cef918ba100b7, /*  726 */
128'hfed608e3fff7c683fff7460307850705, /*  727 */
128'hc55c4bdc611cbf75dfdff0ef85264581, /*  728 */
128'h0004bc232501a85ff0ef85264581b791, /*  729 */
128'h6b026aa26a4269e2790274a2744270e2, /*  730 */
128'hf7578be3bf954709bf1d040580826121, /*  731 */
128'hb7ad02400793943a12f6e06302000693, /*  732 */
128'ha0d1486502000313478145a147014681, /*  733 */
128'h954a9101020695130027e793a8dd0505, /*  734 */
128'h00094503c6ed4711a06d268500e50023, /*  735 */
128'h966300d90023469500d515630e500693, /*  736 */
128'h45850037f6930ff7f7930027979b0165, /*  737 */
128'h00d7946346918bb10107671300b69463, /*  738 */
128'hbdfd00e905a394329201160200876713, /*  739 */
128'h4711c50500b7c783709c4511bf654701, /*  740 */
128'ha623cb890207f7930047f713f4e518e3, /*  741 */
128'hfb0dbf154501e80703e30004bc230004, /*  742 */
128'h8bc100b5c7836c8cfbf58b91b73d4515, /*  743 */
128'hbdb9c4c8af2ff0ef0007c503609cdbe5, /*  744 */
128'h45ad46a10ff7f7930027979b05659a63, /*  745 */
128'h000747039722930117020017061b8732, /*  746 */
128'hfd370ae3f95704e3f94706e3f4e374e3, /*  747 */
128'h00054c634185551b0187151b02b6f263, /*  748 */
128'h0008866300054883cf05051300008517, /*  749 */
128'h0ff57513fbf7051bbd6d4519f11710e3, /*  750 */
128'heea866e30ff57513f9f7051beea87ae3, /*  751 */
128'hf0227179bdf90ff777130017e7933701, /*  752 */
128'h0913451184aef406842ae44ee84aec26, /*  753 */
128'hf0ef6008a0b1c90de199484c49bd0e50, /*  754 */
128'hc783c3210007c7036c1ce1292501afaf, /*  755 */
128'h8bfd033780630327026303f7f79300b7, /*  756 */
128'h740270a2450100979a630017b79317e1, /*  757 */
128'hf0ef852245818082614569a2694264e2, /*  758 */
128'hbfe54511b7cd00042a23d9452501c13f, /*  759 */
128'h88fff0ef842ae426ec06e82245811101, /*  760 */
128'ha8cff0ef6008484c0e500493e50d2501, /*  761 */
128'hcb9900978d630007c7836c1ced092501, /*  762 */
128'h13634791dd792501bcdff0ef85224585, /*  763 */
128'h11018082610564a2644260e2451d00f5, /*  764 */
128'h0005049bfa9ff0ef842aec06e426e822, /*  765 */
128'he0850005049ba42ff0ef6008484ce49d, /*  766 */
128'h6c08700c84cff0ef4581020006136c08, /*  767 */
128'h60e200e782234705601c82aff0ef462d, /*  768 */
128'h00b7ed6347858082610564a285266442, /*  769 */
128'h69a2694264e2740270a2450980824509, /*  770 */
128'hf406ec26f02271794d1c808261456a02, /*  771 */
128'h4a05fcf5fde384ae842ae052e44ee84a, /*  772 */
128'hec8ff0ef852285a600f4fa634c1c59fd, /*  773 */
128'hfb490ce3bf754501000914630005091b, /*  774 */
128'h25018afff0ef852285a6460103390763, /*  775 */
128'h00544783c81c278501378a63481cf15d, /*  776 */
128'h4505bf5d0009049b00f402a30017e793, /*  777 */
128'hf42ee432e82efc061028ec2a7139b759, /*  778 */
128'h8c078793000097970405426383eff0ef, /*  779 */
128'h00070023c3196622631800a78733050e, /*  780 */
128'hcb114501e39897aa00070023c3196762, /*  781 */
128'ha0eff0ef0828080c460100f618634785, /*  782 */
128'hf8ca7175bfe5452d8082612170e22501, /*  783 */
128'he42ee8daecd6f0d2f4cefca6e122e506, /*  784 */
128'h8a7984aa89b20005302314050d634925, /*  785 */
128'h140910630005091b9d6ff0ef1028002c, /*  786 */
128'h64062501b6dff0efe4be1028083c65a2, /*  787 */
128'hc3e101f9fa1301c9f7934519e011e119, /*  788 */
128'h2501e75ff0ef102800f516634791c54d, /*  789 */
128'h7aa2cfcd008a77936406e949008a6a13, /*  790 */
128'h00f40ca300f408a30210071304600793, /*  791 */
128'h00040b2300e40823000407a300040723, /*  792 */
128'h00040e23000405a300e40c2300040ba3, /*  793 */
128'h000ac50300040fa300040f2300040ea3, /*  794 */
128'h00040da300040d234785fc9fe0ef85a2, /*  795 */
128'h00fa82230005099b00040aa300040a23, /*  796 */
128'he3fff0ef030aab03855685ce04098b63, /*  797 */
128'hf0ef0135262385da39fd7522e9112501, /*  798 */
128'h8bc500b44783a895892ac90d250183af, /*  799 */
128'hf565a0854921f60981e30049f993e3d9, /*  800 */
128'h84630029f993e72d0107f71300b44783, /*  801 */
128'h020a6a13c399008a7793e3ad8b850009, /*  802 */
128'hd09c01448523f4800309a78385a279a2, /*  803 */
128'h0513c8c8f33fe0ef0009c503000485a3, /*  804 */
128'h0004a623c8880069d783dbbfe0ef01c4, /*  805 */
128'h640a60aa00f494230134b0230004ae23, /*  806 */
128'h61496b466ae67a0679a6794674e6854a, /*  807 */
128'heccef8a27119b7d5491db7e549118082, /*  808 */
128'hf862fc5ee0daf0caf4a6fc86e4d6e8d2, /*  809 */
128'he4328a2e842a0006a023ec6ef06af466, /*  810 */
128'h4783000998630005099be91fe0ef8ab6, /*  811 */
128'h854e744670e60007899bc39d662200b4, /*  812 */
128'h7c427be26b066aa66a4669e6790674a6, /*  813 */
128'h8b8500a44783808261096de27d027ca2, /*  814 */
128'h893e40f907bb445c0104290316078963, /*  815 */
128'h03040b1320000b930006091b00f67463, /*  816 */
128'h120790631ff777934458fa090ce35c7d, /*  817 */
128'h0197fcb337fd0025478300975c9b6008, /*  818 */
128'hec6347854848eb11020c99630ffcfc93, /*  819 */
128'hf0ef4c0cb741498900f405a3478900a7, /*  820 */
128'h00f405a3478501851763b7e52501bd6f, /*  821 */
128'hf0ef856e4c0c00043d83cc08b7a54985, /*  822 */
128'h073b0099579b000c861bd5792501b98f, /*  823 */
128'h9fb1002dc683c4b58d3a0007849b00a6, /*  824 */
128'h863a86a6001dc503419684bb00f6f463, /*  825 */
128'hf79300a44783f94d25010a6050ef85d2, /*  826 */
128'h951b0097fc6341a507bb4c48c3850407, /*  827 */
128'he0ef955285da20000613910115020097, /*  828 */
128'h445c9a3e9381020497930094949bc5ff, /*  829 */
128'ha0239fa5000aa783c45c9fa54099093b, /*  830 */
128'hf79300a4478304e601634c50b70500fa, /*  831 */
128'h50efe43a85da4685001dc503c38d0407, /*  832 */
128'hfbf7f793672200a44783f139250106c0, /*  833 */
128'h85da0017c503863a4685601c00f40523, /*  834 */
128'h049b444c01a42e23f1152501018050ef, /*  835 */
128'h849b0127f46340bb87bb1ff5f5930009, /*  836 */
128'hbd1fe0ef855295a28626030585930007, /*  837 */
128'he0d2e4cee8caf0a27159b59d499dbf9d, /*  838 */
128'he86aec66f062f45ef85aeca6f486fc56, /*  839 */
128'he0ef8ab689328a2e842a0006a023e46e, /*  840 */
128'hc39d00b44783000997630005099bcb5f, /*  841 */
128'h69a6694664e6854e740670a60007899b, /*  842 */
128'h6da26d426ce27c027ba27b427ae26a06, /*  843 */
128'h445c18078f638b8900a4478380826165, /*  844 */
128'h03040b1320000b9304f76c630127873b, /*  845 */
128'h140793631ff777930409046344585c7d, /*  846 */
128'h0197fcb337fd0025478300975c9b6008, /*  847 */
128'hcb914581485cef01040c9a630ffcfc93, /*  848 */
128'hb759498900f405a3478902e798634705, /*  849 */
128'h4818445cf3fd0005079bd86ff0ef4c0c, /*  850 */
128'h00f405230207e79300a4478312f76a63, /*  851 */
128'hbf99498500f405a3478501879763b795, /*  852 */
128'h0407f79300a44783c85ce311cc1c4858, /*  853 */
128'h40ef85da0017c50346854c50601cc38d, /*  854 */
128'h0523fbf7f79300a44783f969250170d0, /*  855 */
128'h250197cff0ef856e4c0c00043d8300f4, /*  856 */
128'h849b00a6863b0099579b000c869bd159, /*  857 */
128'h00f774639fb5002dc703c4b58d320007, /*  858 */
128'h6bf040ef85d286a6001dc503419704bb, /*  859 */
128'h959b0297f26341a587bb4c4cf1512501, /*  860 */
128'he0ef855a95d220000613918115820097, /*  861 */
128'h949b00f40523fbf7f79300a44783a4ff, /*  862 */
128'h4099093b445c9a3e9381020497930094, /*  863 */
128'hbdd100faa0239fa5000aa783c45c9fa5, /*  864 */
128'hc50300e7fa63445c481800c78e634c5c, /*  865 */
128'h2e23fd092501623040ef85da4685001d, /*  866 */
128'h40ab87bb1ff575130009049b444801a4, /*  867 */
128'h85d28626030505130007849b0127f463, /*  868 */
128'h05230407e79300a447839dbfe0ef9522, /*  869 */
128'he0221141bd2d499db5f9c81cbf4100f4, /*  870 */
128'h00a44783e1752501acffe0ef842ae406, /*  871 */
128'h4c50601cc3950407f793cf690207f713, /*  872 */
128'h25015e1040ef030405930017c5034685, /*  873 */
128'h500c00f40523fbf7f79300a44783ed55, /*  874 */
128'h00b7c703741ce15d2501b77fe0ef6008, /*  875 */
128'hd69b0107169b481800e785a302076713, /*  876 */
128'h569b00d78ea300e78e230086d69b0106, /*  877 */
128'h485800e78fa300d78f230187571b0107, /*  878 */
128'h0107169b00e78d2300078ba300078b23, /*  879 */
128'h571b0107171b00e78a2327010107571b, /*  880 */
128'h07130106d69b00e78aa30087571b0107, /*  881 */
128'h8da3046007130086d69b00e78c230210, /*  882 */
128'h4783000789a30007892300e78ca300d7, /*  883 */
128'h0223478500f40523fdf7f793600800a4, /*  884 */
128'h60a24505ebbfe06f014160a2640200f5, /*  885 */
128'hf0ef842ae406e0221141808201416402, /*  886 */
128'he11925019cbfe0ef8522e9012501efff, /*  887 */
128'he42a110180820141640260a200043023, /*  888 */
128'h0000879700054a6395bfe0efec060028, /*  889 */
128'hbfe5452d8082610560e245011ea78623, /*  890 */
128'heca6f486f0a21028002c4601e42a7159, /*  891 */
128'h1028083c65a2ec190005041bb3bfe0ef, /*  892 */
128'he9916586e41d0005041bcd2ff0efe4be, /*  893 */
128'h616564e6740670a68522cbd8575277a2, /*  894 */
128'h0004c50374a2cb998bc100b5c7838082, /*  895 */
128'h4415fcf41ee34791b7c5c8c897bfe0ef, /*  896 */
128'hf4cef8cae122e506e42afca67175bfd9, /*  897 */
128'he0ef1828002c460184ae00050023f0d2, /*  898 */
128'h597d842677e2ecbe081ce5292501acdf, /*  899 */
128'h4501040a12634a16c2be02f009934bdc, /*  900 */
128'h0307071b1347470300008717e50567a2, /*  901 */
128'h0e94186300e780a303a0071300e78023, /*  902 */
128'h60aa00078023078d00e7812302f00713, /*  903 */
128'h4585808261497a0679a6794674e6640a, /*  904 */
128'hf0ef18284581fd452501f89fe0ef1828, /*  905 */
128'he0ef0007c50365c677e2f5552501e6ef, /*  906 */
128'hf9492501f63fe0ef18284581c2aa8cdf, /*  907 */
128'h65c677e2e1052501e48ff0ef18284581, /*  908 */
128'h458101450e6325018a7fe0ef0007c503, /*  909 */
128'h16e367a24711dd612501a9eff0ef1828, /*  910 */
128'h4781f5cfe0ef1828100cb7594509f8e5, /*  911 */
128'heb05fc97470397361094930102079713, /*  912 */
128'h40f405bbfff7871b04e462630037871b, /*  913 */
128'h1a6396b2920166a20206961300e586bb, /*  914 */
128'h2785b7319c3d01368023fff7c7930127, /*  915 */
128'hfc964603962a1088920102071613b7c1, /*  916 */
128'h67220789bddd4545b7e900c68023377d, /*  917 */
128'h24050785000747039736928102041693, /*  918 */
128'hf426f8227139b709fe9465e3fee78fa3, /*  919 */
128'he0ef84ae842ae456e852ec4efc06f04a, /*  920 */
128'hcf8900b44783000917630005091bfb4f, /*  921 */
128'h69e2790274a2854a744270e20007891b, /*  922 */
128'h4783009777634818808261216aa26a42, /*  923 */
128'he4bd00042623445884bae3918b8900a4, /*  924 */
128'he79300a44783c81cfcf778e34818445c, /*  925 */
128'h1ff7f793445c4481bf7d00f405230207, /*  926 */
128'h0304099300a44783fc960ee34c50d3e5, /*  927 */
128'h0017c50385ce4685601cc3850407f793, /*  928 */
128'hfbf7f79300a44783ed51250126b040ef, /*  929 */
128'h85ce0017c50386264685601c00f40523, /*  930 */
128'h47836008bf59cc44ed352501219040ef, /*  931 */
128'hd6bbfff4869b377dc7290097999b0025, /*  932 */
128'h8ff9413007bb02c6ed630337563b0336, /*  933 */
128'hea634a855a7dd1c19c9dc45c27814c0c, /*  934 */
128'h6008d7b51ff4f793c45c9fa5445c0499, /*  935 */
128'hbfb19ca90094d49bcd112501c87fe0ef, /*  936 */
128'h976347850005059b814ff0efe595484c, /*  937 */
128'h976357fdbded490900f405a3478900f5, /*  938 */
128'hcc0cc84cb5ed490500f405a3478500f5, /*  939 */
128'hfddfe0efcb818b89600800a44783b765, /*  940 */
128'h059bc4bfe0efbf6984cee5990005059b, /*  941 */
128'hfae34f9c601cfabafee3fd4588e30005, /*  942 */
128'hc45c013787bb413484bbcc0c445cfaf5, /*  943 */
128'h4601842ac52de42ef822fc067139b7bd, /*  944 */
128'h65a267e2e1152501fe6fe0ef0828002c, /*  945 */
128'he529250197cff0eff01c101ce01c8522, /*  946 */
128'h30234515e7898bc100b5c783cd996c0c, /*  947 */
128'hc448e30fe0ef0007c50367e2a02d0004, /*  948 */
128'he0ef00f414230067d7838522458167e2, /*  949 */
128'h744270e2f971fcf50be347912501cbdf, /*  950 */
128'hb7c1fcf501e34791bfdd452580826121, /*  951 */
128'he1192501dbafe0ef842ae406e0221141, /*  952 */
128'hf022717980820141640260a200043023, /*  953 */
128'h049bd98fe0ef892e842af406e84aec26, /*  954 */
128'hc5ffe0ef8522458100091f63e8890005, /*  955 */
128'h614564e269428526740270a20005049b, /*  956 */
128'h2501b32ff0ef85224581022430238082, /*  957 */
128'he0ef852285ca00042a2302f513634791, /*  958 */
128'h166347912501f8bfe0ef85224581c68f, /*  959 */
128'h7159bf6584aad16dbf7d00042a2300f5, /*  960 */
128'hf486f0a21028002c460184aee42aeca6, /*  961 */
128'h1028083c65a2e00d0005041bedafe0ef, /*  962 */
128'hcf816786e8010005041b872ff0efe4be, /*  963 */
128'h740670a68522c10fe0ef102885a6c489, /*  964 */
128'h8432f0a27159bfcd44198082616564e6, /*  965 */
128'hf486e0d28522002c46018b2ee42af85a, /*  966 */
128'he0efec66f062f45efc56e4cee8caeca6, /*  967 */
128'h01842c836000000a1c6300050a1be7cf, /*  968 */
128'h70a600fb202302f76263ffec871b481c, /*  969 */
128'h7b427ae26a0669a6694664e685527406, /*  970 */
128'h478500044b83808261656ce27c027ba2, /*  971 */
128'h852285ca4a8559fd4481490902fb9f63, /*  972 */
128'he11109550863093508632501a55fe0ef, /*  973 */
128'hc80400544783fef963e329054c1c2485, /*  974 */
128'h504cb74d009b202300f402a30017e793, /*  975 */
128'h9e631afd4c0944814981490110000ab7, /*  976 */
128'he9212501d10fe0ef0015899b85220009, /*  977 */
128'h4783038b9163200009930344091385ce, /*  978 */
128'h2485e3918fd90087979b000947030019, /*  979 */
128'he02e854ab745fc0c94e33cfd39f90909, /*  980 */
128'h2485e1116582015575332501abcfe0ef, /*  981 */
128'h8a2abfbd4a09b7494a05b7c539f10911, /*  982 */
128'he0ef842ae04aec06e426e8221101bfad, /*  983 */
128'h849bcb9100b44783e4910005049bbc4f, /*  984 */
128'h8082610564a269028526644260e20007, /*  985 */
128'h72e348144458cf390027f71300a44783, /*  986 */
128'hef01600800f40523c8180207e793fed7, /*  987 */
128'h05a3c53900042a232501a58ff0ef484c, /*  988 */
128'h0005091b94dfe0ef4c0cbf7d84aa00a4, /*  989 */
128'h100006374c0cb7dd450502f9146357fd, /*  990 */
128'hf0ef85ca6008f9792501b37fe0ef167d, /*  991 */
128'h00e345094785b769449db7e12501a1cf, /*  992 */
128'hf79300a44783fcf96ae34d1c6008fcf9, /*  993 */
128'h05930017c50346854c50601cdba50407, /*  994 */
128'hf79300a44783f55d2501648040ef0304, /*  995 */
128'h002c4605e42a7175b7b100f40523fbf7, /*  996 */
128'h2501ca0fe0eff8cafca6e122e5061008, /*  997 */
128'h2501e3bfe0efe0be1008081c65a2e905, /*  998 */
128'heb890207f79300b7c78345196786e105, /*  999 */
128'h451dcb810014f79300b5c483c59975e2, /* 1000 */
128'h4503790280826149794674e6640a60aa, /* 1001 */
128'hc89d88c1cc0d0005041bad8fe0ef0009, /* 1002 */
128'h00a8100c02800613fc878de301492783, /* 1003 */
128'h2501951fe0efcaa200a8458996cfe0ef, /* 1004 */
128'h4791d94d2501836ff0ef00a84581f161, /* 1005 */
128'he411f15525019f5fe0ef1008faf518e3, /* 1006 */
128'hf0ef85a27502bf612501f20fe0ef7502, /* 1007 */
128'h002c4605e42a7171b769d575250191cf, /* 1008 */
128'hfcd6e152e54ee94aed26f506f1221028, /* 1009 */
128'h041bbd0fe0efe8eaece6f0e2f4def8da, /* 1010 */
128'he0efe4be1028083c65a21c0414630005, /* 1011 */
128'h1af4176347911c0409630005041bd67f, /* 1012 */
128'h18079f630207f79300b7c783441967a6, /* 1013 */
128'h180902630005091bb45fe0ef45817522, /* 1014 */
128'h16f90b63440557fd16f90f6344094785, /* 1015 */
128'h7422160414630005041ba98fe0ef7522, /* 1016 */
128'h03440a13f6efe0ef85220109549b85ca, /* 1017 */
128'h898fe0ef855200050c1b458120000613, /* 1018 */
128'h47c1248188cfe0ef855202000593462d, /* 1019 */
128'h02f40fa30104949b0109199b0ff4fb13, /* 1020 */
128'h02e00b930104d49b021007930109d99b, /* 1021 */
128'h0089d99b046007930ff97a9304f40623, /* 1022 */
128'h03740a230200061304f406a30084d49b, /* 1023 */
128'h053407a305540723040405a304040523, /* 1024 */
128'he0ef0544051385d2049404a305640423, /* 1025 */
128'h57d200074603468d05740aa3772280ef, /* 1026 */
128'h06f40723478100f69363571400d61663, /* 1027 */
128'h979b06f4042327810107d79b0107969b, /* 1028 */
128'hd79b0086d69b0107d79b0106d69b0107, /* 1029 */
128'h4c8500274b8306f404a306d407a30087, /* 1030 */
128'he8350005041bf59fe0ef1028040b9963, /* 1031 */
128'h8c230210071300e785a3752247416786, /* 1032 */
128'h8ca300078ba300078b230460071300e7, /* 1033 */
128'h8aa301678a2301378da301578d2300e7, /* 1034 */
128'h0005041bd5afe0ef00f5022347850097, /* 1035 */
128'h0195022303852823001c0d1b7522a82d, /* 1036 */
128'h458120000613ec090005041b8dcfe0ef, /* 1037 */
128'hb7498c6a0ffbfb93f61fd0ef3bfd8552, /* 1038 */
128'h740a70aa8522f25fe0ef85ca7522441d, /* 1039 */
128'h7c067ba67b467ae66a0a69aa694a64ea, /* 1040 */
128'hf0a27159b7c544218082614d6d466ce6, /* 1041 */
128'hf48610284605002c843284aee42aeca6, /* 1042 */
128'he4be1028083c65a2e13125019cafe0ef, /* 1043 */
128'h00b7c783451967a6e9152501b65fe0ef, /* 1044 */
128'h752200b74783c30d6706e39d0207f793, /* 1045 */
128'h4785008705a38c3d027474138c658cbd, /* 1046 */
128'h64e6740670a62501c9efe0ef00f50223, /* 1047 */
128'h0088002c4605e02ee42a717180826165, /* 1048 */
128'h96630005079b964fe0efed26f122f506, /* 1049 */
128'he0eff0be083cf4be008865a267861207, /* 1050 */
128'h00b7c703778610079a630005079baf7f, /* 1051 */
128'h8e63479165e610071263020777134799, /* 1052 */
128'h02800613e55fd0ef102805ad46550e05, /* 1053 */
128'h47adf05fd0ef850ae49fd0ef10a8008c, /* 1054 */
128'h0005079baadfe0ef10a865820c054d63, /* 1055 */
128'h079bdc5fe0ef10a80ce793634711cbf9, /* 1056 */
128'h00d4851302a10593464d648aefc50005, /* 1057 */
128'h85a30207e793640602814783e0dfd0ef, /* 1058 */
128'hcbbd8bc100b4c78300f40223478500f4, /* 1059 */
128'hd0ef85a60004450306f7086357d64736, /* 1060 */
128'h0005059bcaefe0ef85220005059bf2df, /* 1061 */
128'hefb10005079bfc3fd0ef8522c5a54789, /* 1062 */
128'h57d602f69d630557468302e007936706, /* 1063 */
128'h042327810107d79b06f707230107969b, /* 1064 */
128'hd69b0087d79b0107d79b0107979b06f7, /* 1065 */
128'h06d707a3478506f704a30086d69b0106, /* 1066 */
128'he7910005079be24fe0ef008800f70223, /* 1067 */
128'h64ea740a70aa0005079bb50fe0ef6506, /* 1068 */
128'he42ae8a2711dbfcd47a18082614d853e, /* 1069 */
128'h2501810fe0efec861028002c4605842e, /* 1070 */
128'h25019abfe0efe4be1028083c65a2e929, /* 1071 */
128'heb950207f79300b7c783451967a6e129, /* 1072 */
128'h571b00e78b23752200645703cb856786, /* 1073 */
128'h571b00e78c230044570300e78ba30087, /* 1074 */
128'had6fe0ef00f50223478500e78ca30087, /* 1075 */
128'he0cae4a6711d80826125644660e62501, /* 1076 */
128'hec86e8a208284601002c893284aee42a, /* 1077 */
128'h08284581c4b9e0510005041bf9bfd0ef, /* 1078 */
128'he0ef08284585e5592501ca8fe0efd202, /* 1079 */
128'hca1fd0ef8526462d75c2e93d2501b8ff, /* 1080 */
128'hce89000700230200061346ad00b48713, /* 1081 */
128'hc78397a6938117820007869bfff6879b, /* 1082 */
128'h510c656202090a63fec783e3177d0007, /* 1083 */
128'h0793470d6562e0150005041be69fd0ef, /* 1084 */
128'h87930270079300e68463000546830430, /* 1085 */
128'h60e6852200a92023c29fd0ef953e0347, /* 1086 */
128'h00f51563479180826125690664a66446, /* 1087 */
128'h4605e42a711db7d5842abf5500048023, /* 1088 */
128'h0005041bee3fd0efec86e8a21028002c, /* 1089 */
128'h938102061793460100010c2366a2ec55, /* 1090 */
128'h4581ea2902000593eba10007c78397b6, /* 1091 */
128'h4585e8410005041bbd6fe0efda021028, /* 1092 */
128'h650601814783e1792501abbfe0ef1028, /* 1093 */
128'h021007136786bc7fd0ef082c462dc3dd, /* 1094 */
128'h00078ba300078b230460071300e78c23, /* 1095 */
128'h079bbf45863eb74d2605a06100e78ca3, /* 1096 */
128'h06e3000747039736930102079713fff6, /* 1097 */
128'h48b107f00e9343658e2e4781082cfeb7, /* 1098 */
128'h6c6391411542f9f7051b27850006c703, /* 1099 */
128'h708505130000651793411742370100a3, /* 1100 */
128'h60e68522441900eef863a82100070f1b, /* 1101 */
128'h000548030505bfcdf36d808261256446, /* 1102 */
128'h802300fe06b3b7cdffe81be306080563, /* 1103 */
128'h4785752200f500235795a885078500c6, /* 1104 */
128'h4791b7c10005041b8fefe0ef00f50223, /* 1105 */
128'ha55fe0ef1028dbd50181478302f51b63, /* 1106 */
128'hd0ef4581020006136506f4450005041b, /* 1107 */
128'h47216786ae5fd0ef082c462d6506b07f, /* 1108 */
128'h8023f91780e3b751842abf1900e785a3, /* 1109 */
128'h472993811782f4c7e5e30585068500e5, /* 1110 */
128'h01814703f8d771e30007869b02000613, /* 1111 */
128'h2e0305052e83bf89eaf71de30e500793, /* 1112 */
128'he826ec22110105c52883058523030545, /* 1113 */
128'h887687f2869a8646040502938f2ae44a, /* 1114 */
128'h47338dfd00c6c5b3250f8f9300005f97, /* 1115 */
128'h0fc1008fa403000f2583000fa38300b6, /* 1116 */
128'h883b004f2703ff4fa3839db9007585bb, /* 1117 */
128'h073b0105e8330198581b0078159b0105, /* 1118 */
128'h8e358e6d00f6c6339f3100f805bb0077, /* 1119 */
128'h8e590146561b00c6171b9e39008f2383, /* 1120 */
128'h00b7c6b300d383bb00c5873b008383bb, /* 1121 */
128'h00f6d39b007686bb8ebd00cf24038ef9, /* 1122 */
128'h03bbffcfa4039fa100d3e6b30116969b, /* 1123 */
128'h8f2d9fa1007777338f2d0007061b00d7, /* 1124 */
128'h881b0f418f5d0167171b00a7579b9f3d, /* 1125 */
128'h5597f45f17e300e387bb0003869b0005, /* 1126 */
128'h52971caf8f9300005f97292585930000, /* 1127 */
128'hc73300cf7f3300d7cf33292282930000, /* 1128 */
128'h0f3b0025c4030015c383000faf0301e6, /* 1129 */
128'h4318972a070a93aa038a0005c70300ef, /* 1130 */
128'h010f083b004fa70300ef0f3b942a040a, /* 1131 */
128'h68330003a70301b8581b9e3900581f1b, /* 1132 */
128'h8e3d8e7501e7c6339f3100f80f3b010f, /* 1133 */
128'h9eb90176561b0096139b008fa7039e39, /* 1134 */
128'h46b305919f3500cf03bb00c3e6334018, /* 1135 */
128'h9eb90fc101e6c6b3fff5c4838efd007f, /* 1136 */
128'hd69b9fb900e6941b94aa048affcfa703, /* 1137 */
128'h0083c7339fb900d3843b8ec140980126, /* 1138 */
128'h171b00c7579b9f3d0077473301e77733, /* 1139 */
128'h0004069b0003861b000f081b8f5d0147, /* 1140 */
128'h1a8f0f1300005f17f25599e300e407bb, /* 1141 */
128'ha703010fc40311e38393000053978ffa, /* 1142 */
128'h400000c2c4b3942a040a00d7c2b30003, /* 1143 */
128'h94aa048a0043a4039f21011fc4839f25, /* 1144 */
128'h0048171b012fc4830107083b40809e21, /* 1145 */
128'h073b0083a4039e210107683301c8581b, /* 1146 */
128'h00c2863b9ea194aa00e2c2b3048a00f8, /* 1147 */
128'he6330156561b013fc90300b6129b4080, /* 1148 */
128'hc6b3ffc3a4839c3500c702bb03c100c2, /* 1149 */
128'h0106941b992a9ea1090a0056c6b300e7, /* 1150 */
128'h00d2843b8ec1000924830106d69b9fa5, /* 1151 */
128'h579b9f3d8f219fa5005747330007081b, /* 1152 */
128'h069b0002861b0f918f5d0177171b0097, /* 1153 */
128'h829300005297f5f592e300e407bb0004, /* 1154 */
128'h0002a70300d745b38f5dfff647130962, /* 1155 */
128'h038a020f45839f2d022f4403021f4383, /* 1156 */
128'ha5839f2d942a040a418c95aa058a93aa, /* 1157 */
128'h0003a5839e2d0068171b0107083b0042, /* 1158 */
128'hc6139db100f8073b0107683301a8581b, /* 1159 */
128'h00a6139b0082a5839e2d8e3d8e59fff6, /* 1160 */
128'h00c703bb00c3e633400c9ead0166561b, /* 1161 */
128'h02c10075e5b3fff7c593023f44839ead, /* 1162 */
128'h94aa00f5969b048a9db5ffc2a4038db9, /* 1163 */
128'h081b00b385bb40809fa18dd50115d59b, /* 1164 */
128'h9f3d007747339fa18f4dfff747130007, /* 1165 */
128'h0003861b0f118f5d0157171b00b7579b, /* 1166 */
128'h883b6462f3ef9de300e587bb0005869b, /* 1167 */
128'h282300c8863b00d306bb00fe07bb010e, /* 1168 */
128'h80826105692264c2cd70cd34c97c0505, /* 1169 */
128'he45ee85af44ef84afc26e0a2715d653c, /* 1170 */
128'h89ae84aa97b203f7f413ec56f052e486, /* 1171 */
128'h408b07bb04000b9304000b13e53c8932, /* 1172 */
128'h00090a1b00f974639381178200078a1b, /* 1173 */
128'h86560084853385ce020ada93020a1a93, /* 1174 */
128'h176399d641590933481020ef0144043b, /* 1175 */
128'h640660a6b7c997824401852660bc0174, /* 1176 */
128'h61616ba26b426ae27a0279a2794274e2, /* 1177 */
128'hec26842a03f7f793f0227179653c8082, /* 1178 */
128'h97a2f800071300178513e84af406e44e, /* 1179 */
128'h091b40a9863b449d0400099300e78023, /* 1180 */
128'hf5633c9020ef95224581920116020006, /* 1181 */
128'h450197828522603cfc1c078e643c0124, /* 1182 */
128'h614569a2694264e2740270a2fd24fde3, /* 1183 */
128'h04053423639cd4e78793000077978082, /* 1184 */
128'h0797ed3c639cd467879300007797e93c, /* 1185 */
128'h0505059311018082e13cb6c787930000, /* 1186 */
128'h0000769747013bf020efec06850a4641, /* 1187 */
128'h07b3454119c5859300006597f5468693, /* 1188 */
128'h962e0047d613070506890007c78300e1, /* 1189 */
128'hfec68f230007c78397ae000646038bbd, /* 1190 */
128'h05130000751760e2fca71de3fef68fa3, /* 1191 */
128'he5060808842ae122717580826105f165, /* 1192 */
128'he85ff0ef080885a26622f71ff0efe42e, /* 1193 */
128'h640a60aaf83ff0ef0808f01ff0ef0808, /* 1194 */
128'h469100d70d63711c46a1595880826149, /* 1195 */
128'hac2380824501cf980200071300d71763, /* 1196 */
128'hec06e426e82211018082556dbfe50007, /* 1197 */
128'h0000569702f5026384ae842a200007b7, /* 1198 */
128'h100585930000659708800613e4468693, /* 1199 */
128'h60e2fc240f7030ef1105051300006517, /* 1200 */
128'he4266100e82211018082610564a26442, /* 1201 */
128'h0000569702f4026384ae200007b7ec06, /* 1202 */
128'h0c0585930000659702f00613e1c68693, /* 1203 */
128'h60e2e0040b7030ef0d05051300006517, /* 1204 */
128'he4266100e82211018082610564a26442, /* 1205 */
128'h0000569702f4026384ae200007b7ec06, /* 1206 */
128'h080585930000659703600613dec68693, /* 1207 */
128'h60e2e404077030ef0905051300006517, /* 1208 */
128'he8226104e42611018082610564a26442, /* 1209 */
128'h0000769702f48263842e200007b7ec06, /* 1210 */
128'h040585930000659703e00613c9468693, /* 1211 */
128'h90011402037030ef0505051300006517, /* 1212 */
128'he42611018082610564a2644260e2e880, /* 1213 */
128'h02f48263842e200007b7ec06e8226104, /* 1214 */
128'h0000659704500613c486869300007697, /* 1215 */
128'h7f2030ef00c5051300006517ffc58593, /* 1216 */
128'h8082610564a2644260e2ec8090011402, /* 1217 */
128'h84ae200007b7ec06e4266100e8221101, /* 1218 */
128'h04c00613d34686930000569702f40263, /* 1219 */
128'hfc85051300006517fb85859300006597, /* 1220 */
128'h8082610564a2644260e2f0047ae030ef, /* 1221 */
128'h84ae200007b7ec06e4266100e8221101, /* 1222 */
128'h05300613d04686930000569702f40263, /* 1223 */
128'hf885051300006517f785859300006597, /* 1224 */
128'h8082610564a2644260e2f40476e030ef, /* 1225 */
128'hfc06f04af426f82200053983ec4e7139, /* 1226 */
128'h569702f984638436893284ae200007b7, /* 1227 */
128'h85930000659705a00613cca686930000, /* 1228 */
128'h722030efe43af3e5051300006517f2e5, /* 1229 */
128'h79130029191b8b0589890014159b6722, /* 1230 */
128'h70e288a10125e5b30034949b8dd90049, /* 1231 */
128'h612169e2790274a202b9b8238dc57442, /* 1232 */
128'h85224605468147057100e02211418082, /* 1233 */
128'hf35ff0ef45818522f7dff0efe4064581, /* 1234 */
128'h6008f67ff0ef45814605468547058522, /* 1235 */
128'h808201414501640260a2d97ff0ef4581, /* 1236 */
128'h02053c23460546814705e022e4061141, /* 1237 */
128'h45818522f39ff0ef842a458104053023, /* 1238 */
128'hf0ef46054685470545818522ef1ff0ef, /* 1239 */
128'hd4dff06f0141458160a264026008f23f, /* 1240 */
128'h842e200007b7ec06e8226104e4261101, /* 1241 */
128'h06100613bf4686930000569702f48263, /* 1242 */
128'he585051300006517e485859300006597, /* 1243 */
128'h64a2644260e2fc809041144263e030ef, /* 1244 */
128'h07b7ec06e8226104e426110180826105, /* 1245 */
128'hbc0686930000569702f48263842e2000, /* 1246 */
128'h00006517e04585930000659706800613, /* 1247 */
128'he0a08c7d17fd67855fa030efe1450513, /* 1248 */
128'h6100e82211018082610564a2644260e2, /* 1249 */
128'h569702f4026384ae200007b7ec06e426, /* 1250 */
128'h85930000659706f00613b8a686930000, /* 1251 */
128'he4245b4030efdce5051300006517dbe5, /* 1252 */
128'h3903e04a11018082610564a2644260e2, /* 1253 */
128'h84ae842a200007b7ec06e426e8220005, /* 1254 */
128'h07600613b54686930000569702f90263, /* 1255 */
128'hd885051300006517d785859300006597, /* 1256 */
128'h64a2644260e2c84404993c2356e030ef, /* 1257 */
128'he8caeca67100f0a27159808261056902, /* 1258 */
128'hec66f062f45ef85afc56e0d2e4cef486, /* 1259 */
128'hd01ce03084b2892e0005d783020408a3, /* 1260 */
128'h0e049c636ca020ef00c9051345814611, /* 1261 */
128'h200007b700043983bf5ff0ef45856008, /* 1262 */
128'hf71344810049278316f99a6304043a03, /* 1263 */
128'h3c234c1c4485e391448d8b89c7090017, /* 1264 */
128'h86638b85008a2783000a09638cdd0324, /* 1265 */
128'h852245814605468147050144e4931607, /* 1266 */
128'h00892583be1ff0ef85224581d71ff0ef, /* 1267 */
128'h5583c4fff0efacec0c1300005c178522, /* 1268 */
128'hc81ff0efca4a0a1300006a1785220009, /* 1269 */
128'hcf5ff0ef85224581cbdff0ef852285a6, /* 1270 */
128'h45b7d27ff0ef85224581460546854705, /* 1271 */
128'h85224585e93ff0ef852224058593000f, /* 1272 */
128'he593009899b785220d89b583cd1ff0ef, /* 1273 */
128'h00006a9768198993eb7ff0ef25810015, /* 1274 */
128'h694664e6740670a6efe9485cc64a8a93, /* 1275 */
128'h45016ce27c027ba27b427ae26a0669a6, /* 1276 */
128'h488cdb7ff0efe024852244cc80826165, /* 1277 */
128'h603cee079be38b85449cdf3ff0ef8522, /* 1278 */
128'h4781458163900107e683654100043883, /* 1279 */
128'h89e36e89f005051300ff0e3743114701, /* 1280 */
128'h01e8183b070500371f1b00064803ec06, /* 1281 */
128'hf2e50067036316fd060527810107e7b3, /* 1282 */
128'h0087981b010767330187971b0187d81b, /* 1283 */
128'h8fd98fe9010767330087d79b01c87833, /* 1284 */
128'he31c9746938183751782170200be873b, /* 1285 */
128'h9706869300005697b765470147812585, /* 1286 */
128'h00006517b84585930000659714900613, /* 1287 */
128'hbd6100c4e493bd8537a030efb9450513, /* 1288 */
128'h00005597000b1d633b7d20000bb78b4e, /* 1289 */
128'h6f6000efb84505130000651795458593, /* 1290 */
128'h0f20061386e20179096300043903b711, /* 1291 */
128'h4c81485c0709348333a030ef855685d2, /* 1292 */
128'h0c8937830209370312048e6324818cfd, /* 1293 */
128'h4581cc5cf9200793c7817c1c00f76f63, /* 1294 */
128'hf793b27ff0ef85224581b6fff0ef8522, /* 1295 */
128'h6913ff397913852201442903c3950044, /* 1296 */
128'h05130000651785cad47ff0ef85ca0089, /* 1297 */
128'h01442903c3950084f793680000efb265, /* 1298 */
128'hd1fff0ef85ca00496913ff3979138522, /* 1299 */
128'hf793658000efb26505130000651785ca, /* 1300 */
128'h017c8c630384390300043c83cfb50014, /* 1301 */
128'h855685d209c006138c06869300005697, /* 1302 */
128'h02043c2300492783cba97c1c28e030ef, /* 1303 */
128'h0793018c871308e69f630037f693470d, /* 1304 */
128'h161bff87051363104591480d468100c9, /* 1305 */
128'h8f518361ff87370301068763c3900086, /* 1306 */
128'hcbb5603cfeb690e30791872a2685c398, /* 1307 */
128'h8889c85c9bf9485cc85c0027e793485c, /* 1308 */
128'h569701748c63040439036004cc9d4c85, /* 1309 */
128'h30ef855685d20ca0061385a686930000, /* 1310 */
128'h8b850089278300090963040430232100, /* 1311 */
128'hc85c9bf54c85485cb4dff0ef8522ef8d, /* 1312 */
128'h20ef4505d80c8ee3c47ff0ef8522484c, /* 1313 */
128'h00f92623000cb783dbd98b85bd9560f0, /* 1314 */
128'h648397a667a1bf41b1dff0ef8522b771, /* 1315 */
128'h00878913fa978de394be00093c830109, /* 1316 */
128'h0ca139a020efe43e002c46218566639c, /* 1317 */
128'h04800513717908b041635535b7dd87ca, /* 1318 */
128'h30ef892e84b2e44ef406e84aec26f022, /* 1319 */
128'h05130000451785a2cc1d5551842a1000, /* 1320 */
128'h00006517862285aa89aa785010ef7c65, /* 1321 */
128'h200007b702098b634fe000ef9f450513, /* 1322 */
128'h4789cb990024f793f40401242423e01c, /* 1323 */
128'h614569a2694264e2740270a24501c45c, /* 1324 */
128'h8522b7e5c45c4785d4fd450188858082, /* 1325 */
128'h0537458146098082bff9557d0e8030ef, /* 1326 */
128'h6108953e050e200007b7f73ff06f2000, /* 1327 */
128'h07b7e4066380e0221141711c80822501, /* 1328 */
128'h0613762686930000469702f402632000, /* 1329 */
128'h0513000065178d6585930000659734c0, /* 1330 */
128'h60a2557de3914505703c0cc030ef8e65, /* 1331 */
128'hec064501842ae8221101808201416402, /* 1332 */
128'h468560e26622644285a24d3010efe42e, /* 1333 */
128'hf022f4062000051371797940006f6105, /* 1334 */
128'h651784aa006030efe052e44ee84aec26, /* 1335 */
128'h10ef0001b50310e030ef94a505130000, /* 1336 */
128'h681c206010ef842a491010ef450144b0, /* 1337 */
128'h45833f8000ef638c9305051300006517, /* 1338 */
128'h546c3e8000ef92e505130000651706f4, /* 1339 */
128'h91c115c20085d59b9385051300006517, /* 1340 */
128'h05130000651706c44583583c3d2000ef, /* 1341 */
128'h77130187d61b0107d69b0087d71b92e5, /* 1342 */
128'h3a6000ef26010ff6f6930ff7f7930ff7, /* 1343 */
128'h545c398000ef91e50513000065175c0c, /* 1344 */
128'h859300006597c7898a85859300006597, /* 1345 */
128'h6517378000ef90e50513000065178965, /* 1346 */
128'h00006597744805e030ef91a505130000, /* 1347 */
128'h6617584c19c42783db5fb0efe8c58593, /* 1348 */
128'hbd06061300006617e789872606130000, /* 1349 */
128'h4581852633a000ef8f85051300006517, /* 1350 */
128'h8f8a0a1300006a174481ed5ff0ef8426, /* 1351 */
128'h01f4f793200009138f89899300006997, /* 1352 */
128'h854e0004458330c000ef855285a6e789, /* 1353 */
128'h9fe304052fa000ef819100f5f6132485, /* 1354 */
128'h70a22e8000efe165051300006517fd24, /* 1355 */
128'h8082614545016a0269a2694264e27402, /* 1356 */
128'h40f707b30003b6830083b7830103b703, /* 1357 */
128'hb8230017079300d7fe63938117822785, /* 1358 */
128'h0007802345050103b78300a7002300f3, /* 1359 */
128'h96130103b7830083b703808245018082, /* 1360 */
128'h8e9dfff706930003b7038f9992010205, /* 1361 */
128'h40a786bb87aa9d9dfff7059b00c6f563, /* 1362 */
128'h8082852e0007002300b6e6630103b703, /* 1363 */
128'h002307850007c68300d3b82300170693, /* 1364 */
128'h40a0053be681000556634881bfe900d7, /* 1365 */
128'h0ff6f81304100693c219061006934885, /* 1366 */
128'h751302b6733b0005061b385986ba4e25, /* 1367 */
128'h751302b6563b0305051b046e67630ff3, /* 1368 */
128'h40e685bbfe718532fea68fa306850ff5, /* 1369 */
128'h02d007930008876302f5e96303000513, /* 1370 */
128'h80230015559b40e6853b068500f68023, /* 1371 */
128'h808200b61b63fff5081b86ba25810006, /* 1372 */
128'hb7d92585fea68fa30685bf5d00a8053b, /* 1373 */
128'hc8830007c30397ba9381178240c807bb, /* 1374 */
128'hb7f10685011780230066802326050006, /* 1375 */
128'he8d2eccef4a6f8a2597d011cf0ca7119, /* 1376 */
128'hf02ef42afc3e843684b2e0dafc86e4d6, /* 1377 */
128'h591303000a9306c00a1302500993f82a, /* 1378 */
128'h079bc52d8f1d0004c50377a277420209, /* 1379 */
128'h0135086304d7ff639381178276820017, /* 1380 */
128'h0014c503bfe1e7bff0ef020103930485, /* 1381 */
128'h0004c783035510634781048905450f63, /* 1382 */
128'h00f6f36346a50ff7f793fd07879bcb9d, /* 1383 */
128'h06d50f630640069304890014c5034781, /* 1384 */
128'h0630079304d50f630580069302a6eb63, /* 1385 */
128'h69e6790674a6744670e6f55d08f50963, /* 1386 */
128'hc503808261090007051b6b066aa66a46, /* 1387 */
128'h6c6306e50e6307300713b74d048d0024, /* 1388 */
128'h003800840b13f6e51ee30700071300a7, /* 1389 */
128'h071302e5006307500713a00d46014685, /* 1390 */
128'h003800840b13fa850613f6e510e30780, /* 1391 */
128'h0b13f8b50693a81145c1001636134685, /* 1392 */
128'hf0ef400845a946010016b69300380084, /* 1393 */
128'hddbff0ef0028020103930005059be37f, /* 1394 */
128'hf0ef00840b130201039300044503a809, /* 1395 */
128'h01247433600000840b13b5fd845ad93f, /* 1396 */
128'h8522020103930005059b4db010ef8522, /* 1397 */
128'he0c2fc3ef83aec061034f436715db7f1, /* 1398 */
128'h715d8082616160e2e8dff0efe436e4c6, /* 1399 */
128'hf83aec06100005931014862ef436f032, /* 1400 */
128'h616160e2e69ff0efe436e4c6e0c2fc3e, /* 1401 */
128'h05931234862afe36fa32f62e710d8082, /* 1402 */
128'heec6eac2e6bee2baea22ee0608081000, /* 1403 */
128'h85220f7020ef0808842ae3fff0efe436, /* 1404 */
128'h0087b303679c691c80826135645260f2, /* 1405 */
128'h04b7ee63479d80824501830200030363, /* 1406 */
128'h97ba83f92bc707130000471702059793, /* 1407 */
128'h795c878297bae426e822ec061101439c, /* 1408 */
128'h020497930c5010ef7540f55c08c52483, /* 1409 */
128'h4501e91c64a2644260e202f457b39381, /* 1410 */
128'h05e135f1bfd9617cbfe97d5c80826105, /* 1411 */
128'h8082557d8082557db7e9659c95aa058e, /* 1412 */
128'h00055e63ff5ff0ef842ae406e0221141, /* 1413 */
128'h64028522000307630207b303679c681c, /* 1414 */
128'h80820141640260a245018302014160a2, /* 1415 */
128'h00004797150200a7eb6347ad8082557d, /* 1416 */
128'h0000551780826108953e817524478793, /* 1417 */
128'h83020007b303679c691c80824f450513, /* 1418 */
128'h17824785d23e47d502f1102347a1715d, /* 1419 */
128'he486100c200007930030e83ee42e0785, /* 1420 */
128'h4d148082616160a6fd3ff0efcc3ed402, /* 1421 */
128'h308345018082450100e6fe6340040737, /* 1422 */
128'h80822401011322813483230134032381, /* 1423 */
128'h85a2980101f1041322813823dc010113, /* 1424 */
128'hf95ff0ef1a05348322113c2322913423, /* 1425 */
128'hc70302f71c630a0447830a04c703f579, /* 1426 */
128'h47830c04c70302f716630dd447830dd4, /* 1427 */
128'h1a630e0447830e04c70302f710630c04, /* 1428 */
128'h56f010ef0d4485130d440593461100f7, /* 1429 */
128'h0513842af0227179b761fb600513d551, /* 1430 */
128'h1023858a460185226b8020eff4063e80, /* 1431 */
128'h0513e509842af21ff0efc202c4020001, /* 1432 */
128'h80826145740270a2852269a020ef7d00, /* 1433 */
128'hc23ef406f022478500f1102347857179, /* 1434 */
128'h4ad4008007b745386914c195842ac402, /* 1435 */
128'h06b78f75600006b78ff58ff9f8078793, /* 1436 */
128'hf0ef8522858a4601c43e8fd98f554000, /* 1437 */
128'h80826145740270a2c43c47b2e119ec9f, /* 1438 */
128'h07c55783c23e47d500f1102347b5711d, /* 1439 */
128'h6989fdf949370107979bf852fc4ee0ca, /* 1440 */
128'hc43e842e8aaaec86f456e4a6e8a26a05, /* 1441 */
128'h4601e00a0a13e0098993080909134495, /* 1442 */
128'h1005f79345b2ed0de73ff0ef8556858a, /* 1443 */
128'hc78d0125f7b3054793630135f7b3c789, /* 1444 */
128'hfba00513d4bff0ef3505051300005517, /* 1445 */
128'h61257aa27a4279e2690664a6644660e6, /* 1446 */
128'h57630014079b347dfe04c6e334fd8082, /* 1447 */
128'h49e34501b7555a6020ef3e80051300f0, /* 1448 */
128'h0513d09ff0ef3265051300005517fc80, /* 1449 */
128'h102347c17139e7a919c52783bf7df920, /* 1450 */
128'hf426fc06f822858a460147d5c42e00f1, /* 1451 */
128'h8b891b842783c11dde3ff0efc23e842a, /* 1452 */
128'hc901dcdff0ef8522858a46014495cb91, /* 1453 */
128'h45018082612174a2744270e2f8ed34fd, /* 1454 */
128'he8a2ec86e0cae4a6711d80824501bfd5, /* 1455 */
128'h02c9270347c906d7f66384b6892a4785, /* 1456 */
128'h4755d432cf3108c92783260102f11023, /* 1457 */
128'hca26d23a854a100c47850030cc3ee42e, /* 1458 */
128'h0497f0634785e529842ad75ff0efc83e, /* 1459 */
128'hd402854a100c47f5460102f1102347b1, /* 1460 */
128'h2805051300005517c11dd55ff0efd23e, /* 1461 */
128'h6125690664a6644660e68522c43ff0ef, /* 1462 */
128'h0004841bb74d02f6063bbf6147c58082, /* 1463 */
128'hf04af426f822fc067139b7c54401b7d5, /* 1464 */
128'h84b28a2e4148842ace05e456e852ec4e, /* 1465 */
128'h852200b44583c11d892a482010ef8ab6, /* 1466 */
128'h7a63014485b3681000054d638c5fa0ef, /* 1467 */
128'h4481bd9ff0ef236505130000551700b6, /* 1468 */
128'h89a6f96decdff0ef854a08c92583a089, /* 1469 */
128'h86a2844e0089f3630207e40301093783, /* 1470 */
128'h6783fc851ae3f01ff0ef854a85d68652, /* 1471 */
128'h99e39aa2028784339a22408989b308c9, /* 1472 */
128'h6a4269e274a279028526744270e2fc09, /* 1473 */
128'h47f500f1102347997139808261216aa2, /* 1474 */
128'h0106161b8edd030007b70086969bc23e, /* 1475 */
128'h4601440dc43684aafc06f426f8228ed1, /* 1476 */
128'h85263e800593e919c53ff0ef8526858a, /* 1477 */
128'h347d8082612174a2744270e2d91ff0ef, /* 1478 */
128'h3823bffc07b7db0101134d18bfcdfc79, /* 1479 */
128'h22913c2324813023241134239fb92321, /* 1480 */
128'h04131ce7f56349013ffc073723313423, /* 1481 */
128'h1863892ac09ff0ef84aa85a2980101f1, /* 1482 */
128'h6c2020ef20000513e7991a04b7831e05, /* 1483 */
128'h200006131e0503631a04b5031aa4b023, /* 1484 */
128'h1cf76b6347210c044783123010ef85a2, /* 1485 */
128'h07b753b897ba078adf07071300004717, /* 1486 */
128'h0d44278300e7fd63cc981ff787934004, /* 1487 */
128'h00d773630147d69307a6800707136705, /* 1488 */
128'h8b8506f48f2309b449830a044783f8dc, /* 1489 */
128'h0b344783c7890e244783e7810019f993, /* 1490 */
128'hc7898b890a04478300098a6308f480a3, /* 1491 */
128'h091407130e24478306f48fa309c44783, /* 1492 */
128'h09d405130a844783fcdc07c60c848613, /* 1493 */
128'h979b00074583fff74783e0fc07c64681, /* 1494 */
128'hc39197aeffe745839fad0105959b0087, /* 1495 */
128'h478302f585b30e04458300098c634685, /* 1496 */
128'h14e30621070de21c07ce02b787b30dd4, /* 1497 */
128'h468508d4470308e4478304098f63fca7, /* 1498 */
128'h97ba08c447039fb90087171b0107979b, /* 1499 */
128'h02e787b30dd4478302f707330e044703, /* 1500 */
128'h0187979b08a4470308b44783f8fc07ce, /* 1501 */
128'h9fb90087171b089447039fb90107171b, /* 1502 */
128'hf4fc07a6c319f4fc54d89fb908844703, /* 1503 */
128'he3918bfd09c44783c7898b850a044783, /* 1504 */
128'he0bff0ef852645850af006134685ce81, /* 1505 */
128'h0e0446830af447830af407a34785ed35, /* 1506 */
128'hc79954dc08f4aa2300a6979bc7b98b85, /* 1507 */
128'h0dd44783f8dc07a60d44278300098663, /* 1508 */
128'h0a74478308d4ac2302f686bb00a6969b, /* 1509 */
128'h3483854a240134032481308308f48023, /* 1510 */
128'h80822501011322813983230139032381, /* 1511 */
128'h27058bfd8b7d0057d79b00a7d71b50fc, /* 1512 */
128'hb503892abf4d08f4aa2302f707bb2785, /* 1513 */
128'h5951bf651a04b023524020efd1691a04, /* 1514 */
128'h382322113c23dc010113bf455929bf55, /* 1515 */
128'h02f58863478923213023229134232281, /* 1516 */
128'h34032381308354a9c585468102b7e163, /* 1517 */
128'h24010113228134832201390385262301, /* 1518 */
128'h842e4685fef760e34705ffc5879b8082, /* 1519 */
128'hf57184aad1fff0ef892a45850b900613, /* 1520 */
128'h980101f10413f1e9258199f5ffe4059b, /* 1521 */
128'hf7d50b944783e51998dff0ef854a85a2, /* 1522 */
128'he84aec267179b74d84aab75ddf400493, /* 1523 */
128'hf6930ff5f99308154783f022f406e44e, /* 1524 */
128'h84aa45850b3006138edd892e9be10079, /* 1525 */
128'h1c6300f51e63842a57b5c519cc7ff0ef, /* 1526 */
128'h10ef8526842a875ff0ef852685ca0009, /* 1527 */
128'h694264e2740270a28522013505a315e0, /* 1528 */
128'h382328113c23d60101138082614569a2, /* 1529 */
128'h382327313c2329213023289134232881, /* 1530 */
128'h382325713c2327613023275134232741, /* 1531 */
128'h478923b13c2325a13023259134232581, /* 1532 */
128'h9f3dbff7879bbffc07b74d180ac7e963, /* 1533 */
128'h551784ae8b32892abfe787933ffc07b7, /* 1534 */
128'h779307e9460300e7eb63e3a505130000, /* 1535 */
128'hf96ff0efe5c5051300005517e7b90016, /* 1536 */
128'h348329013403298130838522f8400413, /* 1537 */
128'h3a8327013a0327813983280139032881, /* 1538 */
128'h3c8325013c0325813b8326013b032681, /* 1539 */
128'h80822a01011323813d8324013d032481, /* 1540 */
128'haa83db45e34505130000551709892703, /* 1541 */
128'h0005ac83e79102eaf7bb060a81630045, /* 1542 */
128'hf0efe3a5051300005517cb8902ecf7bb, /* 1543 */
128'h4b8502eadabb02c92783bf415429f24f, /* 1544 */
128'h89d6856200c488138c0a009c9c9be399, /* 1545 */
128'hf33b0017859b000828834e114e854781, /* 1546 */
128'hf0efe32505130000551700030d6302e8, /* 1547 */
128'h02e8d33bb7f14b814a814c81b7c1ee4f, /* 1548 */
128'h0107c78397a6078e0208806300652023, /* 1549 */
128'h0ffbfb9300dbebb300be96bbcb898b85, /* 1550 */
128'h8963fbc596e387ae05110821013309bb, /* 1551 */
128'hf00600e3e1450513000055178a09000b, /* 1552 */
128'hf94ff0ef854a85d2fe0a7a1302f10a13, /* 1553 */
128'h161b09ea478309fa4603ee0519e3842a, /* 1554 */
128'h7a63963e09da47839e3d0087979b0106, /* 1555 */
128'he56ff0efe04505130000551785ce0136, /* 1556 */
128'h89b60017f7130a7a46830084c783b5c1, /* 1557 */
128'h47010016e993c3990fe6f9938b89c719, /* 1558 */
128'h581b4b189726070e0017059b46114505, /* 1559 */
128'h571b00b517bb02080463001878130017, /* 1560 */
128'h4187d79b8b050189999b0187979b0027, /* 1561 */
128'h872e0ff9f99300f9e9b3c70d4189d99b, /* 1562 */
128'hef898b850a6a478302d98263fcc592e3, /* 1563 */
128'hc793b5912cc020efdb85051300005517, /* 1564 */
128'hcb898b8509ba4783bfd100f9f9b3fff7, /* 1565 */
128'hb51d547ddbaff0efde85051300005517, /* 1566 */
128'h06134685e3958b850afa4783e20b02e3, /* 1567 */
128'h07a34785e569a21ff0ef854a45850af0, /* 1568 */
128'h049308f92a2300a7979b0e0a47830afa, /* 1569 */
128'h0ff6f69301acd6bb08c00d934d010880, /* 1570 */
128'hf4932485ed499f1ff0ef854a45858626, /* 1571 */
128'hd6bb08f00d134c81ffb492e32d210ff4, /* 1572 */
128'h9cbff0ef854a458586260ff6f693019a, /* 1573 */
128'h4d61ffa492e32ca10ff4f4932485e935, /* 1574 */
128'h45858656000c26834c818aa609b00d93, /* 1575 */
128'he13999dff0ef854a0ff6f6930196d6bb, /* 1576 */
128'hf493248dffac90e30ffafa932ca12a85, /* 1577 */
128'h458509c0061386defdb498e30c110ff4, /* 1578 */
128'h4783d4fb0de34785ed19975ff0ef854a, /* 1579 */
128'h854a458509b00613468501379b630a7a, /* 1580 */
128'h45850a70061386cebb3d842a957ff0ef, /* 1581 */
128'he0221141b32ddd79842a945ff0ef854a, /* 1582 */
128'h679c681c00055e63810ff0ef842ae406, /* 1583 */
128'h014160a264028522000307630187b303, /* 1584 */
128'hf426713980820141640260a245058302, /* 1585 */
128'h478500f5866384aa4791f04af822fc06, /* 1586 */
128'hd78300f110230370079304f592635529, /* 1587 */
128'h8526858a46010107979b4955842e07c4, /* 1588 */
128'h00f110234799ed19d52ff0efc43ec24a, /* 1589 */
128'h858a4601c43e478900f41f634791c24a, /* 1590 */
128'h6121790274a2744270e2d34ff0ef8526, /* 1591 */
128'h6918ee09b7cdc402fef414e347858082, /* 1592 */
128'hf46385be27814f1887ae00f5f3634f5c, /* 1593 */
128'hc2cff06f02c50823dd0c0007059b00e7, /* 1594 */
128'h070d4b9c711910000737691c80828082, /* 1595 */
128'he0dae4d6e8d2eccef0caf4a6fc86f8a2, /* 1596 */
128'hf11ff0ef842ac17c8fd9f466f862fc5e, /* 1597 */
128'h551702042423eb8d6b9c679c681cc509, /* 1598 */
128'h70e6f8500493bacff0efbfa505130000, /* 1599 */
128'h6b066aa66a4669e674a6790685267446, /* 1600 */
128'hf3e54481541c808261097ca27c427be2, /* 1601 */
128'h02f4082347851af42c23478df93ff0ef, /* 1602 */
128'h10ef7d000513ba2ff0ef852202042c23, /* 1603 */
128'hf94584aa97826b9c679c8522681c3ef0, /* 1604 */
128'h08f422231a04282318042e2308842783, /* 1605 */
128'h852245814601b72ff0ef8522d85c4785, /* 1606 */
128'h8522f14984aacf2ff0ef8522f1dff0ef, /* 1607 */
128'h681c00f1102347a1000505a345d000ef, /* 1608 */
128'h0713e3991aa007138ff94bdc00ff8737, /* 1609 */
128'hf0efc23ec43a8522858a460147d50aa0, /* 1610 */
128'h00f715630aa0079300c14703e911bf8f, /* 1611 */
128'h4a55037009933e900913cc1c800207b7, /* 1612 */
128'h0cb780020c3700ff8bb74b0502900a93, /* 1613 */
128'hc402c252013110238522858a46014000, /* 1614 */
128'h4bdc015110234c18681ce13dbb6ff0ef, /* 1615 */
128'h0197e7b301871563c43e0177f7b3c25a, /* 1616 */
128'h47b2ed1db8eff0ef8522858a4601c43e, /* 1617 */
128'h10ef3e80051306090863397d0007ca63, /* 1618 */
128'h073700e68563800207374c14bf452ff0, /* 1619 */
128'h1e23d45c8b8541e7d79bc43ccc188001, /* 1620 */
128'h1f63f9200793b55d18f40ca347850604, /* 1621 */
128'hc34ff0ef85224581c04ff0ef852202f5, /* 1622 */
128'hbfd118f40c2347850007d663443ced09, /* 1623 */
128'h051300005517d965c1cff0ef85224585, /* 1624 */
128'hb58584aab595fa100493a10ff0efa765, /* 1625 */
128'he352e74eeb4aef26f706f3227161551c, /* 1626 */
128'h4401e6eeeaeaeee6f2e2f6defadafed6, /* 1627 */
128'hc7b1199bc7831cd010ef45018baae3b5, /* 1628 */
128'h04f110234789e7b5180b8ca3198bc783, /* 1629 */
128'habaff0efc482c2be855e008c479d4601, /* 1630 */
128'h4495cf818b851b8ba783120500e3842a, /* 1631 */
128'h100503e3842aaa0ff0ef855e008c4601, /* 1632 */
128'hd99ff0ef855ea031020ba423f4fd34fd, /* 1633 */
128'h69ba695a64fa741a70ba8522d55d842a, /* 1634 */
128'h6db66d566cf67c167bb67b567af66a1a, /* 1635 */
128'h0407c163180b8c23048ba7838082615d, /* 1636 */
128'h0205149313b010ef4501b16ff0ef855e, /* 1637 */
128'h842ab36ff0ef855e45853e8009139081, /* 1638 */
128'h117010ef85260007cc63048ba783f155, /* 1639 */
128'h07b7bfe91a5010ef0640051312a96ee3, /* 1640 */
128'h8b8541e7d79b048ba78300fbac234000, /* 1641 */
128'h0f63450dbf0506fb9e23478502fba623, /* 1642 */
128'h0637a029400406370ea61ee345111aa6, /* 1643 */
128'h8a9d0036d61b00cbac234006061b4001, /* 1644 */
128'h96ce964e068a8a3d4009899300003997, /* 1645 */
128'h06bb018ba88345051086a6830f864603, /* 1646 */
128'h180bae231a0ba8238a0500c7d61b02d6, /* 1647 */
128'h0107d69b08dba22308dba42304cba823, /* 1648 */
128'ha8231408dc63090ba62300d5183b8abd, /* 1649 */
128'h06b70107979b14068e6302cba683090b, /* 1650 */
128'h4721938117828fd98ff50107571b003f, /* 1651 */
128'h0a0bbc23030787b300e797b307090785, /* 1652 */
128'h0c0bbc230c0bb8230c0bb4230c0bb023, /* 1653 */
128'h0107d463200007930afbb8230e0bb023, /* 1654 */
128'h00e7f46320000793090ba70308fba623, /* 1655 */
128'h00e78e63577d04cba783c21508fba823, /* 1656 */
128'h04e11023855e008c46010107979b4711, /* 1657 */
128'hd78304f11023479d902ff0efc282c4be, /* 1658 */
128'hc2ca855e008c0107979b4601495507cb, /* 1659 */
128'haa234785e40516e3842a8e4ff0efc4be, /* 1660 */
128'h842ac9aff0ef855e08fb80a357fd08fb, /* 1661 */
128'h855e00b545830f7000ef855ee2051ae3, /* 1662 */
128'h5a63018ba703e0051fe3842affbfe0ef, /* 1663 */
128'h0370079304fba0232789100007b75407, /* 1664 */
128'h0107979b108c460107cbd78306f11023, /* 1665 */
128'h4905d2caed05880ff0efd4bed2ca855e, /* 1666 */
128'h1023988102091a93033007930bf10493, /* 1667 */
128'h855e108c08104b210a854a11d48206f1, /* 1668 */
128'h16e33a7dc131850ff0efd05aec56e826, /* 1669 */
128'h40030637a7a940020637bb45842afe0a, /* 1670 */
128'h08bba82300b515bb89bd0165d59bbd99, /* 1671 */
128'h01e7569b8ff50027979b16f16685b54d, /* 1672 */
128'h4098b5558b1d938100f7571b17828fd5, /* 1673 */
128'h0087161b0187179b0187569b00ff0537, /* 1674 */
128'hf00706138fd167410087569b8e698fd5, /* 1675 */
128'h0187559b40d804fbaa2327818fd58ef1, /* 1676 */
128'h0087571b8de90087159b8ecd0187169b, /* 1677 */
128'h8b3d0187d71b04ebac238f558f718ecd, /* 1678 */
128'hac238001073720d70263468921270063, /* 1679 */
128'h0737040ba7830007596302d7971300eb, /* 1680 */
128'h800107b7018ba70304fba0238fd92000, /* 1681 */
128'ha903639ce3c78793000057971ef71863, /* 1682 */
128'h3497020d1a13044ba783f0be4d05040b, /* 1683 */
128'h79130ff1079300f9793321a484930000, /* 1684 */
128'h00e797bb478540980a05fe07fc1383f9, /* 1685 */
128'h4a81017d8b3716078563278100f977b3, /* 1686 */
128'h77b340dc0007ac8397d6109c840b0b1b, /* 1687 */
128'h45a1400007b7140781630197f7b300f9, /* 1688 */
128'h05b700fc88634591200007b700fc8d63, /* 1689 */
128'h971ff0ef855e0015b59340bc85b31000, /* 1690 */
128'h00ec8d6347a1400007370e051c638daa, /* 1691 */
128'h8cb3100007b700ec8863479120000737, /* 1692 */
128'hdfdfe0ef855e02fbaa23001cb79340fc, /* 1693 */
128'h47994d850ce79163470d01a78663409c, /* 1694 */
128'h17c12d81810007b7d33e47d50af11023, /* 1695 */
128'h855e110c040007930110d53e00fde7b3, /* 1696 */
128'h010c4783e941e91fe0efc93ee552e162, /* 1697 */
128'h14079a631afba823409c09b794638bbd, /* 1698 */
128'hae2308bba2230017b79317ed088ba583, /* 1699 */
128'hfd930ff10793947ff0ef855e460118fb, /* 1700 */
128'h475507cbd7830af1102303700793fe07, /* 1701 */
128'he03ad33a8cee855e110c0107979b4601, /* 1702 */
128'h0af1102347b56702e915e35fe0efd53e, /* 1703 */
128'h855e110c0110040007134791d502d33a, /* 1704 */
128'h0c63e0dfe0efe03ac93ae552e16ee43e, /* 1705 */
128'h017d85b74785f3ed37fd670267a20e05, /* 1706 */
128'h85934601180bae23096ba2231afba823, /* 1707 */
128'heafa94e347a10a918c9ff0ef855e8405, /* 1708 */
128'h4517e6f49fe3096787930000379704a1, /* 1709 */
128'hb61ddf400413cbdfe0ef552505130000, /* 1710 */
128'hac2380020737b519a007071b80011737, /* 1711 */
128'hbbc580030737de075ee30307971300eb, /* 1712 */
128'h4a159881190201000ab70ff104934905, /* 1713 */
128'h08f110234799020a08633a7d09053ac5, /* 1714 */
128'hc556855e010c040007931030c33e47d5, /* 1715 */
128'h4cdcd0051ce3d61fe0efdc3ef84af426, /* 1716 */
128'h961bf006869366c144dcfbe18b8583a5, /* 1717 */
128'ha70302e796938fd18ff50087d79b0087, /* 1718 */
128'hb35d04fba02300876793da06d9e3040b, /* 1719 */
128'h974e837902079713eaf768e34581472d, /* 1720 */
128'h00ff0537040d859366c1b54511872583, /* 1721 */
128'h971b0187d61b0d91000da783f0068693, /* 1722 */
128'h8f510087d79b8e690087961b8f510187, /* 1723 */
128'h008ca703fdb59ee3fefdae238fd98ff5, /* 1724 */
128'h018ba60300f6f8638bbd00c7579b46a5, /* 1725 */
128'hee8686930000369704d61c63800306b7, /* 1726 */
128'h08fbae230087171b1487a78397b6078a, /* 1727 */
128'h8fd10186d61b8ff917fd67c100cca683, /* 1728 */
128'h0613c305c38d03f7771327810126d71b, /* 1729 */
128'h02f757bb8a8d0106d69b02e6073b3e80, /* 1730 */
128'h1b0ba7830adba2230afba02302d606bb, /* 1731 */
128'ha62320000793c79919cba7831afbaa23, /* 1732 */
128'h00051523484000ef855e08fba82308fb, /* 1733 */
128'hccccd6b7aaaab7b708cba70300050623, /* 1734 */
128'h36b327818ef98ff9ccc68693aaa78793, /* 1735 */
128'h8693f0f0f6b79fb500f037b3068600d0, /* 1736 */
128'hff0106b79fb5068a00d036b38ef90f06, /* 1737 */
128'h76c19fb5068e00d036b38ef9f0068693, /* 1738 */
128'hd11c9fb9071200e037338f7502071613, /* 1739 */
128'h07abd70302c7d7b3ed1092010a8bb783, /* 1740 */
128'h85930000459784aa06fbc603074bd683, /* 1741 */
128'ha803a95fe0effef536230245051338e5, /* 1742 */
128'h571b0088579b06cbc603077bc883070b, /* 1743 */
128'h77130ff878130ff7f7930188569b0108, /* 1744 */
128'h04d4851336c585930000459726810ff7, /* 1745 */
128'h3685859300004597074ba603a5ffe0ef, /* 1746 */
128'h8a3d8abd0146561b0106569b06248513, /* 1747 */
128'h02fba4234785740010ef8526a3ffe0ef, /* 1748 */
128'h400407b704fba0232785100007b7b8d1, /* 1749 */
128'h051300004517e691ecf76ce31a0bb683, /* 1750 */
128'h04fba0230017079b70000737bb952e65, /* 1751 */
128'h0027f6931adba42303f7f6930c46c783, /* 1752 */
128'h04eba0230217071bc68900c7f693ce91, /* 1753 */
128'hc7998b8504eba02301076713040ba703, /* 1754 */
128'h040baa0304fba02300c7e793040ba783, /* 1755 */
128'h00fa7a33855e4601088ba583044ba783, /* 1756 */
128'h3b174a85db4ff0efd984849300003497, /* 1757 */
128'hddcc8c9300003c974c2ddaab0b130000, /* 1758 */
128'h3917cbb5278100fa77b300fa97bb409c, /* 1759 */
128'h409c10000db720000d37d8a909130000, /* 1760 */
128'h40dc04f718630017b79317ed00494703, /* 1761 */
128'h00894683c3a18ff900fa77b300092703, /* 1762 */
128'hdebfe0ef855e0fb6f69345850b700613, /* 1763 */
128'hddbfe0ef855e45850b7006134681c131, /* 1764 */
128'h08fba223180bae231a0ba823088ba783, /* 1765 */
128'hfb9911e30931973fe0ef855e035baa23, /* 1766 */
128'he0ef1ba5051300004517f7649fe304a1, /* 1767 */
128'h89634721400006b700092783bb6d925f, /* 1768 */
128'h0017b71341b787b301a78663471100d7, /* 1769 */
128'hf0ef855e408c933fe0ef855e02ebaa23, /* 1770 */
128'h409ce79d0046f79300892683f941808f, /* 1771 */
128'h0017b79317ed088ba583ef8d1afba823, /* 1772 */
128'hcb0ff0ef855e460118fbae2308bba223, /* 1773 */
128'h06130ff6f693bb91fd319fdfe0ef855e, /* 1774 */
128'h4581b7c9f521d31fe0ef855e45850b70, /* 1775 */
128'h11872583974e837902079713fcfc65e3, /* 1776 */
128'h478d6da000ef06cb851300ec4641bf6d, /* 1777 */
128'h0107979b008c460107cbd78304f11023, /* 1778 */
128'h1b63842a96ffe0efc2be47d5855ec4be, /* 1779 */
128'h9e2304e157830007d663018ba783ec05, /* 1780 */
128'h07cbd783c2be479d04f1102347a506fb, /* 1781 */
128'h93bfe0efc4be855e0107979b008c4601, /* 1782 */
128'ha50345e6475647c646b6ea051163842a, /* 1783 */
128'ha42306eba22306fba02304dbae23018b, /* 1784 */
128'h8a3d01a6d61bf2c51a634000063706bb, /* 1785 */
128'hf0a609634505f0c543638ca602e34509, /* 1786 */
128'hfa100413f0eff06f2006061b40010637, /* 1787 */
128'h557d8082557d80824501c56ce54ff06f, /* 1788 */
128'h9dc7879300005797808218b50d238082, /* 1789 */
128'h5717842ae406e02247851141ef9d439c, /* 1790 */
128'haeefe0ef852212a000ef9cf723230000, /* 1791 */
128'h00ef02c00513fc5ff0ef852200055563, /* 1792 */
128'h808201414501640260a20dc000ef13e0, /* 1793 */
128'h6394631c994707130000571780824501, /* 1794 */
128'h168505130000451785aa114102e79063, /* 1795 */
128'h80820141853e478160a2f60fe0efe406, /* 1796 */
128'h8082853ebfd187b600a604630fc7a603, /* 1797 */
128'h4703c105fbdff0efe42eec0611014148, /* 1798 */
128'h0ff007930815470302b7006365a21035, /* 1799 */
128'h60e25535eb3fe06f610560e200f70c63, /* 1800 */
128'h1101bfcdf8400513bfe5450180826105, /* 1801 */
128'h842acd09f7dff0ef84aee822ec06e426, /* 1802 */
128'h644260e2e0800f840413e501cf0ff0ef, /* 1803 */
128'h879300004797bfd555358082610564a2, /* 1804 */
128'h0f8505138082c3980015071b438877e7, /* 1805 */
128'h11018082438876678793000047978082, /* 1806 */
128'hec06e4266380e8228c87879300005797, /* 1807 */
128'h8082610564a2644260e20094176384be, /* 1808 */
128'hb7d56000a9cff0ef8522c78119a44783, /* 1809 */
128'h00004797e79ce39c8987879300005797, /* 1810 */
128'h8807879300005797e50880827007ae23, /* 1811 */
128'he4a6711d8082e308e518e11ce7886798, /* 1812 */
128'hf852fc4e6080e8a28684849300005497, /* 1813 */
128'he0caec86e06ae466e862ec5ef05af456, /* 1814 */
128'h8a9300004a97056a0a1300004a1789aa, /* 1815 */
128'h8b9300004b9704eb0b1300004b17046a, /* 1816 */
128'h4d295e2c8c9300003c9700050c1b04eb, /* 1817 */
128'h7a4279e2690664a660e6644602941563, /* 1818 */
128'h000045176d026ca26c426be27b027aa2, /* 1819 */
128'hc7914901541cddcfe06f612510c50513, /* 1820 */
128'h0fc42603681c89560007c36389524c1c, /* 1821 */
128'h855e85ca00090663dbefe0ef638c855a, /* 1822 */
128'he0ef856685e200978e63601cdb2fe0ef, /* 1823 */
128'h10ef56a505130000351701a98863da4f, /* 1824 */
128'he04ae426ec06e8221101b77160002860, /* 1825 */
128'h511ccbbd4d5ccfad44014d1cc1414401, /* 1826 */
128'h059384aa892ec7ad639cc7bd651ccbad, /* 1827 */
128'hc57c57fdcd21842a15c010ef45051c00, /* 1828 */
128'h3023e90410f502a347850ef52c234799, /* 1829 */
128'h8793fffff797e65ff0ef040528230325, /* 1830 */
128'h302321a787930000179716f43c2391c7, /* 1831 */
128'h681c18f4342320a787930000179718f4, /* 1832 */
128'hf0ef10f400230247c78385220ea42e23, /* 1833 */
128'h80826105690264a2644260e28522e99f, /* 1834 */
128'h6294611c4b468693000046971180106f, /* 1835 */
128'hd713e11897360017671302d786b36518, /* 1836 */
128'h40f007b300f7553b93ed836d8f3d0127, /* 1837 */
128'h051300004517808225018d5d00f717bb, /* 1838 */
128'hfefff0efe022e4061141fc3ff06f6de5, /* 1839 */
128'h640260a28d410105151bfe9ff0ef842a, /* 1840 */
128'hfdbff0efe022e4061141808201412501, /* 1841 */
128'h8d4115029001fd1ff0ef14020005041b, /* 1842 */
128'hfff5c703058587aa80820141640260a2, /* 1843 */
128'h896387aa962a8082fb75fee78fa30785, /* 1844 */
128'hfb65fee78fa30785fff5c703058500c7, /* 1845 */
128'h0585eb09001786930007c70387aa8082, /* 1846 */
128'h87b68082fb75fee78fa30785fff5c703, /* 1847 */
128'h86930007c70387b68082e21987aab7d5, /* 1848 */
128'h00178713fff5c6830585963efb7d0017, /* 1849 */
128'h000780a300c715638082e291fed70fa3, /* 1850 */
128'hfff5c783000547030585b7cd87ba8082, /* 1851 */
128'h0505e3994187d79b0187979b40f707bb, /* 1852 */
128'ha839478100c59463962e8082853ef37d, /* 1853 */
128'h979b40f707bbfff5c783000547030585, /* 1854 */
128'h8082853eff790505e3994187d79b0187, /* 1855 */
128'hc399808200b79363000547830ff5f593, /* 1856 */
128'h000547830ff5f59380824501bfcd0505, /* 1857 */
128'hc70387aabfcd0505dffd808200b79363, /* 1858 */
128'h1101bfcd0785808240a78533e7010007, /* 1859 */
128'h952265a2fe5ff0efec06842ae42ee822, /* 1860 */
128'h7be3157d00b78663000547830ff5f593, /* 1861 */
128'h87aa95aa80826105644260e24501fe85, /* 1862 */
128'h808240a78533e7010007c70300b78563, /* 1863 */
128'h40c785330007c68387aa862ab7fd0785, /* 1864 */
128'h1be3000748030705fed80fe38082ea99, /* 1865 */
128'hc60387aa86aabfcd872eb7d50785fe08, /* 1866 */
128'h070500c80a638082ea1140d785330007, /* 1867 */
128'h0785bfd5872e8082fe081be300074803, /* 1868 */
128'hfee68fe380824501eb1900054703bff9, /* 1869 */
128'hbfd587aeb7e50505fafd0007c6830785, /* 1870 */
128'h4797e519842a84aeec06e426e8221101, /* 1871 */
128'hf0ef85a68522cc1163804da787930000, /* 1872 */
128'hbf2300004797ef8100044783942af9df, /* 1873 */
128'h8082610564a2644260e2852244014a07, /* 1874 */
128'hc78100054783c519f9fff0ef852285a6, /* 1875 */
128'hbfd948a7b92300004797050500050023, /* 1876 */
128'h8526842ac891e822ec066104e4261101, /* 1877 */
128'h60e2e008050500050023c501f73ff0ef, /* 1878 */
128'h00054783c11d8082610564a285266442, /* 1879 */
128'he3110017c703ce810007c68387aacf99, /* 1880 */
128'h4501b7e5078900d780a300e780238082, /* 1881 */
128'h04c79063963e87aacb9d007577938082, /* 1882 */
128'h00c508b3872aff6d377d8fd507a28082, /* 1883 */
128'h5761003657930106ef6340e88833469d, /* 1884 */
128'hf6934725bfc1963a97aa078e02e78733, /* 1885 */
128'h8fa30785bfe1fef73c230721bfd10ff5, /* 1886 */
128'hcb9d8b9d00a5e7b300b50a63bf6dfeb7, /* 1887 */
128'hff8738030721808202c79e63963e87aa, /* 1888 */
128'h5713ff06e8e340f88833ff07bc2307a1, /* 1889 */
128'h07b3963e95ba070e02f707b357e10036, /* 1890 */
128'hbfe1469d00c508b387aa872ebfc100e5, /* 1891 */
128'h7179bf65fee78fa30785fff5c7030585, /* 1892 */
128'he02ee84af406e432ec26852e842af022, /* 1893 */
128'h64636582892ace1184aa6622dcdff0ef, /* 1894 */
128'hf79ff0ef944a864a8522fff6091300c5, /* 1895 */
128'h614564e269428526740270a200040023, /* 1896 */
128'hf0ef00a5e963842ae406e02211418082, /* 1897 */
128'h06b395b280820141640260a28522f57f, /* 1898 */
128'hc78315fdd7e500e587b340b6073300c5, /* 1899 */
128'h00c51563962ab7fd00f6802316fd0005, /* 1900 */
128'h9f990005c703000547838082853e4781, /* 1901 */
128'h808200c51363962ab7dd05850505fbed, /* 1902 */
128'hf0227179bfc50505feb78de300054783, /* 1903 */
128'hf0ef89aee84af406e44eec26852e842a, /* 1904 */
128'h091bd13ff0ef8522c8890005049bd1ff, /* 1905 */
128'h64e2740270a28522440100995b630005, /* 1906 */
128'h397d852285ce86268082614569a26942, /* 1907 */
128'h0ff5f593962abfe90405d175f8bff0ef, /* 1908 */
128'h00150793000547038082450100c51463, /* 1909 */
128'hef630ff5f59347c1b7ed853efeb70be3, /* 1910 */
128'hc7038082853e4781e60187aa260100c7, /* 1911 */
128'h00757713b7f5367d0785feb71ce30007, /* 1912 */
128'hc80387aa0007069b40e7873b47a1c31d, /* 1913 */
128'h02071793faf5078536fdfcb81ce30007, /* 1914 */
128'h179300b7e733008597938e1d953e9381, /* 1915 */
128'h27018edd00365713020796938fd90107, /* 1916 */
128'hf8b71fe30007c703d24d8a1deb1187aa, /* 1917 */
128'h0a63008785130007b803bfcd367d0785, /* 1918 */
128'hfef51be30785f8b712e30007c70300d8, /* 1919 */
128'h00054703e7a9419cb7f1377d87aabfa5, /* 1920 */
128'h000027970015470308f7116303000793, /* 1921 */
128'hc6898a850006c68300e786b3ee478793, /* 1922 */
128'h04d71b63078006930ff777130207071b, /* 1923 */
128'hc3b10447f7930007c78397ba00254703, /* 1924 */
128'h0005470302f71c6347c14198c19c47c1, /* 1925 */
128'h000027170015478302f7166303000793, /* 1926 */
128'h879bc7098b0500074703973ee9470713, /* 1927 */
128'h050900e79363078007130ff7f7930207, /* 1928 */
128'h842ee8221101bf6d47a9bf7d47a18082, /* 1929 */
128'h468100c16583f63ff0efc632ec06006c, /* 1930 */
128'h0007079b00054703e508081300002817, /* 1931 */
128'h00089863044678930006460300f80633, /* 1932 */
128'h00467893808261058536644260e2ec05, /* 1933 */
128'h02d586b3feb7f4e3fd07879b00088b63, /* 1934 */
128'hf793fe07079bc6098a09b7d196be0505, /* 1935 */
128'hf8227139b7e1e008b7cdfc97879b0ff7, /* 1936 */
128'h84b2842ae42e00063023f04afc06f426, /* 1937 */
128'h74a2744270e25529e90165a2b0dff0ef, /* 1938 */
128'hf0ef8522082c892a862e808261217902, /* 1939 */
128'h8f81cb010007c703fe8782e367e2f5df, /* 1940 */
128'h4501e088fcf718e347a9fd279be30785, /* 1941 */
128'hf06f00e6846302d0071300054683b7e9, /* 1942 */
128'h053360a2f23ff0efe40605051141f2df, /* 1943 */
128'hf0ef842ee406e02211418082014140a0, /* 1944 */
128'h02d704630007c70304b00693601cf0df, /* 1945 */
128'h640260a202d70e630470069300e6ea63, /* 1946 */
128'h06b0069302d7076304d0069380820141, /* 1947 */
128'h9fe3052a069007130017c683fed716e3, /* 1948 */
128'h078d00e69863042007130027c683fce6, /* 1949 */
128'h1101bfd50789bff1052a052ab7e9e01c, /* 1950 */
128'h6583e0fff0efc632ec06006c842ee822, /* 1951 */
128'h00054703cfc8081300002817468100c1, /* 1952 */
128'h044678930006460300f806330007079b, /* 1953 */
128'h808261058536644260e2ec0500089863, /* 1954 */
128'hfeb7f4e3fd07879b00088b6300467893, /* 1955 */
128'h079bc6098a09b7d196be050502d586b3, /* 1956 */
128'hb7e1e008b7cdfc97879b0ff7f793fe07, /* 1957 */
128'h0693601cf87ff0ef842ee406e0221141, /* 1958 */
128'h069300e6ea6302d704630007c70304b0, /* 1959 */
128'h069380820141640260a202d70e630470, /* 1960 */
128'hc683fed716e306b0069302d7076304d0, /* 1961 */
128'h0027c683fce69fe3052a069007130017, /* 1962 */
128'h052ab7e9e01c078d00e6986304200713, /* 1963 */
128'h842ae406e0221141bfd50789bff1052a, /* 1964 */
128'h2797fff5c70300a405b395bff0efe589, /* 1965 */
128'h00074703973efff58513c22787930000, /* 1966 */
128'h157d80820141557d640260a2e7198b11, /* 1967 */
128'h8b1100074703973e00054703fea47ae3, /* 1968 */
128'hf06f014105054581462960a26402f77d, /* 1969 */
128'h812100a107a31141fa5ff06f4581d7df, /* 1970 */
128'h462547818082014100e1550300a10723, /* 1971 */
128'hfd07069b8082853ee3190005470345a9, /* 1972 */
128'h879b9fb902f587bb00d667630ff6f693, /* 1973 */
128'h4563842ee406e0221141bff90505fd07, /* 1974 */
128'h357d02b455bb45a900b7f86347a500a0, /* 1975 */
128'h014160a2640202a4753b4529fe7ff0ef, /* 1976 */
128'h0000471707fe47854e60006f03050513, /* 1977 */
128'h1101808204f73a230000471704f73a23, /* 1978 */
128'h84ae862ee4260464041300004417e822, /* 1979 */
128'h95a660e2600ca2fff0efec06600885aa, /* 1980 */
128'h4797e42611018082610564a26442e00c, /* 1981 */
128'he82200a484930000449701a787930000, /* 1982 */
128'h5f050513000035170004b9036380e04a, /* 1983 */
128'h85a26088b9bfd0ef85a24124043bec06, /* 1984 */
128'h051300003517862286aa608ce77fc0ef, /* 1985 */
128'h25730ff0000f0000100fb81fd0ef5e65, /* 1986 */
128'h000025976902834a64a260e26442f140, /* 1987 */
128'he406e022114183026105250105458593, /* 1988 */
128'h640260a2557d008503638c0fa0ef8432, /* 1989 */
128'h01258413f22271698082450180820141, /* 1990 */
128'hf0ef892eea4aee26f606852289aae64e, /* 1991 */
128'h0505fa2ff0ef852600a404b30505faef, /* 1992 */
128'hee631ff00793fff5071beabff0ef9526, /* 1993 */
128'hf80ff0ef8522f4a7a3230000479704e7, /* 1994 */
128'h9526f72ff0ef376505130000351784aa, /* 1995 */
128'h842af62ff0ef852204a7f2630ff00793, /* 1996 */
128'h00a405b3f54ff0ef3585051300003517, /* 1997 */
128'h741270b2abbfd0ef5385051300003517, /* 1998 */
128'h4717200007938082615569b2695264f2, /* 1999 */
128'h850a458110000613b755eef725230000, /* 2000 */
128'hf0ef850a3145859300003597893ff0ef, /* 2001 */
128'h359700f7096302f0079301294703e1af, /* 2002 */
128'h850a85a2e2aff0ef850a50a585930000, /* 2003 */
128'h858a4390ea47879300004797e22ff0ef, /* 2004 */
128'h17934405a4bfd0ef4f05051300003517, /* 2005 */
128'h00004717e8f7362300004717451101f4, /* 2006 */
128'hc6a7942300004797db5ff0efe8f73623, /* 2007 */
128'h4611c4a79e2300004797da7ff0ef4501, /* 2008 */
128'h4797eb1ff0ef854ec505859300004597, /* 2009 */
128'he426ec06e8221101b799e48797230000, /* 2010 */
128'h84ae450d892a08c7df638432478de04a, /* 2011 */
128'h451708a7956325010004d783d69ff0ef, /* 2012 */
128'h25010024d783d53ff0efe1e555030000, /* 2013 */
128'hdc3ff0ef00448513ffc4059b06a79a63, /* 2014 */
128'h4517bea7952300004797d37ff0ef4511, /* 2015 */
128'h000047974611d23ff0efdee555030000, /* 2016 */
128'hf0ef854abcc5859300004597bca79b23, /* 2017 */
128'hdc45d58300004597256000ef4535e2df, /* 2018 */
128'h4797240000ef02000513d35ff0ef4515, /* 2019 */
128'h0000471727850007d783dae787930000, /* 2020 */
128'h278d439cd947879300004797daf71023, /* 2021 */
128'h937fd0ef3fc50513000035170087cf63, /* 2022 */
128'h60e2d61ff06f6105690264a260e26442, /* 2023 */
128'hf022f406717980826105690264a26442, /* 2024 */
128'h0f230115c78300f10fa347090105c783, /* 2025 */
128'h02e78a63470d00e78e6301e1578300f1, /* 2026 */
128'hd06f61453dc505130000351770a27402, /* 2027 */
128'hd0efe42e3b45051300003517842a8e5f, /* 2028 */
128'hd8dff06f614570a265a2740285228d5f, /* 2029 */
128'h0113ebfff06f614505c170a241907402, /* 2030 */
128'h842a232130232291342322813823dc01, /* 2031 */
128'h22113c230028218006134581893284ae, /* 2032 */
128'he802c44a08282040061385a6e92ff0ef, /* 2033 */
128'h23813083f63ff0ef8522002ced4ff0ef, /* 2034 */
128'h24010113220139032281348323013403, /* 2035 */
128'h45974611cb81caa7d783000047978082, /* 2036 */
128'he40611418082cf5ff06fa92585930000, /* 2037 */
128'ha70300e57763878e1041e703492000ef, /* 2038 */
128'h1007e78310a7a22310e1a02327051001, /* 2039 */
128'h4501808201418d5d91011782150260a2, /* 2040 */
128'hfc1ff0ef84aae426e822ec0611018082, /* 2041 */
128'h150202f407b33e8007933ce000ef842a, /* 2042 */
128'h610564a28d0502a7d533644260e29101, /* 2043 */
128'h00ef842af95ff0efe022e40611418082, /* 2044 */
128'h60a202f407b324078793000f47b73a20, /* 2045 */
128'h1101808202a7d5330141910115026402, /* 2046 */
128'h892af63ff0ef84aae04ae426e822ec06, /* 2047 */
128'h24040413000f443702a48533370000ef, /* 2048 */
128'hfe856ee3f45ff0ef0405944a02855433, /* 2049 */
128'he426110180826105690264a2644260e2, /* 2050 */
128'h68048493842ae04aec06e822009894b7, /* 2051 */
128'hf0ef41240433854a89260084f3638922, /* 2052 */
128'h80826105690264a2644260e2f47dfa1f, /* 2053 */
128'h100007b7808200054503808200b50023, /* 2054 */
128'h4783100007378082020575130147c503, /* 2055 */
128'h07b7808200a70023dfe50207f7930147, /* 2056 */
128'h476d00e78623f8000713000782231000, /* 2057 */
128'h071300e78623470d0007822300e78023, /* 2058 */
128'h808200e788230200071300e78423fc70, /* 2059 */
128'h60a2e50900044503842ae406e0221141, /* 2060 */
128'h2797b7f50405fa5ff0ef808201416402, /* 2061 */
128'h97aa973e811100f57713b7a787930000, /* 2062 */
128'h00f5802300e580a30007c78300074703, /* 2063 */
128'hf0efec068121842a002ce82211018082, /* 2064 */
128'hf0ef00914503f65ff0ef00814503fd1f, /* 2065 */
128'h00814503fb7ff0ef0ff47513002cf5df, /* 2066 */
128'h644260e2f43ff0ef00914503f4bff0ef, /* 2067 */
128'h892af406e84aec26f022717980826105, /* 2068 */
128'hf0ef0ff57513002c0089553b54e14461, /* 2069 */
128'h00914503f13ff0ef346100814503f81f, /* 2070 */
128'h694264e2740270a2fe9410e3f0bff0ef, /* 2071 */
128'h892af406e84aec26f022717980826145, /* 2072 */
128'h0ff57513002c0089553354e103800413, /* 2073 */
128'h4503ed1ff0ef346100814503f3fff0ef, /* 2074 */
128'h64e2740270a2fe9410e3ec9ff0ef0091, /* 2075 */
128'hf13ff0efec06002c1101808261456942, /* 2076 */
128'he9fff0ef00914503ea7ff0ef00814503, /* 2077 */
128'h25730ff0000f0000100f8082610560e2, /* 2078 */
128'h8302037ea9c58593000025974305f140, /* 2079 */
128'h4517e2258593000035974605d9010113, /* 2080 */
128'h3c2326813023261134239fa505130000, /* 2081 */
128'ha0ef2541302325313423252138232491, /* 2082 */
128'hd0ef07a5051300003517c5152501e75f, /* 2083 */
128'h3903258134832601340326813083d64f, /* 2084 */
128'h80822701011324013a03248139832501, /* 2085 */
128'h35974605d3afd0ef0705051300003517, /* 2086 */
128'h44812501e85fa0ef0808082585930000, /* 2087 */
128'h140a0a1300003a1709620bf00913e12d, /* 2088 */
128'ha0ef080895ca66050074918102049593, /* 2089 */
128'h45210004099b00c4d41be5052501fedf, /* 2090 */
128'hdbfff0ef000445039452dc9ff0ef880d, /* 2091 */
128'h54020808f3f99cbd47b2286010ef854e, /* 2092 */
128'h0405051300003517c9192501c96fb0ef, /* 2093 */
128'h35974605bf9101e5051300003517bfb9, /* 2094 */
128'hc5112501dabfa0ef4501d3a585930000, /* 2095 */
128'h86a20bf00493bf1d0305051300003517, /* 2096 */
128'hd0ef032505130000351785a201849613, /* 2097 */
128'h85a2c78fd0ef06e5051300003517c84f, /* 2098 */
128'hc981c62e0005059b962f90ef01849513, /* 2099 */
128'h3517bdddc5afd0ef0685051300003517, /* 2100 */
128'h0023e8dff0efc4cfd0ef83a505130000, /* 2101 */
128'ha001ddbff0efe4062501114190020000, /* 2102 */
128'h471780824501808224050513000f4537, /* 2103 */
128'h869300756513157d631c882707130000, /* 2104 */
128'h8082953e055e10d00513e30895360017, /* 2105 */
128'hf0efe4328532ec06e822110102b50633, /* 2106 */
128'h85229e8ff0ef45816622c509842afd1f, /* 2107 */
128'h000035171141808280826105644260e2, /* 2108 */
128'hc0ef20000537bccfd0efe40600450513, /* 2109 */
128'h45018082450180820141450160a2f89f, /* 2110 */
128'h1141808202f5553347a9b00025738082, /* 2111 */
128'hff0505130000351785aa862e86b28736, /* 2112 */
128'h1141a001d2dff0ef4505b90fd0efe406, /* 2113 */
128'h408007b3f57ff0efe406952e842ae022, /* 2114 */
128'h80824505808201418d7d640260a29522, /* 2115 */
128'hf406ec26f02271798082450580824505, /* 2116 */
128'h64e2740270a20096186300c684bb842e, /* 2117 */
128'hedbfc0efe432852285b2808261454501, /* 2118 */
128'h450980824509bff92605200404136622, /* 2119 */
128'h80824501808280828082808245098082, /* 2120 */
128'he426e822ec061101c2dff06f80824501, /* 2121 */
128'h986300d5043300d584b3003796934781, /* 2122 */
128'h380380826105450164a2644260e200c7, /* 2123 */
128'h000035176090600c02e8036360980004, /* 2124 */
128'h0000351785a28626acefd0eff6450513, /* 2125 */
128'h711dbf5d0785a001abefd0eff7c50513, /* 2126 */
128'hfc4ee8a2f7c5051300003517892ae0ca, /* 2127 */
128'he466e4a6ec86e862ec5ef05af456f852, /* 2128 */
128'hf68a0a1300003a17a8efd0ef44018b2e, /* 2129 */
128'h00003c17fff94993f70b8b9300003b97, /* 2130 */
128'h00040c9ba6afd0ef85524ac1f74c0c13, /* 2131 */
128'h03649863448187caa5efd0ef855e85e6, /* 2132 */
128'h87caa48fd0ef856285e6a50fd0ef8552, /* 2133 */
128'h00003517fd5417e3040502b49b634581, /* 2134 */
128'h008486b3a8894501a2efd0eff9c50513, /* 2135 */
128'he39840e9873300349713c689873e8a85, /* 2136 */
128'h8a856390008586b3bf5d07a104856398, /* 2137 */
128'h02e60d6340e9873300359713c689873e, /* 2138 */
128'h35179e8fd0efefe5051300003517058e, /* 2139 */
128'h644660e6557d9dcfd0eff2a505130000, /* 2140 */
128'h6c426be27b027aa27a4279e2690664a6, /* 2141 */
128'he0d27159bfa507a10585808261256ca2, /* 2142 */
128'hf85ae4ceeca6020005138aaa6a05fc56, /* 2143 */
128'he46ee86aec66e8caf0a2f486f062f45e, /* 2144 */
128'h9c4a0a134981bb1ff0ef44818bb28b2e, /* 2145 */
128'h00fa8db300349793238c0c1300003c17, /* 2146 */
128'hef8505130000351703749b6300fb0cb3, /* 2147 */
128'h7ba26a0669a6694670a67406962fd0ef, /* 2148 */
128'h7b4264e685da86266da26d426ce27c02, /* 2149 */
128'h842ac81fe0efe33ff06f61657ae28556, /* 2150 */
128'hc6ffe0ef892ac75fe0ef8d2ac7bfe0ef, /* 2151 */
128'h00a96533010d1d1b0105151b0344f7b3, /* 2152 */
128'h00acb0238d4191011402150201a46433, /* 2153 */
128'hf7930985b1fff0ef4521ef8100adb023, /* 2154 */
128'hb7ad0485b0fff0ef0007c50397e20039, /* 2155 */
128'hec4ef04af426f822fc06e032e42e7139, /* 2156 */
128'he0ef892ac13fe0ef842ac19fe0ef89aa, /* 2157 */
128'h0109179b0105151bc07fe0ef84aac0df, /* 2158 */
128'h8d5d9101178265a2660215028fc18d45, /* 2159 */
128'h00c79c63974e00e58833003797134781, /* 2160 */
128'h6121863e69e2854e790274a270e27442, /* 2161 */
128'h00083703e3148ea907856314d79ff06f, /* 2162 */
128'hfc06e032e42e7139b7f100e830238f29, /* 2163 */
128'h842aba1fe0ef89aaec4ef04af426f822, /* 2164 */
128'hb8ffe0ef84aab95fe0ef892ab9bfe0ef, /* 2165 */
128'h660215028fc18d450109179b0105151b, /* 2166 */
128'h88330037971347818d5d9101178265a2, /* 2167 */
128'h790274a270e2744200c79c63974e00e5, /* 2168 */
128'h07856314d01ff06f6121863e69e2854e, /* 2169 */
128'hb7f100e830238f0900083703e3148e89, /* 2170 */
128'hec4ef04af426f822fc06e032e42e7139, /* 2171 */
128'he0ef892ab23fe0ef842ab29fe0ef89aa, /* 2172 */
128'h0109179b0105151bb17fe0ef84aab1df, /* 2173 */
128'h8d5d9101178265a2660215028fc18d45, /* 2174 */
128'h00c79c63974e00e58833003797134781, /* 2175 */
128'h6121863e69e2854e790274a270e27442, /* 2176 */
128'h3703e31402a686b307856314c89ff06f, /* 2177 */
128'he42e7139b7e100e8302302a707330008, /* 2178 */
128'he0ef89aaec4ef04af426f822fc06e032, /* 2179 */
128'h84aaaa1fe0ef892aaa7fe0ef842aaadf, /* 2180 */
128'h8fc18d450109179b0105151ba9bfe0ef, /* 2181 */
128'h971347818d5d9101178265a266021502, /* 2182 */
128'h70e2744200c79c63974e00e588330037, /* 2183 */
128'hc0dff06f6121863e69e2854e790274a2, /* 2184 */
128'h3703e31402a6d6b3078563144505e111, /* 2185 */
128'he42e7139b7d100e8302302a757330008, /* 2186 */
128'he0ef89aaec4ef04af426f822fc06e032, /* 2187 */
128'h84aaa21fe0ef892aa27fe0ef842aa2df, /* 2188 */
128'h8fc18d450109179b0105151ba1bfe0ef, /* 2189 */
128'h971347818d5d9101178265a266021502, /* 2190 */
128'h70e2744200c79c63974e00e588330037, /* 2191 */
128'hb8dff06f6121863e69e2854e790274a2, /* 2192 */
128'h30238f4900083703e3148ec907856314, /* 2193 */
128'hf426f822fc06e032e42e7139b7f100e8, /* 2194 */
128'h9affe0ef842a9b5fe0ef89aaec4ef04a, /* 2195 */
128'h0105151b9a3fe0ef84aa9a9fe0ef892a, /* 2196 */
128'h178265a2660215028fc18d450109179b, /* 2197 */
128'h974e00e588330037971347818d5d9101, /* 2198 */
128'h69e2854e790274a270e2744200c79c63, /* 2199 */
128'he3148ee907856314b15ff06f6121863e, /* 2200 */
128'he42e7139b7f100e830238f6900083703, /* 2201 */
128'he0ef89aaec4ef04af426f822fc06e032, /* 2202 */
128'h84aa931fe0ef892a937fe0ef842a93df, /* 2203 */
128'h8fc18cc90109179b0105151b92bfe0ef, /* 2204 */
128'h169347018fc59081178265a266021482, /* 2205 */
128'h70e2744200c71c6396ae00d988330037, /* 2206 */
128'ha9dff06f6121863a69e2854e790274a2, /* 2207 */
128'h7159bfc9070500a83023e28800f70533, /* 2208 */
128'he4cef0a2a5c5051300003517892ae8ca, /* 2209 */
128'hec66eca6f486f062f45ef85afc56e0d2, /* 2210 */
128'h0a1300003a17d6dfc0ef44018b3289ae, /* 2211 */
128'h0c1300003c17a4eb8b9300003b97a46a, /* 2212 */
128'hfff44493d4bfc0ef855204000a93a56c, /* 2213 */
128'h460140900cb3d3dfc0ef8885855e85a2, /* 2214 */
128'h0566186397ce00f905b30036179314fd, /* 2215 */
128'hd17fc0ef856285a2d1ffc0efe4328552, /* 2216 */
128'h2405e12984aaa03ff0ef854a85ce6622, /* 2217 */
128'hcf7fc0efa645051300003517fb541be3, /* 2218 */
128'h7ae26a0669a664e669468526740670a6, /* 2219 */
128'h00167693808261656ce27c027ba27b42, /* 2220 */
128'h54fdbf590605e198e3988726c2918766, /* 2221 */
128'h988505130000351784aaeca67159bfc1, /* 2222 */
128'hf062f45ef85afc56e0d2e4cee8caf0a2, /* 2223 */
128'hc97fc0ef44018ab2892ee86af486ec66, /* 2224 */
128'hc58b0b1300003b179709899300003997, /* 2225 */
128'h968c0c1300003c17c58b8b9300003b97, /* 2226 */
128'hc0ef854e04000a13970c8c9300003c97, /* 2227 */
128'h856285a2000bbd03cba500147793c65f, /* 2228 */
128'h85b300361793fffd45134601c53fc0ef, /* 2229 */
128'hc37fc0efe432854e05561c6397ca00f4, /* 2230 */
128'hf0ef852685ca6622c2ffc0ef856685a2, /* 2231 */
128'h00003517fb441ae32405e5298d2a91bf, /* 2232 */
128'h64e6856a740670a6c0ffc0ef97c50513, /* 2233 */
128'h6ce27c027ba27b427ae26a0669a66946, /* 2234 */
128'h00167693bf49000b3d03808261656d42, /* 2235 */
128'h5d7db7790605e198e398872ac291876a, /* 2236 */
128'h8985051300003517842ae8a2711db7e1, /* 2237 */
128'hec86e862ec5ef05af456f852e0cae4a6, /* 2238 */
128'h00003917babfc0ef4c018ab284aefc4e, /* 2239 */
128'h00003b9788cb0b1300003b1788490913, /* 2240 */
128'h099bb89fc0ef854a10000a13894b8b93, /* 2241 */
128'h1793008c1713b7dfc0ef855a85ce000c, /* 2242 */
128'h17138fd9018c17130187e7b38fd9010c, /* 2243 */
128'h8fd9030c17138fd9028c17138fd9020c, /* 2244 */
128'h00e406b30036171346018fd9038c1713, /* 2245 */
128'h85ceb39fc0efe432854a055617639726, /* 2246 */
128'h81dff0ef852285a66622b31fc0ef855e, /* 2247 */
128'h051300003517f94c19e30c05e91d89aa, /* 2248 */
128'h690664a6854e644660e6b11fc0ef87e5, /* 2249 */
128'h808261256c426be27b027aa27a4279e2, /* 2250 */
128'hf4a67119bff159fdb74d0605e29ce31c, /* 2251 */
128'heccef0caf8a27ae505130000251784aa, /* 2252 */
128'hfc86f06af466f862fc5ee0dae4d6e8d2, /* 2253 */
128'h00002a17abbfc0ef44018b32892eec6e, /* 2254 */
128'h07f00b9379cc8c9300002c97794a0a13, /* 2255 */
128'h0a9379ad0d1300002d1703f00c134985, /* 2256 */
128'ha87fc0ef856685a2a8ffc0ef85520800, /* 2257 */
128'h17934601008995b300e99733408b873b, /* 2258 */
128'he432855205661a6397ca00f486b30036, /* 2259 */
128'h85ca6622a5bfc0ef856a85a2a63fc0ef, /* 2260 */
128'hfb541be32405e1398daaf46ff0ef8526, /* 2261 */
128'h744670e6a3bfc0ef7a85051300002517, /* 2262 */
128'h7be26b066aa66a4669e6790674a6856e, /* 2263 */
128'h008c6663808261096de27d027ca27c42, /* 2264 */
128'h5dfdbfe5e298e398bf610605e28ce38c, /* 2265 */
128'h6c8505130000251784aaf4a67119b7f1, /* 2266 */
128'hf862fc5ee0dae4d6e8d2eccef0caf8a2, /* 2267 */
128'hc0ef44018b32892eec6efc86f06af466, /* 2268 */
128'h8c9300002c976aea0a1300002a179d5f, /* 2269 */
128'h00002d1703f00c13498507f00b936b6c, /* 2270 */
128'h85a29a9fc0ef855208000a936b4d0d13, /* 2271 */
128'h96b300f997b3408b87bb9a1fc0ef8566, /* 2272 */
128'h003617134601fff6c693fff7c7930089, /* 2273 */
128'hc0efe432855205661a63974a00e485b3, /* 2274 */
128'h852685ca662296dfc0ef856a85a2975f, /* 2275 */
128'h2517fb5417e32405e1398daae58ff0ef, /* 2276 */
128'h856e744670e694dfc0ef6ba505130000, /* 2277 */
128'h7c427be26b066aa66a4669e6790674a6, /* 2278 */
128'he314008c6663808261096de27d027ca2, /* 2279 */
128'hb7f15dfdbfe5e19ce31cbf610605e194, /* 2280 */
128'hf8a25da505130000251784aaf4a67119, /* 2281 */
128'hf466f862fc5ee0dae4d6e8d2eccef0ca, /* 2282 */
128'h8e7fc0ef44018a32892eec6efc86f06a, /* 2283 */
128'h5c8c0c1300002c175c09899300002997, /* 2284 */
128'h2c9703f00b9308100b134d0507f00a93, /* 2285 */
128'h856285a28bbfc0ef854e5c2c8c930000, /* 2286 */
128'h00fd17b3408b07bb408a873b8b3fc0ef, /* 2287 */
128'h16b300fd17b30024079b8f5d00ed1733, /* 2288 */
128'h16934601fff7c313fff748938fd5008d, /* 2289 */
128'he432854e05461c6396ca00d485330036, /* 2290 */
128'h85ca662286bfc0ef856685a2873fc0ef, /* 2291 */
128'h080007932405ed298daad56ff0ef8526, /* 2292 */
128'h847fc0ef5b45051300002517f8f41be3, /* 2293 */
128'h6aa66a4669e6790674a6856e744670e6, /* 2294 */
128'h808261096de27d027ca27c427be26b06, /* 2295 */
128'h85be00081363859a008bea6300167813, /* 2296 */
128'h85bafe081be385c6b7610605e10ce28c, /* 2297 */
128'h00002517892af0ca7119bf755dfdbfc5, /* 2298 */
128'hec6ef06af466fc5ee8d2ecce4c450513, /* 2299 */
128'he03289aef862e0dae4d6f4a6f8a2fc86, /* 2300 */
128'h2c974aaa0a1300002a17fd0fc0ef4b81, /* 2301 */
128'h4da14bad0d1300002d174b2c8c930000, /* 2302 */
128'hc0ef85524401003b949b01779c334785, /* 2303 */
128'h4a93f98fc0ef856685da00848b3bfa4f, /* 2304 */
128'h974e00e908330036171367824601fffc, /* 2305 */
128'h856a85daf7afc0efe432855206f61063, /* 2306 */
128'h8b2ac5eff0ef854a85ce6622f72fc0ef, /* 2307 */
128'h040007932b85fbb41be38c562405e931, /* 2308 */
128'hf46fc0ef4b45051300002517fafb90e3, /* 2309 */
128'h6aa66a4669e6790674a6855a744670e6, /* 2310 */
128'h808261096de27d027ca27c427be26b06, /* 2311 */
128'h00b83023e30c85d6e11185e200167513, /* 2312 */
128'hf4cef8cafca67175b7e95b7db7490605, /* 2313 */
128'he8daecd6f0d2698502000513892e84aa, /* 2314 */
128'he032f46ef86ae122e506fc66e0e2e4de, /* 2315 */
128'hd90c0c1300003c174a01904ff0ef4a81, /* 2316 */
128'h8bca8b26784c8c9300002c979c498993, /* 2317 */
128'h04fd956396da003d969367824d214d81, /* 2318 */
128'h0863ed45842aba2ff0ef852685ca866e, /* 2319 */
128'h8522e98fc0ef42e5051300002517020a, /* 2320 */
128'h6b466ae67a0679a6794674e6640a60aa, /* 2321 */
128'h4a05808261497da27d427ce26c066ba6, /* 2322 */
128'he0ef842a9b2fe0efec36b7758ba68b4a, /* 2323 */
128'h67a29a0fe0efe42a9a6fe0efe82a9acf, /* 2324 */
128'h15028c510106161b8d5d0105151b6642, /* 2325 */
128'hcea7b823000037978d4166e291011402, /* 2326 */
128'h00fb86330006c683018786b34781e288, /* 2327 */
128'hf7b3ffa795e300d600230ff6f6930785, /* 2328 */
128'h001a879b82eff0ef4521ef910ba1033d, /* 2329 */
128'h81aff0ef0007c50397e68b8d00078a9b, /* 2330 */
128'hf0d2f4cef8ca7175bfa1547dbf0d0d85, /* 2331 */
128'he8daecd6fca66a050200051389ae892a, /* 2332 */
128'h8cb2f46ee122e506f86afc66e0e2e4de, /* 2333 */
128'hc7848493000034974a81fe5fe0ef4b01, /* 2334 */
128'h8c4e8bca664d0d1300002d179c4a0a13, /* 2335 */
128'h059d956397de00fc06b3003d97934d81, /* 2336 */
128'h8863e579842aa82ff0ef854a85ce866e, /* 2337 */
128'h8522d78fc0ef30e5051300002517020a, /* 2338 */
128'h6b466ae67a0679a6794674e6640a60aa, /* 2339 */
128'h4a85808261497da27d427ce26c066ba6, /* 2340 */
128'h842a890fe0efe836ec3eb7758c4a8bce, /* 2341 */
128'h87efe0efe02a884fe0efe42a88afe0ef, /* 2342 */
128'h8c518d590106161b0105151b67026622, /* 2343 */
128'hbca7bc23000037978d41910114021502, /* 2344 */
128'h902393c117c20004d783e38866c267e2, /* 2345 */
128'hd78300f6912393c117c20024d78300f6, /* 2346 */
128'h17c20064d78300f6922393c117c20044, /* 2347 */
128'he0ef4521ef91034df7b300f6932393c1, /* 2348 */
128'hc50397ea8b8d00078b1b001b079bef9f, /* 2349 */
128'h6505b789547dbf290d85ee5fe0ef0007, /* 2350 */
128'hfca6e122fff586138932f8ca71758082, /* 2351 */
128'h230505130000251785aa962a84ae842a, /* 2352 */
128'hf86afc66e0e2e4dee8daecd6f0d2f4ce, /* 2353 */
128'hd9930044d793c7cfc0efec36e506f46e, /* 2354 */
128'h44854a81e43e99a20034d793e83e0014, /* 2355 */
128'h218b8b9300002b97218b0b1300002b17, /* 2356 */
128'h218c8c9300002c97218c0c1300002c17, /* 2357 */
128'h220d8d9300002d97220d0d1300002d17, /* 2358 */
128'h0000251702997863ad0a0a1300003a17, /* 2359 */
128'h74e68556640a60aac1efc0ef21450513, /* 2360 */
128'h7ce26c066ba66b466ae67a0679a67946, /* 2361 */
128'hbf6fc0ef855a85a6808261497da27d42, /* 2362 */
128'hc0ef8562beafc0ef855e85ca00090663, /* 2363 */
128'hf0ef852265a2bdcfc0ef856a85e6be4f, /* 2364 */
128'h6762010a2783bccfc0ef856eed15920f, /* 2365 */
128'h051300002517c58d000a358302f74963, /* 2366 */
128'h852285ce6642008a3783bb0fc0ef1965, /* 2367 */
128'h4a89b98fc0ef18650513000025179782, /* 2368 */
128'h0485b88fc0efeb65051300002517b7e9, /* 2369 */
128'hf022f40617450513000025177179bfa1, /* 2370 */
128'h251704000593c8bfe0efe44ee84aec26, /* 2371 */
128'h051300002517b5cfc0ef172505130000, /* 2372 */
128'hc0ef1b25051300002517b50fc0ef18e5, /* 2373 */
128'hb36fc0ef4485e665051300002517b44f, /* 2374 */
128'h46054685008495b3497901f499934441, /* 2375 */
128'h70a2ff2417e3e6dff0ef240501358533, /* 2376 */
128'h460580828082614569a2694264e27402, /* 2377 */
128'h45a901f61e1346814881470100c5131b, /* 2378 */
128'h0007802397aa000780234000081387f2, /* 2379 */
128'h97aa387d0007802397aa0007802397aa, /* 2380 */
128'h8e15c020267302b71d632705fe0813e3, /* 2381 */
128'h02a68733411686b33e800513c00026f3, /* 2382 */
128'h02a767b302b345bb02c7473340000593, /* 2383 */
128'ha96fc06f14c505130000251702a74733, /* 2384 */
128'h1141bf51c00028f3c02026f3fac710e3, /* 2385 */
128'h4509f75ff0ef4505f7bff0ef4501e406, /* 2386 */
128'hf63ff0ef4521f69ff0ef4511f6fff0ef, /* 2387 */
128'h400007b791011502bff1f5dff0ef4541, /* 2388 */
128'h07b7808225016388400007b78082e388, /* 2389 */
128'h400007b7808225016b880007b8234000, /* 2390 */
128'h0106161b8d5d0085979b808225017b88, /* 2391 */
128'h4000073747812581f7888d51400007b7, /* 2392 */
128'h8b097a98400006b73e80079300b7ef63, /* 2393 */
128'he60380827388400007b7ffe537fdc319, /* 2394 */
128'h051300002517bfe1f710069127850006, /* 2395 */
128'hf14af526f922fd067131afffe06f1865, /* 2396 */
128'h00002517ab7fe0efe15ae556e952ed4e, /* 2397 */
128'h2917080009b74401addfe0ef0bc50513, /* 2398 */
128'h6390078e013407b344950ba909130000, /* 2399 */
128'hfe9416e399afc0ef0405854a0004059b, /* 2400 */
128'h44990a29091300002917020009b74401, /* 2401 */
128'h051345854601868a0137e7b30204079b, /* 2402 */
128'h2405854a85a2862af43ff0efc03e04b0, /* 2403 */
128'h0b1300002b174901fc941ee3962fc0ef, /* 2404 */
128'h2a1707aa8a9300002a97400004b7216b, /* 2405 */
128'h0007c783016907b3499108aa0a130000, /* 2406 */
128'h8622240125816080608ce09c09058556, /* 2407 */
128'hc0ef25818552688c0004b823922fc0ef, /* 2408 */
128'h4709006457930ff47413fd391be3914f, /* 2409 */
128'h00e78c63470504e78163470d02e78b63, /* 2410 */
128'he0ef85228eafc0ef0505051300002517, /* 2411 */
128'h8d6fc0ef04c5051300002517a001b43f, /* 2412 */
128'hc0ef04a5051300002517b7fdd53ff0ef, /* 2413 */
128'h0485051300002517bff1ec0f80ef8c4f, /* 2414 */
128'h000000000000b7e9e2bff0ef8b2fc0ef, /* 2415 */
128'h08082828282828080808080808080808, /* 2416 */
128'h08080808080808080808080808080808, /* 2417 */
128'h101010101010101010101010101010a0, /* 2418 */
128'h10101010101004040404040404040404, /* 2419 */
128'h01010101010101010141414141414110, /* 2420 */
128'h10101010100101010101010101010101, /* 2421 */
128'h02020202020202020242424242424210, /* 2422 */
128'h08101010100202020202020202020202, /* 2423 */
128'h00000000000000000000000000000000, /* 2424 */
128'h00000000000000000000000000000000, /* 2425 */
128'h101010101010101010101010101010a0, /* 2426 */
128'h10101010101010101010101010101010, /* 2427 */
128'h01010101010101010101010101010101, /* 2428 */
128'h02010101010101011001010101010101, /* 2429 */
128'h02020202020202020202020202020202, /* 2430 */
128'h02020202020202021002020202020202, /* 2431 */
128'hc1bdceee242070dbe8c7b756d76aa478, /* 2432 */
128'hfd469501a83046134787c62af57c0faf, /* 2433 */
128'h895cd7beffff5bb18b44f7af698098d8, /* 2434 */
128'h49b40821a679438efd9871936b901122, /* 2435 */
128'he9b6c7aa265e5a51c040b340f61e2562, /* 2436 */
128'he7d3fbc8d8a1e68102441453d62f105d, /* 2437 */
128'h455a14edf4d50d87c33707d621e1cde6, /* 2438 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /* 2439 */
128'hfde5380c6d9d61228771f681fffa3942, /* 2440 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /* 2441 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /* 2442 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /* 2443 */
128'hfc93a039ab9423a7432aff97f4292244, /* 2444 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /* 2445 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /* 2446 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /* 2447 */
128'h0c07020d08030e09040f0a05000b0601, /* 2448 */
128'h020f0c090603000d0a0704010e0b0805, /* 2449 */
128'h09020b040d060f08010a030c050e0700, /* 2450 */
128'h6c5f7465735f64735f63736972776f6c, /* 2451 */
128'h6e67696c615f64730000000000006465, /* 2452 */
128'h645f6b6c635f64730000000000000000, /* 2453 */
128'h69747465735f64730000000000007669, /* 2454 */
128'h735f646d635f6473000000000000676e, /* 2455 */
128'h74657365725f64730000000074726174, /* 2456 */
128'h6e636b6c625f64730000000000000000, /* 2457 */
128'h69736b6c625f64730000000000000074, /* 2458 */
128'h6f656d69745f6473000000000000657a, /* 2459 */
128'h655f7172695f64730000000000007475, /* 2460 */
128'h5f63736972776f6c000000000000006e, /* 2461 */
128'h00000000646d635f74726174735f6473, /* 2462 */
128'h746e695f746961775f63736972776f6c, /* 2463 */
128'h000000000067616c665f747075727265, /* 2464 */
128'h00007172695f64735f63736972776f6c, /* 2465 */
128'h695f646d635f64735f63736972776f6c, /* 2466 */
128'h5f63736972776f6c0000000000007172, /* 2467 */
128'h007172695f646e655f617461645f6473, /* 2468 */
128'h00000000bffe9a8800000000bffead80, /* 2469 */
128'h004c4b40004c4b400030000020000000, /* 2470 */
128'h6d6d5f6472616f62000000020000ffff, /* 2471 */
128'h00000000bffe4ea60064637465675f63, /* 2472 */
128'h00000000bffe4d1200000000bffe4ab4, /* 2473 */
128'h00000000000000000000000000000000, /* 2474 */
128'hffffbd88ffffbd84ffffbd84ffffbd5e, /* 2475 */
128'hffffbd8cffffbd8cffffbd8cffffbd8c, /* 2476 */
128'h00000000bffeb0a800000000bffeb098, /* 2477 */
128'h00000000bffeb0d000000000bffeb0b8, /* 2478 */
128'h00000000bffeb10000000000bffeb0e8, /* 2479 */
128'h00000000bffeb13000000000bffeb118, /* 2480 */
128'h00000000bffeb16000000000bffeb148, /* 2481 */
128'h00000000bffeb19000000000bffeb178, /* 2482 */
128'h40040300400402004004010040040000, /* 2483 */
128'h40050000400405004004040140040400, /* 2484 */
128'h30000000000000030000000040050100, /* 2485 */
128'h60000000000000053000000000000001, /* 2486 */
128'h70000000000000027000000000000004, /* 2487 */
128'h00000001400000007000000000000000, /* 2488 */
128'h00000005000000012000000000000006, /* 2489 */
128'h20000000000000020000000040000000, /* 2490 */
128'h00000000100000000000000100000000, /* 2491 */
128'h1e19140f0d0c0a000000000000000000, /* 2492 */
128'h000186a00000271050463c37322d2823, /* 2493 */
128'h017d7840017d784000989680000f4240, /* 2494 */
128'h031975000319750002faf080018cba80, /* 2495 */
128'h02faf08005f5e10002faf080017d7840, /* 2496 */
128'h00000020000000000bebc2000c65d400, /* 2497 */
128'h00000200000001000000008000000040, /* 2498 */
128'h00002000000010000000080000000400, /* 2499 */
128'h0000c000000080000000600000004000, /* 2500 */
128'h37363534333231300002000000010000, /* 2501 */
128'h2043534952776f4c4645444342413938, /* 2502 */
128'h746f6f622d7520646573696d696e696d, /* 2503 */
128'h00000000647261432d445320726f6620, /* 2504 */
128'he00600003800000039080000edfe0dd0, /* 2505 */
128'h00000000100000001100000028000000, /* 2506 */
128'h0000000000000000a806000059010000, /* 2507 */
128'h00000000010000000000000000000000, /* 2508 */
128'h02000000000000000400000003000000, /* 2509 */
128'h020000000f0000000400000003000000, /* 2510 */
128'h2c6874651b0000001400000003000000, /* 2511 */
128'h007665642d657261622d656e61697261, /* 2512 */
128'h2c687465260000001000000003000000, /* 2513 */
128'h0100000000657261622d656e61697261, /* 2514 */
128'h1a0000000300000000006e65736f6863, /* 2515 */
128'h303140747261752f636f732f2c000000, /* 2516 */
128'h0000003030323531313a303030303030, /* 2517 */
128'h00000000737570630100000002000000, /* 2518 */
128'h01000000000000000400000003000000, /* 2519 */
128'h000000000f0000000400000003000000, /* 2520 */
128'h40787d01380000000400000003000000, /* 2521 */
128'h03000000000000304075706301000000, /* 2522 */
128'h0300000080f0fa024b00000004000000, /* 2523 */
128'h03000000007570635b00000004000000, /* 2524 */
128'h03000000000000006700000004000000, /* 2525 */
128'h0000000079616b6f6b00000005000000, /* 2526 */
128'h7a6874651b0000001300000003000000, /* 2527 */
128'h0000766373697200656e61697261202c, /* 2528 */
128'h34367672720000000b00000003000000, /* 2529 */
128'h0b000000030000000000636466616d69, /* 2530 */
128'h0000393376732c76637369727c000000, /* 2531 */
128'h01000000850000000000000003000000, /* 2532 */
128'h6f72746e6f632d747075727265746e69, /* 2533 */
128'h04000000030000000000000072656c6c, /* 2534 */
128'h0000000003000000010000008f000000, /* 2535 */
128'h1b0000000f00000003000000a0000000, /* 2536 */
128'h000063746e692d7570632c7663736972, /* 2537 */
128'h01000000b50000000400000003000000, /* 2538 */
128'h01000000bb0000000400000003000000, /* 2539 */
128'h01000000020000000200000002000000, /* 2540 */
128'h0030303030303030384079726f6d656d, /* 2541 */
128'h6f6d656d5b0000000700000003000000, /* 2542 */
128'h67000000100000000300000000007972, /* 2543 */
128'h00000040000000000000008000000000, /* 2544 */
128'h0300000000636f730100000002000000, /* 2545 */
128'h03000000020000000000000004000000, /* 2546 */
128'h03000000020000000f00000004000000, /* 2547 */
128'h616972612c6874651b0000001f000000, /* 2548 */
128'h706d697300636f732d657261622d656e, /* 2549 */
128'h000000000300000000007375622d656c, /* 2550 */
128'h303240746e696c6301000000c3000000, /* 2551 */
128'h0d000000030000000000003030303030, /* 2552 */
128'h30746e696c632c76637369721b000000, /* 2553 */
128'hca000000100000000300000000000000, /* 2554 */
128'h07000000010000000300000001000000, /* 2555 */
128'h00000000670000001000000003000000, /* 2556 */
128'h0300000000000c000000000000000002, /* 2557 */
128'h006c6f72746e6f63de00000008000000, /* 2558 */
128'h7075727265746e690100000002000000, /* 2559 */
128'h3030634072656c6c6f72746e6f632d74, /* 2560 */
128'h04000000030000000000000030303030, /* 2561 */
128'h04000000030000000000000000000000, /* 2562 */
128'h0c00000003000000010000008f000000, /* 2563 */
128'h003063696c702c76637369721b000000, /* 2564 */
128'h03000000a00000000000000003000000, /* 2565 */
128'h0b00000001000000ca00000010000000, /* 2566 */
128'h10000000030000000900000001000000, /* 2567 */
128'h000000000000000c0000000067000000, /* 2568 */
128'he8000000040000000300000000000004, /* 2569 */
128'hfb000000040000000300000007000000, /* 2570 */
128'hb5000000040000000300000003000000, /* 2571 */
128'hbb000000040000000300000002000000, /* 2572 */
128'h75626564010000000200000002000000, /* 2573 */
128'h0000304072656c6c6f72746e6f632d67, /* 2574 */
128'h637369721b0000001000000003000000, /* 2575 */
128'h03000000003331302d67756265642c76, /* 2576 */
128'hffff000001000000ca00000008000000, /* 2577 */
128'h00000000670000001000000003000000, /* 2578 */
128'h03000000001000000000000000000000, /* 2579 */
128'h006c6f72746e6f63de00000008000000, /* 2580 */
128'h30303140747261750100000002000000, /* 2581 */
128'h08000000030000000000003030303030, /* 2582 */
128'h03000000003035373631736e1b000000, /* 2583 */
128'h00000010000000006700000010000000, /* 2584 */
128'h04000000030000000010000000000000, /* 2585 */
128'h040000000300000080f0fa024b000000, /* 2586 */
128'h040000000300000000c2010006010000, /* 2587 */
128'h04000000030000000200000014010000, /* 2588 */
128'h04000000030000000100000025010000, /* 2589 */
128'h04000000030000000200000030010000, /* 2590 */
128'h0100000002000000040000003a010000, /* 2591 */
128'h3030303240636d6d2d63736972776f6c, /* 2592 */
128'h10000000030000000000000030303030, /* 2593 */
128'h00000000000000200000000067000000, /* 2594 */
128'h14010000040000000300000000000100, /* 2595 */
128'h25010000040000000300000002000000, /* 2596 */
128'h1b0000000c0000000300000002000000, /* 2597 */
128'h0200000000636d6d2d63736972776f6c, /* 2598 */
128'h406874652d63736972776f6c01000000, /* 2599 */
128'h03000000000000003030303030303033, /* 2600 */
128'h2d63736972776f6c1b0000000c000000, /* 2601 */
128'h5b000000080000000300000000687465, /* 2602 */
128'h0400000003000000006b726f7774656e, /* 2603 */
128'h04000000030000000200000014010000, /* 2604 */
128'h06000000030000000300000025010000, /* 2605 */
128'h0300000000007fe3023e180047010000, /* 2606 */
128'h00000030000000006700000010000000, /* 2607 */
128'h01000000020000000080000000000000, /* 2608 */
128'h303440646e7277682d63736972776f6c, /* 2609 */
128'h0e000000030000000000303030303030, /* 2610 */
128'h6e7277682d63736972776f6c1b000000, /* 2611 */
128'h67000000100000000300000000000064, /* 2612 */
128'h00100000000000000000004000000000, /* 2613 */
128'h09000000020000000200000002000000, /* 2614 */
128'h2300736c6c65632d7373657264646123, /* 2615 */
128'h61706d6f6300736c6c65632d657a6973, /* 2616 */
128'h6f647473006c65646f6d00656c626974, /* 2617 */
128'h65736162656d697400687461702d7475, /* 2618 */
128'h6b636f6c630079636e6575716572662d, /* 2619 */
128'h63697665640079636e6575716572662d, /* 2620 */
128'h75746174730067657200657079745f65, /* 2621 */
128'h2d756d6d006173692c76637369720073, /* 2622 */
128'h230074696c70732d626c740065707974, /* 2623 */
128'h00736c6c65632d747075727265746e69, /* 2624 */
128'h6f72746e6f632d747075727265746e69, /* 2625 */
128'h646e6168702c78756e696c0072656c6c, /* 2626 */
128'h727265746e69007365676e617200656c, /* 2627 */
128'h6572006465646e657478652d73747075, /* 2628 */
128'h616d2c76637369720073656d616e2d67, /* 2629 */
128'h766373697200797469726f6972702d78, /* 2630 */
128'h70732d746e6572727563007665646e2c, /* 2631 */
128'h61702d747075727265746e6900646565, /* 2632 */
128'h0073747075727265746e6900746e6572, /* 2633 */
128'h6f692d6765720074666968732d676572, /* 2634 */
128'h63616d2d6c61636f6c0068746469772d, /* 2635 */
128'h0000000000000000737365726464612d, /* 2636 */
128'h0000000000203a642520656369766544, /* 2637 */
128'h00203a6425206563697665642073250a, /* 2638 */
128'h00000000203a6425206563697665440a, /* 2639 */
128'h000a656369766564206e776f6e6b6e75, /* 2640 */
128'h00000a2973252c73252870756b6f6f6c, /* 2641 */
128'h7265206c616e7265746e692070636864, /* 2642 */
128'h00000000000000000a7025202c726f72, /* 2643 */
128'h5145525f5043484420676e69646e6553, /* 2644 */
128'h4b434120504348440000000a54534555, /* 2645 */
128'h696c432050434844000000000000000a, /* 2646 */
128'h203a7373657264644120504920746e65, /* 2647 */
128'h0000000a64252e64252e64252e642520, /* 2648 */
128'h73657264644120504920726576726553, /* 2649 */
128'h0a64252e64252e64252e642520203a73, /* 2650 */
128'h6120726574756f520000000000000000, /* 2651 */
128'h252e64252e642520203a737365726464, /* 2652 */
128'h6b73616d2074654e0000000a64252e64, /* 2653 */
128'h64252e642520203a7373657264646120, /* 2654 */
128'h697420657361654c000a64252e64252e, /* 2655 */
128'h7364253a6d64253a686425203d20656d, /* 2656 */
128'h3d206e69616d6f44000000000000000a, /* 2657 */
128'h4820746e65696c4300000a2273252220, /* 2658 */
128'h000a22732522203d20656d616e74736f, /* 2659 */
128'h000000000a44455050494b53204b4341, /* 2660 */
128'h000000000000000a4b414e2050434844, /* 2661 */
128'h73657264646120646574736575716552, /* 2662 */
128'h0000000000000a646573756665722073, /* 2663 */
128'h000000000000000a732520726f727245, /* 2664 */
128'h6e6f6974706f2064656c646e61686e75, /* 2665 */
128'h656c646e61686e55000000000a642520, /* 2666 */
128'h64252065646f63706f20504348442064, /* 2667 */
128'h20676e69646e6553000000000000000a, /* 2668 */
128'h000a595245564f435349445f50434844, /* 2669 */
128'h00000000000a29732528726f72726570, /* 2670 */
128'h3a2043414d2073250000000030687465, /* 2671 */
128'h3a583230253a583230253a5832302520, /* 2672 */
128'h000a583230253a583230253a58323025, /* 2673 */
128'h484420646e65732074276e646c756f43, /* 2674 */
128'h206e6f20595245564f43534944205043, /* 2675 */
128'h00000a7325203a732520656369766564, /* 2676 */
128'h5043484420726f6620676e6974696157, /* 2677 */
128'h2020202020202020000a524546464f5f, /* 2678 */
128'h00000000000063250000000000000020, /* 2679 */
128'h0000005832302520000000000000002e, /* 2680 */
128'h00000000732573250000000000000a0a, /* 2681 */
128'h00000000007325203a646c697542202c, /* 2682 */
128'h73257a4820756c250000000000007325, /* 2683 */
128'h0000000000756c250000000000000000, /* 2684 */
128'h0073257a4863252000000000646c252e, /* 2685 */
128'h00000000007325736574794220756c25, /* 2686 */
128'h00003a786c3830250073254269632520, /* 2687 */
128'h000a73252020202000786c6c2a302520, /* 2688 */
128'h000000203a5d64255b6e6f6974636553, /* 2689 */
128'h25203d206465726975716572206e656c, /* 2690 */
128'h000a7825203d206c6175746361202c58, /* 2691 */
128'h302c782578302c7825287970636d656d, /* 2692 */
128'h25287465736d656d00000a3b29782578, /* 2693 */
128'h00000000000a3b29782578302c302c78, /* 2694 */
128'h0000000054455346464f5f4f4c43414d, /* 2695 */
128'h0000000054455346464f5f494843414d, /* 2696 */
128'h000000000054455346464f5f524c5054, /* 2697 */
128'h000000000054455346464f5f53434654, /* 2698 */
128'h0054455346464f5f4c5254434f49444d, /* 2699 */
128'h000000000054455346464f5f53434652, /* 2700 */
128'h00000000000054455346464f5f525352, /* 2701 */
128'h000000000054455346464f5f44414252, /* 2702 */
128'h000000000054455346464f5f524c5052, /* 2703 */
128'h46464f5f524c5052000000003f3f3f3f, /* 2704 */
128'h0000000000000047000064252b544553, /* 2705 */
128'h0a50495049203d206f746f7250205049, /* 2706 */
128'h00000000000000540000000000000000, /* 2707 */
128'h000a504745203d206f746f7250205049, /* 2708 */
128'h000a505550203d206f746f7250205049, /* 2709 */
128'h0000000a3a7265646165682074736574, /* 2710 */
128'h000a3a73746e65746e6f632074736574, /* 2711 */
128'h000a504449203d206f746f7250205049, /* 2712 */
128'h00000a5054203d206f746f7250205049, /* 2713 */
128'h0a50434344203d206f746f7250205049, /* 2714 */
128'h00000000000000360000000000000000, /* 2715 */
128'h0a50565352203d206f746f7250205049, /* 2716 */
128'h6f746f72502050490000000000000000, /* 2717 */
128'h6f746f7250205049000a455247203d20, /* 2718 */
128'h6f746f7250205049000a505345203d20, /* 2719 */
128'h6f746f725020504900000a4841203d20, /* 2720 */
128'h6f746f7250205049000a50544d203d20, /* 2721 */
128'h0000000000000a485054454542203d20, /* 2722 */
128'h5041434e45203d206f746f7250205049, /* 2723 */
128'h000000000000004d000000000000000a, /* 2724 */
128'h0a504d4f43203d206f746f7250205049, /* 2725 */
128'h6f746f72502050490000000000000000, /* 2726 */
128'h00000000000000000a50544353203d20, /* 2727 */
128'h494c504455203d206f746f7250205049, /* 2728 */
128'h6f746f725020504900000000000a4554, /* 2729 */
128'h00000000000000000a534c504d203d20, /* 2730 */
128'h000a574152203d206f746f7250205049, /* 2731 */
128'h7075736e75203d206f746f7270205049, /* 2732 */
128'h000000000a2978252820646574726f70, /* 2733 */
128'h257830203d20657079745f6f746f7270, /* 2734 */
128'h656c646e61686e750000000000000a78, /* 2735 */
128'h0000000a21747075727265746e692064, /* 2736 */
128'h000a726464612043414d207075746553, /* 2737 */
128'h00000a786c253a786c25203d2043414d, /* 2738 */
128'h3025203d20737365726464612043414d, /* 2739 */
128'h3230253a783230253a783230253a7832, /* 2740 */
128'h0000000a2e783230253a783230253a78, /* 2741 */
128'h75727265746e692074656e7265687445, /* 2742 */
128'h0a646c25203d20737574617473207470, /* 2743 */
128'h65687420746f6f420000000000000000, /* 2744 */
128'h2e6d6172676f727020646564616f6c20, /* 2745 */
128'h2c657962646f6f4700000000000a2e2e, /* 2746 */
128'h000000000a2e2e2e207265746f6f6220, /* 2747 */
128'h00007f7c5d5b3f3e3d3c3b3a2c2b2a22, /* 2748 */
128'h007f7c5d5b3f3e3d3c3b3a2e2c2b2a22, /* 2749 */
128'h66656463626139383736353433323130, /* 2750 */
128'h72776f6c2f6372730000000000000000, /* 2751 */
128'h00000000000000632e636d6d5f637369, /* 2752 */
128'h61625f6473203d3d20657361625f6473, /* 2753 */
128'h5f63736972776f6c00726464615f6573, /* 2754 */
128'h000a74756f656d6974207325203a6473, /* 2755 */
128'h616d202c6465766f6d65722064726143, /* 2756 */
128'h6425206f74206465676e616863206b73, /* 2757 */
128'h736e692064726143000000000000000a, /* 2758 */
128'h6e616863206b73616d202c6465747265, /* 2759 */
128'h0000000000000a6425206f7420646567, /* 2760 */
128'h25207461206465746165726320636d6d, /* 2761 */
128'h0000000a7825203d2074736f68202c78, /* 2762 */
128'h0000000000006f4e0000000000736559, /* 2763 */
128'h002020203a434d4d0000000052444420, /* 2764 */
128'h00000000000a7325203a656369766544, /* 2765 */
128'h3a4449207265727574636166756e614d, /* 2766 */
128'h0a7825203a4d454f000000000a782520, /* 2767 */
128'h6325203a656d614e0000000000000000, /* 2768 */
128'h0000000000000a206325632563256325, /* 2769 */
128'h00000a6425203a646565705320737542, /* 2770 */
128'h25203a79746963617061432068676948, /* 2771 */
128'h79746963617061430000000000000a73, /* 2772 */
128'h7464695720737542000000000000203a, /* 2773 */
128'h000000000a73257469622d6425203a68, /* 2774 */
128'h0000007825782520000000203a78250a, /* 2775 */
128'h00000000000064735f63736972776f6c, /* 2776 */
128'h0000000065646f6d206e776f6e6b6e55, /* 2777 */
128'h7830203a726f72724520737574617453, /* 2778 */
128'h2074756f656d69540000000a58383025, /* 2779 */
128'h616572206472616320676e6974696177, /* 2780 */
128'h6c69616620636d6d00000000000a7964, /* 2781 */
128'h6d6320706f747320646e6573206f7420, /* 2782 */
128'h6f6c62203a434d4d0000000000000a64, /* 2783 */
128'h20786c257830207265626d756e206b63, /* 2784 */
128'h6c2578302878616d2073646565637865, /* 2785 */
128'h203d3e20434d4d6500000000000a2978, /* 2786 */
128'h726f6620646572697571657220342e34, /* 2787 */
128'h642072657375206465636e61686e6520, /* 2788 */
128'h000000000000000a6165726120617461, /* 2789 */
128'h757320746f6e2073656f642064726143, /* 2790 */
128'h696e6f697469747261702074726f7070, /* 2791 */
128'h656f64206472614300000000000a676e, /* 2792 */
128'h20434820656e6966656420746f6e2073, /* 2793 */
128'h00000a657a69732070756f7267205057, /* 2794 */
128'h636e61686e6520617461642072657355, /* 2795 */
128'h5720434820746f6e2061657261206465, /* 2796 */
128'h696c6120657a69732070756f72672050, /* 2797 */
128'h72617020692550470000000a64656e67, /* 2798 */
128'h505720434820746f6e206e6f69746974, /* 2799 */
128'h67696c6120657a69732070756f726720, /* 2800 */
128'h656f642064726143000000000a64656e, /* 2801 */
128'h6e652074726f7070757320746f6e2073, /* 2802 */
128'h657475626972747461206465636e6168, /* 2803 */
128'h6e65206c61746f54000000000000000a, /* 2804 */
128'h6563786520657a6973206465636e6168, /* 2805 */
128'h20752528206d756d6978616d20736465, /* 2806 */
128'h656f64206472614300000a297525203e, /* 2807 */
128'h6f682074726f7070757320746f6e2073, /* 2808 */
128'h61702064656c6c6f72746e6f63207473, /* 2809 */
128'h6572206574697277206e6f6974697472, /* 2810 */
128'h6e6974746573207974696c696261696c, /* 2811 */
128'h726c61206472614300000000000a7367, /* 2812 */
128'h64656e6f697469747261702079646165, /* 2813 */
128'h206f6e203a434d4d000000000000000a, /* 2814 */
128'h0000000a746e65736572702064726163, /* 2815 */
128'h73657220746f6e206469642064726143, /* 2816 */
128'h20656761746c6f76206f7420646e6f70, /* 2817 */
128'h00000000000000000a217463656c6573, /* 2818 */
128'h7463656c6573206f7420656c62616e75, /* 2819 */
128'h00000000000000000a65646f6d206120, /* 2820 */
128'h646e756f66206473635f747865206f4e, /* 2821 */
128'h78363025206e614d0000000000000a21, /* 2822 */
128'h000000783430257834302520726e5320, /* 2823 */
128'h00000000632563256325632563256325, /* 2824 */
128'h6167656c20434d4d00000064252e6425, /* 2825 */
128'h636167654c2044530000000000007963, /* 2826 */
128'h6867694820434d4d0000000000000079, /* 2827 */
128'h0000297a484d36322820646565705320, /* 2828 */
128'h35282064656570532068676948204453, /* 2829 */
128'h6867694820434d4d000000297a484d30, /* 2830 */
128'h0000297a484d32352820646565705320, /* 2831 */
128'h7a484d32352820323552444420434d4d, /* 2832 */
128'h31524453205348550000000000000029, /* 2833 */
128'h00000000000000297a484d3532282032, /* 2834 */
128'h7a484d30352820353252445320534855, /* 2835 */
128'h35524453205348550000000000000029, /* 2836 */
128'h000000000000297a484d303031282030, /* 2837 */
128'h7a484d30352820303552444420534855, /* 2838 */
128'h31524453205348550000000000000029, /* 2839 */
128'h0000000000297a484d38303228203430, /* 2840 */
128'h0000297a484d30303228203030325348, /* 2841 */
128'h6f6e2064252065636976654420434d4d, /* 2842 */
128'h00000000000000000a646e756f662074, /* 2843 */
128'h000000000000445300000000434d4d65, /* 2844 */
128'h000000297325282000006425203a7325, /* 2845 */
128'h6e656c20656c69460000000000636d6d, /* 2846 */
128'h000000000000000a6425203d20687467, /* 2847 */
128'h0a7325203d202964252c70252835646d, /* 2848 */
128'h20747365757165520000000000000000, /* 2849 */
128'h25202e676e6f6c206f6f742068746170, /* 2850 */
128'h000000000000002f00000000000a646c, /* 2851 */
128'h6b636f6c62202c22732522203a717277, /* 2852 */
128'h00000000000000000a64253d657a6973, /* 2853 */
128'h646e6520656c69662065766965636552, /* 2854 */
128'h775f656c646e61680000000000000a2e, /* 2855 */
128'h00000000000a2e64656c6c6163207172, /* 2856 */
128'h65706f2050544654206c6167656c6c49, /* 2857 */
128'h00000000000000000a2e6e6f69746172, /* 2858 */
128'h445320746e756f6d206f74206c696146, /* 2859 */
128'h000000000000000a2172657669726420, /* 2860 */
128'h6e69206e69622e746f6f622064616f4c, /* 2861 */
128'h0000000000000a79726f6d656d206f74, /* 2862 */
128'h00000000000000006e69622e746f6f62, /* 2863 */
128'h62206e65706f206f742064656c696146, /* 2864 */
128'h206f74206c6961660000000a21746f6f, /* 2865 */
128'h000000000021656c69662065736f6c63, /* 2866 */
128'h6420746e756f6d75206f74206c696166, /* 2867 */
128'h2520646564616f4c00000000216b7369, /* 2868 */
128'h726f6d656d206f742073657479622064, /* 2869 */
128'h6f726620782520737365726464612079, /* 2870 */
128'h642520666f206e69622e746f6f62206d, /* 2871 */
128'h00000000000000000a2e736574796220, /* 2872 */
128'h20524444206f7420666c652064616f6c, /* 2873 */
128'h6461657220666c65000a79726f6d656d, /* 2874 */
128'h646f6320687469772064656c69616620, /* 2875 */
128'h000000005c2d2f7c0000000064252065, /* 2876 */
128'h696620646573616220746f6f622d750a, /* 2877 */
128'h6c20746f6f6220656761747320747372, /* 2878 */
128'h6f6974726573736100000a726564616f, /* 2879 */
128'h6c6966202c64656c696166207325206e, /* 2880 */
128'h66202c642520656e696c202c73252065, /* 2881 */
128'h00000000000a7325206e6f6974636e75, /* 2882 */
128'h3d212078257830203a4552554c494146, /* 2883 */
128'h2074657366666f207461207825783020, /* 2884 */
128'h2c7025203d20317000000a2e78257830, /* 2885 */
128'h000000000000000a7025203d20327020, /* 2886 */
128'h00000000002020202020202020202020, /* 2887 */
128'h00000000000808080808080808080808, /* 2888 */
128'h000000000000752520676e6974746573, /* 2889 */
128'h000000000000752520676e6974736574, /* 2890 */
128'h6c626973736f70203a4552554c494146, /* 2891 */
128'h696c2073736572646461206461622065, /* 2892 */
128'h2578302074657366666f20746120656e, /* 2893 */
128'h676e697070696b5300000000000a2e78, /* 2894 */
128'h2e2e2e74736574207478656e206f7420, /* 2895 */
128'h0808080808080808000000000000000a, /* 2896 */
128'h08082020202020202020202020080808, /* 2897 */
128'h00000000000000080808080808080808, /* 2898 */
128'h6e617220747365740000000000082008, /* 2899 */
128'h7830206f742070257830207369206567, /* 2900 */
128'h00752520706f6f4c00000000000a7025, /* 2901 */
128'h0000000000000a3a000000000075252f, /* 2902 */
128'h00000073736572646441206b63757453, /* 2903 */
128'h00000000000a6b6f0000203a73252020, /* 2904 */
128'h656d20657261420a00000a2e656e6f44, /* 2905 */
128'h00000a74736574204d415244206c6174, /* 2906 */
128'h6f6973726576207265747365746d656d, /* 2907 */
128'h297469622d64252820302e332e34206e, /* 2908 */
128'h6867697279706f43000000000000000a, /* 2909 */
128'h20323130322d31303032202943282074, /* 2910 */
128'h2e6e6f62617a61432073656c72616843, /* 2911 */
128'h6465736e6563694c000000000000000a, /* 2912 */
128'h4720554e4720656874207265646e7520, /* 2913 */
128'h694c2063696c627550206c6172656e65, /* 2914 */
128'h2032206e6f69737265762065736e6563, /* 2915 */
128'h00000000000000000a2e29796c6e6f28, /* 2916 */
128'h6425203d207465735f676e696b726f77, /* 2917 */
128'h7463757274736e6920646c25202c424b, /* 2918 */
128'h73656c63796320646c25202c736e6f69, /* 2919 */
128'h0a646c252e646c25203d20495043202c, /* 2920 */
128'h6f57206f6c6c65480000000000000000, /* 2921 */
128'h205d64255b70777300000a0d21646c72, /* 2922 */
128'h4d454f20495053510000000a5825203d, /* 2923 */
128'h0000000000000a7825203d205d64255b, /* 2924 */
128'h3d20676e697474657320686374697753, /* 2925 */
128'h73206d6f646e6152000a58252c582520, /* 2926 */
128'h000000000000000a5825203d20646565, /* 2927 */
128'h00000000000000000a746f6f62204453, /* 2928 */
128'h0000000000000a74736574204d415244, /* 2929 */
128'h0000000000000a746f6f622050544654, /* 2930 */
128'h00000000000a74736574206568636143, /* 2931 */
128'hcccccccccccccccd00000a0d70617274, /* 2932 */
128'h1032547698badcfeefcdab8967452301, /* 2933 */
128'h5851f42d4c957f2d1000000020000000, /* 2934 */
128'haaaaaaaaaaaaaaaa5555555555555555, /* 2935 */
128'h00000000000000000000000000000000, /* 2936 */
128'h00000000000000000000000000000000, /* 2937 */
128'h00000000000000000000000000000000, /* 2938 */
128'h00000000000000000000000000000000, /* 2939 */
128'h00000000000000000000000000000000, /* 2940 */
128'h00000000000000000000000000000000, /* 2941 */
128'h00000000000000000000000000000000, /* 2942 */
128'h00000000000000000000000000000000, /* 2943 */
128'h00004b4d47545045000000030f060301, /* 2944 */
128'h000000003000000000000000004b4d47, /* 2945 */
128'h00000000ffffffff0000000000000000, /* 2946 */
128'h0000646d635f6473000000000c000000, /* 2947 */
128'h00000000ffffffff00006772615f6473, /* 2948 */
128'h000000002f7c5c2d00000000bffeb028, /* 2949 */
128'h0000000600000000bffeb1e0cc33aa55, /* 2950 */
128'hbffe709e0000000000000000ffffffff, /* 2951 */
128'h00000000000000000000000000000000, /* 2952 */
128'h00000000000000000000000000000000, /* 2953 */
128'h00000000000000000000000000000000, /* 2954 */
128'h00000000000000000000000000000000, /* 2955 */
128'h00000000000000000000000000000000, /* 2956 */
128'h00000000000000000000000000000000, /* 2957 */
128'h00000000000000000000000000000000, /* 2958 */
128'h00000000000000000000000000000000, /* 2959 */
128'h00000000000000000000000000000000, /* 2960 */
128'h00000000000000000000000000000000, /* 2961 */
128'h00000000000000000000000000000000, /* 2962 */
128'h00000000000000000000000000000000, /* 2963 */
128'h00000000000000000000000000000000, /* 2964 */
128'h00000000000000000000000000000000, /* 2965 */
128'h00000000000000000000000000000000, /* 2966 */
128'h00000000000000000000000000000000, /* 2967 */
128'h00000000000000000000000000000000, /* 2968 */
128'h00000000000000000000000000000000, /* 2969 */
128'h00000000000000000000000000000000, /* 2970 */
128'h00000000000000000000000000000000, /* 2971 */
128'h00000000000000000000000000000000, /* 2972 */
128'h00000000000000000000000000000000, /* 2973 */
128'h00000000000000000000000000000000, /* 2974 */
128'h00000000000000000000000000000000, /* 2975 */
128'h00000000000000000000000000000000, /* 2976 */
128'h00000000000000000000000000000000, /* 2977 */
128'h00000000000000000000000000000000, /* 2978 */
128'h00000000000000000000000000000000, /* 2979 */
128'h00000000000000000000000000000000, /* 2980 */
128'h00000000000000000000000000000000, /* 2981 */
128'h00000000000000000000000000000000, /* 2982 */
128'h00000000000000000000000000000000, /* 2983 */
128'h00000000000000000000000000000000, /* 2984 */
128'h00000000000000000000000000000000, /* 2985 */
128'h00000000000000000000000000000000, /* 2986 */
128'h00000000000000000000000000000000, /* 2987 */
128'h00000000000000000000000000000000, /* 2988 */
128'h00000000000000000000000000000000, /* 2989 */
128'h00000000000000000000000000000000, /* 2990 */
128'h00000000000000000000000000000000, /* 2991 */
128'h00000000000000000000000000000000, /* 2992 */
128'h00000000000000000000000000000000, /* 2993 */
128'h00000000000000000000000000000000, /* 2994 */
128'h00000000000000000000000000000000, /* 2995 */
128'h00000000000000000000000000000000, /* 2996 */
128'h00000000000000000000000000000000, /* 2997 */
128'h00000000000000000000000000000000, /* 2998 */
128'h00000000000000000000000000000000, /* 2999 */
128'h00000000000000000000000000000000, /* 3000 */
128'h00000000000000000000000000000000, /* 3001 */
128'h00000000000000000000000000000000, /* 3002 */
128'h00000000000000000000000000000000, /* 3003 */
128'h00000000000000000000000000000000, /* 3004 */
128'h00000000000000000000000000000000, /* 3005 */
128'h00000000000000000000000000000000, /* 3006 */
128'h00000000000000000000000000000000, /* 3007 */
128'h00000000000000000000000000000000, /* 3008 */
128'h00000000000000000000000000000000, /* 3009 */
128'h00000000000000000000000000000000, /* 3010 */
128'h00000000000000000000000000000000, /* 3011 */
128'h00000000000000000000000000000000, /* 3012 */
128'h00000000000000000000000000000000, /* 3013 */
128'h00000000000000000000000000000000, /* 3014 */
128'h00000000000000000000000000000000, /* 3015 */
128'h00000000000000000000000000000000, /* 3016 */
128'h00000000000000000000000000000000, /* 3017 */
128'h00000000000000000000000000000000, /* 3018 */
128'h00000000000000000000000000000000, /* 3019 */
128'h00000000000000000000000000000000, /* 3020 */
128'h00000000000000000000000000000000, /* 3021 */
128'h00000000000000000000000000000000, /* 3022 */
128'h00000000000000000000000000000000, /* 3023 */
128'h00000000000000000000000000000000, /* 3024 */
128'h00000000000000000000000000000000, /* 3025 */
128'h00000000000000000000000000000000, /* 3026 */
128'h00000000000000000000000000000000, /* 3027 */
128'h00000000000000000000000000000000, /* 3028 */
128'h00000000000000000000000000000000, /* 3029 */
128'h00000000000000000000000000000000, /* 3030 */
128'h00000000000000000000000000000000, /* 3031 */
128'h00000000000000000000000000000000, /* 3032 */
128'h00000000000000000000000000000000, /* 3033 */
128'h00000000000000000000000000000000, /* 3034 */
128'h00000000000000000000000000000000, /* 3035 */
128'h00000000000000000000000000000000, /* 3036 */
128'h00000000000000000000000000000000, /* 3037 */
128'h00000000000000000000000000000000, /* 3038 */
128'h00000000000000000000000000000000, /* 3039 */
128'h00000000000000000000000000000000, /* 3040 */
128'h00000000000000000000000000000000, /* 3041 */
128'h00000000000000000000000000000000, /* 3042 */
128'h00000000000000000000000000000000, /* 3043 */
128'h00000000000000000000000000000000, /* 3044 */
128'h00000000000000000000000000000000, /* 3045 */
128'h00000000000000000000000000000000, /* 3046 */
128'h00000000000000000000000000000000, /* 3047 */
128'h00000000000000000000000000000000, /* 3048 */
128'h00000000000000000000000000000000, /* 3049 */
128'h00000000000000000000000000000000, /* 3050 */
128'h00000000000000000000000000000000, /* 3051 */
128'h00000000000000000000000000000000, /* 3052 */
128'h00000000000000000000000000000000, /* 3053 */
128'h00000000000000000000000000000000, /* 3054 */
128'h00000000000000000000000000000000, /* 3055 */
128'h00000000000000000000000000000000, /* 3056 */
128'h00000000000000000000000000000000, /* 3057 */
128'h00000000000000000000000000000000, /* 3058 */
128'h00000000000000000000000000000000, /* 3059 */
128'h00000000000000000000000000000000, /* 3060 */
128'h00000000000000000000000000000000, /* 3061 */
128'h00000000000000000000000000000000, /* 3062 */
128'h00000000000000000000000000000000, /* 3063 */
128'h00000000000000000000000000000000, /* 3064 */
128'h00000000000000000000000000000000, /* 3065 */
128'h00000000000000000000000000000000, /* 3066 */
128'h00000000000000000000000000000000, /* 3067 */
128'h00000000000000000000000000000000, /* 3068 */
128'h00000000000000000000000000000000, /* 3069 */
128'h00000000000000000000000000000000, /* 3070 */
128'h00000000000000000000000000000000, /* 3071 */
128'h00000000000000000000000000000000, /* 3072 */
128'h00000000000000000000000000000000, /* 3073 */
128'h00000000000000000000000000000000, /* 3074 */
128'h00000000000000000000000000000000, /* 3075 */
128'h00000000000000000000000000000000, /* 3076 */
128'h00000000000000000000000000000000, /* 3077 */
128'h00000000000000000000000000000000, /* 3078 */
128'h00000000000000000000000000000000, /* 3079 */
128'h00000000000000000000000000000000, /* 3080 */
128'h00000000000000000000000000000000, /* 3081 */
128'h00000000000000000000000000000000, /* 3082 */
128'h00000000000000000000000000000000, /* 3083 */
128'h00000000000000000000000000000000, /* 3084 */
128'h00000000000000000000000000000000, /* 3085 */
128'h00000000000000000000000000000000, /* 3086 */
128'h00000000000000000000000000000000, /* 3087 */
128'h00000000000000000000000000000000, /* 3088 */
128'h00000000000000000000000000000000, /* 3089 */
128'h00000000000000000000000000000000, /* 3090 */
128'h00000000000000000000000000000000, /* 3091 */
128'h00000000000000000000000000000000, /* 3092 */
128'h00000000000000000000000000000000, /* 3093 */
128'h00000000000000000000000000000000, /* 3094 */
128'h00000000000000000000000000000000, /* 3095 */
128'h00000000000000000000000000000000, /* 3096 */
128'h00000000000000000000000000000000, /* 3097 */
128'h00000000000000000000000000000000, /* 3098 */
128'h00000000000000000000000000000000, /* 3099 */
128'h00000000000000000000000000000000, /* 3100 */
128'h00000000000000000000000000000000, /* 3101 */
128'h00000000000000000000000000000000, /* 3102 */
128'h00000000000000000000000000000000, /* 3103 */
128'h00000000000000000000000000000000, /* 3104 */
128'h00000000000000000000000000000000, /* 3105 */
128'h00000000000000000000000000000000, /* 3106 */
128'h00000000000000000000000000000000, /* 3107 */
128'h00000000000000000000000000000000, /* 3108 */
128'h00000000000000000000000000000000, /* 3109 */
128'h00000000000000000000000000000000, /* 3110 */
128'h00000000000000000000000000000000, /* 3111 */
128'h00000000000000000000000000000000, /* 3112 */
128'h00000000000000000000000000000000, /* 3113 */
128'h00000000000000000000000000000000, /* 3114 */
128'h00000000000000000000000000000000, /* 3115 */
128'h00000000000000000000000000000000, /* 3116 */
128'h00000000000000000000000000000000, /* 3117 */
128'h00000000000000000000000000000000, /* 3118 */
128'h00000000000000000000000000000000, /* 3119 */
128'h00000000000000000000000000000000, /* 3120 */
128'h00000000000000000000000000000000, /* 3121 */
128'h00000000000000000000000000000000, /* 3122 */
128'h00000000000000000000000000000000, /* 3123 */
128'h00000000000000000000000000000000, /* 3124 */
128'h00000000000000000000000000000000, /* 3125 */
128'h00000000000000000000000000000000, /* 3126 */
128'h00000000000000000000000000000000, /* 3127 */
128'h00000000000000000000000000000000, /* 3128 */
128'h00000000000000000000000000000000, /* 3129 */
128'h00000000000000000000000000000000, /* 3130 */
128'h00000000000000000000000000000000, /* 3131 */
128'h00000000000000000000000000000000, /* 3132 */
128'h00000000000000000000000000000000, /* 3133 */
128'h00000000000000000000000000000000, /* 3134 */
128'h00000000000000000000000000000000, /* 3135 */
128'h00000000000000000000000000000000, /* 3136 */
128'h00000000000000000000000000000000, /* 3137 */
128'h00000000000000000000000000000000, /* 3138 */
128'h00000000000000000000000000000000, /* 3139 */
128'h00000000000000000000000000000000, /* 3140 */
128'h00000000000000000000000000000000, /* 3141 */
128'h00000000000000000000000000000000, /* 3142 */
128'h00000000000000000000000000000000, /* 3143 */
128'h00000000000000000000000000000000, /* 3144 */
128'h00000000000000000000000000000000, /* 3145 */
128'h00000000000000000000000000000000, /* 3146 */
128'h00000000000000000000000000000000, /* 3147 */
128'h00000000000000000000000000000000, /* 3148 */
128'h00000000000000000000000000000000, /* 3149 */
128'h00000000000000000000000000000000, /* 3150 */
128'h00000000000000000000000000000000, /* 3151 */
128'h00000000000000000000000000000000, /* 3152 */
128'h00000000000000000000000000000000, /* 3153 */
128'h00000000000000000000000000000000, /* 3154 */
128'h00000000000000000000000000000000, /* 3155 */
128'h00000000000000000000000000000000, /* 3156 */
128'h00000000000000000000000000000000, /* 3157 */
128'h00000000000000000000000000000000, /* 3158 */
128'h00000000000000000000000000000000, /* 3159 */
128'h00000000000000000000000000000000, /* 3160 */
128'h00000000000000000000000000000000, /* 3161 */
128'h00000000000000000000000000000000, /* 3162 */
128'h00000000000000000000000000000000, /* 3163 */
128'h00000000000000000000000000000000, /* 3164 */
128'h00000000000000000000000000000000, /* 3165 */
128'h00000000000000000000000000000000, /* 3166 */
128'h00000000000000000000000000000000, /* 3167 */
128'h00000000000000000000000000000000, /* 3168 */
128'h00000000000000000000000000000000, /* 3169 */
128'h00000000000000000000000000000000, /* 3170 */
128'h00000000000000000000000000000000, /* 3171 */
128'h00000000000000000000000000000000, /* 3172 */
128'h00000000000000000000000000000000, /* 3173 */
128'h00000000000000000000000000000000, /* 3174 */
128'h00000000000000000000000000000000, /* 3175 */
128'h00000000000000000000000000000000, /* 3176 */
128'h00000000000000000000000000000000, /* 3177 */
128'h00000000000000000000000000000000, /* 3178 */
128'h00000000000000000000000000000000, /* 3179 */
128'h00000000000000000000000000000000, /* 3180 */
128'h00000000000000000000000000000000, /* 3181 */
128'h00000000000000000000000000000000, /* 3182 */
128'h00000000000000000000000000000000, /* 3183 */
128'h00000000000000000000000000000000, /* 3184 */
128'h00000000000000000000000000000000, /* 3185 */
128'h00000000000000000000000000000000, /* 3186 */
128'h00000000000000000000000000000000, /* 3187 */
128'h00000000000000000000000000000000, /* 3188 */
128'h00000000000000000000000000000000, /* 3189 */
128'h00000000000000000000000000000000, /* 3190 */
128'h00000000000000000000000000000000, /* 3191 */
128'h00000000000000000000000000000000, /* 3192 */
128'h00000000000000000000000000000000, /* 3193 */
128'h00000000000000000000000000000000, /* 3194 */
128'h00000000000000000000000000000000, /* 3195 */
128'h00000000000000000000000000000000, /* 3196 */
128'h00000000000000000000000000000000, /* 3197 */
128'h00000000000000000000000000000000, /* 3198 */
128'h00000000000000000000000000000000, /* 3199 */
128'h00000000000000000000000000000000, /* 3200 */
128'h00000000000000000000000000000000, /* 3201 */
128'h00000000000000000000000000000000, /* 3202 */
128'h00000000000000000000000000000000, /* 3203 */
128'h00000000000000000000000000000000, /* 3204 */
128'h00000000000000000000000000000000, /* 3205 */
128'h00000000000000000000000000000000, /* 3206 */
128'h00000000000000000000000000000000, /* 3207 */
128'h00000000000000000000000000000000, /* 3208 */
128'h00000000000000000000000000000000, /* 3209 */
128'h00000000000000000000000000000000, /* 3210 */
128'h00000000000000000000000000000000, /* 3211 */
128'h00000000000000000000000000000000, /* 3212 */
128'h00000000000000000000000000000000, /* 3213 */
128'h00000000000000000000000000000000, /* 3214 */
128'h00000000000000000000000000000000, /* 3215 */
128'h00000000000000000000000000000000, /* 3216 */
128'h00000000000000000000000000000000, /* 3217 */
128'h00000000000000000000000000000000, /* 3218 */
128'h00000000000000000000000000000000, /* 3219 */
128'h00000000000000000000000000000000, /* 3220 */
128'h00000000000000000000000000000000, /* 3221 */
128'h00000000000000000000000000000000, /* 3222 */
128'h00000000000000000000000000000000, /* 3223 */
128'h00000000000000000000000000000000, /* 3224 */
128'h00000000000000000000000000000000, /* 3225 */
128'h00000000000000000000000000000000, /* 3226 */
128'h00000000000000000000000000000000, /* 3227 */
128'h00000000000000000000000000000000, /* 3228 */
128'h00000000000000000000000000000000, /* 3229 */
128'h00000000000000000000000000000000, /* 3230 */
128'h00000000000000000000000000000000, /* 3231 */
128'h00000000000000000000000000000000, /* 3232 */
128'h00000000000000000000000000000000, /* 3233 */
128'h00000000000000000000000000000000, /* 3234 */
128'h00000000000000000000000000000000, /* 3235 */
128'h00000000000000000000000000000000, /* 3236 */
128'h00000000000000000000000000000000, /* 3237 */
128'h00000000000000000000000000000000, /* 3238 */
128'h00000000000000000000000000000000, /* 3239 */
128'h00000000000000000000000000000000, /* 3240 */
128'h00000000000000000000000000000000, /* 3241 */
128'h00000000000000000000000000000000, /* 3242 */
128'h00000000000000000000000000000000, /* 3243 */
128'h00000000000000000000000000000000, /* 3244 */
128'h00000000000000000000000000000000, /* 3245 */
128'h00000000000000000000000000000000, /* 3246 */
128'h00000000000000000000000000000000, /* 3247 */
128'h00000000000000000000000000000000, /* 3248 */
128'h00000000000000000000000000000000, /* 3249 */
128'h00000000000000000000000000000000, /* 3250 */
128'h00000000000000000000000000000000, /* 3251 */
128'h00000000000000000000000000000000, /* 3252 */
128'h00000000000000000000000000000000, /* 3253 */
128'h00000000000000000000000000000000, /* 3254 */
128'h00000000000000000000000000000000, /* 3255 */
128'h00000000000000000000000000000000, /* 3256 */
128'h00000000000000000000000000000000, /* 3257 */
128'h00000000000000000000000000000000, /* 3258 */
128'h00000000000000000000000000000000, /* 3259 */
128'h00000000000000000000000000000000, /* 3260 */
128'h00000000000000000000000000000000, /* 3261 */
128'h00000000000000000000000000000000, /* 3262 */
128'h00000000000000000000000000000000, /* 3263 */
128'h00000000000000000000000000000000, /* 3264 */
128'h00000000000000000000000000000000, /* 3265 */
128'h00000000000000000000000000000000, /* 3266 */
128'h00000000000000000000000000000000, /* 3267 */
128'h00000000000000000000000000000000, /* 3268 */
128'h00000000000000000000000000000000, /* 3269 */
128'h00000000000000000000000000000000, /* 3270 */
128'h00000000000000000000000000000000, /* 3271 */
128'h00000000000000000000000000000000, /* 3272 */
128'h00000000000000000000000000000000, /* 3273 */
128'h00000000000000000000000000000000, /* 3274 */
128'h00000000000000000000000000000000, /* 3275 */
128'h00000000000000000000000000000000, /* 3276 */
128'h00000000000000000000000000000000, /* 3277 */
128'h00000000000000000000000000000000, /* 3278 */
128'h00000000000000000000000000000000, /* 3279 */
128'h00000000000000000000000000000000, /* 3280 */
128'h00000000000000000000000000000000, /* 3281 */
128'h00000000000000000000000000000000, /* 3282 */
128'h00000000000000000000000000000000, /* 3283 */
128'h00000000000000000000000000000000, /* 3284 */
128'h00000000000000000000000000000000, /* 3285 */
128'h00000000000000000000000000000000, /* 3286 */
128'h00000000000000000000000000000000, /* 3287 */
128'h00000000000000000000000000000000, /* 3288 */
128'h00000000000000000000000000000000, /* 3289 */
128'h00000000000000000000000000000000, /* 3290 */
128'h00000000000000000000000000000000, /* 3291 */
128'h00000000000000000000000000000000, /* 3292 */
128'h00000000000000000000000000000000, /* 3293 */
128'h00000000000000000000000000000000, /* 3294 */
128'h00000000000000000000000000000000, /* 3295 */
128'h00000000000000000000000000000000, /* 3296 */
128'h00000000000000000000000000000000, /* 3297 */
128'h00000000000000000000000000000000, /* 3298 */
128'h00000000000000000000000000000000, /* 3299 */
128'h00000000000000000000000000000000, /* 3300 */
128'h00000000000000000000000000000000, /* 3301 */
128'h00000000000000000000000000000000, /* 3302 */
128'h00000000000000000000000000000000, /* 3303 */
128'h00000000000000000000000000000000, /* 3304 */
128'h00000000000000000000000000000000, /* 3305 */
128'h00000000000000000000000000000000, /* 3306 */
128'h00000000000000000000000000000000, /* 3307 */
128'h00000000000000000000000000000000, /* 3308 */
128'h00000000000000000000000000000000, /* 3309 */
128'h00000000000000000000000000000000, /* 3310 */
128'h00000000000000000000000000000000, /* 3311 */
128'h00000000000000000000000000000000, /* 3312 */
128'h00000000000000000000000000000000, /* 3313 */
128'h00000000000000000000000000000000, /* 3314 */
128'h00000000000000000000000000000000, /* 3315 */
128'h00000000000000000000000000000000, /* 3316 */
128'h00000000000000000000000000000000, /* 3317 */
128'h00000000000000000000000000000000, /* 3318 */
128'h00000000000000000000000000000000, /* 3319 */
128'h00000000000000000000000000000000, /* 3320 */
128'h00000000000000000000000000000000, /* 3321 */
128'h00000000000000000000000000000000, /* 3322 */
128'h00000000000000000000000000000000, /* 3323 */
128'h00000000000000000000000000000000, /* 3324 */
128'h00000000000000000000000000000000, /* 3325 */
128'h00000000000000000000000000000000, /* 3326 */
128'h00000000000000000000000000000000, /* 3327 */
128'h00000000000000000000000000000000, /* 3328 */
128'h00000000000000000000000000000000, /* 3329 */
128'h00000000000000000000000000000000, /* 3330 */
128'h00000000000000000000000000000000, /* 3331 */
128'h00000000000000000000000000000000, /* 3332 */
128'h00000000000000000000000000000000, /* 3333 */
128'h00000000000000000000000000000000, /* 3334 */
128'h00000000000000000000000000000000, /* 3335 */
128'h00000000000000000000000000000000, /* 3336 */
128'h00000000000000000000000000000000, /* 3337 */
128'h00000000000000000000000000000000, /* 3338 */
128'h00000000000000000000000000000000, /* 3339 */
128'h00000000000000000000000000000000, /* 3340 */
128'h00000000000000000000000000000000, /* 3341 */
128'h00000000000000000000000000000000, /* 3342 */
128'h00000000000000000000000000000000, /* 3343 */
128'h00000000000000000000000000000000, /* 3344 */
128'h00000000000000000000000000000000, /* 3345 */
128'h00000000000000000000000000000000, /* 3346 */
128'h00000000000000000000000000000000, /* 3347 */
128'h00000000000000000000000000000000, /* 3348 */
128'h00000000000000000000000000000000, /* 3349 */
128'h00000000000000000000000000000000, /* 3350 */
128'h00000000000000000000000000000000, /* 3351 */
128'h00000000000000000000000000000000, /* 3352 */
128'h00000000000000000000000000000000, /* 3353 */
128'h00000000000000000000000000000000, /* 3354 */
128'h00000000000000000000000000000000, /* 3355 */
128'h00000000000000000000000000000000, /* 3356 */
128'h00000000000000000000000000000000, /* 3357 */
128'h00000000000000000000000000000000, /* 3358 */
128'h00000000000000000000000000000000, /* 3359 */
128'h00000000000000000000000000000000, /* 3360 */
128'h00000000000000000000000000000000, /* 3361 */
128'h00000000000000000000000000000000, /* 3362 */
128'h00000000000000000000000000000000, /* 3363 */
128'h00000000000000000000000000000000, /* 3364 */
128'h00000000000000000000000000000000, /* 3365 */
128'h00000000000000000000000000000000, /* 3366 */
128'h00000000000000000000000000000000, /* 3367 */
128'h00000000000000000000000000000000, /* 3368 */
128'h00000000000000000000000000000000, /* 3369 */
128'h00000000000000000000000000000000, /* 3370 */
128'h00000000000000000000000000000000, /* 3371 */
128'h00000000000000000000000000000000, /* 3372 */
128'h00000000000000000000000000000000, /* 3373 */
128'h00000000000000000000000000000000, /* 3374 */
128'h00000000000000000000000000000000, /* 3375 */
128'h00000000000000000000000000000000, /* 3376 */
128'h00000000000000000000000000000000, /* 3377 */
128'h00000000000000000000000000000000, /* 3378 */
128'h00000000000000000000000000000000, /* 3379 */
128'h00000000000000000000000000000000, /* 3380 */
128'h00000000000000000000000000000000, /* 3381 */
128'h00000000000000000000000000000000, /* 3382 */
128'h00000000000000000000000000000000, /* 3383 */
128'h00000000000000000000000000000000, /* 3384 */
128'h00000000000000000000000000000000, /* 3385 */
128'h00000000000000000000000000000000, /* 3386 */
128'h00000000000000000000000000000000, /* 3387 */
128'h00000000000000000000000000000000, /* 3388 */
128'h00000000000000000000000000000000, /* 3389 */
128'h00000000000000000000000000000000, /* 3390 */
128'h00000000000000000000000000000000, /* 3391 */
128'h00000000000000000000000000000000, /* 3392 */
128'h00000000000000000000000000000000, /* 3393 */
128'h00000000000000000000000000000000, /* 3394 */
128'h00000000000000000000000000000000, /* 3395 */
128'h00000000000000000000000000000000, /* 3396 */
128'h00000000000000000000000000000000, /* 3397 */
128'h00000000000000000000000000000000, /* 3398 */
128'h00000000000000000000000000000000, /* 3399 */
128'h00000000000000000000000000000000, /* 3400 */
128'h00000000000000000000000000000000, /* 3401 */
128'h00000000000000000000000000000000, /* 3402 */
128'h00000000000000000000000000000000, /* 3403 */
128'h00000000000000000000000000000000, /* 3404 */
128'h00000000000000000000000000000000, /* 3405 */
128'h00000000000000000000000000000000, /* 3406 */
128'h00000000000000000000000000000000, /* 3407 */
128'h00000000000000000000000000000000, /* 3408 */
128'h00000000000000000000000000000000, /* 3409 */
128'h00000000000000000000000000000000, /* 3410 */
128'h00000000000000000000000000000000, /* 3411 */
128'h00000000000000000000000000000000, /* 3412 */
128'h00000000000000000000000000000000, /* 3413 */
128'h00000000000000000000000000000000, /* 3414 */
128'h00000000000000000000000000000000, /* 3415 */
128'h00000000000000000000000000000000, /* 3416 */
128'h00000000000000000000000000000000, /* 3417 */
128'h00000000000000000000000000000000, /* 3418 */
128'h00000000000000000000000000000000, /* 3419 */
128'h00000000000000000000000000000000, /* 3420 */
128'h00000000000000000000000000000000, /* 3421 */
128'h00000000000000000000000000000000, /* 3422 */
128'h00000000000000000000000000000000, /* 3423 */
128'h00000000000000000000000000000000, /* 3424 */
128'h00000000000000000000000000000000, /* 3425 */
128'h00000000000000000000000000000000, /* 3426 */
128'h00000000000000000000000000000000, /* 3427 */
128'h00000000000000000000000000000000, /* 3428 */
128'h00000000000000000000000000000000, /* 3429 */
128'h00000000000000000000000000000000, /* 3430 */
128'h00000000000000000000000000000000, /* 3431 */
128'h00000000000000000000000000000000, /* 3432 */
128'h00000000000000000000000000000000, /* 3433 */
128'h00000000000000000000000000000000, /* 3434 */
128'h00000000000000000000000000000000, /* 3435 */
128'h00000000000000000000000000000000, /* 3436 */
128'h00000000000000000000000000000000, /* 3437 */
128'h00000000000000000000000000000000, /* 3438 */
128'h00000000000000000000000000000000, /* 3439 */
128'h00000000000000000000000000000000, /* 3440 */
128'h00000000000000000000000000000000, /* 3441 */
128'h00000000000000000000000000000000, /* 3442 */
128'h00000000000000000000000000000000, /* 3443 */
128'h00000000000000000000000000000000, /* 3444 */
128'h00000000000000000000000000000000, /* 3445 */
128'h00000000000000000000000000000000, /* 3446 */
128'h00000000000000000000000000000000, /* 3447 */
128'h00000000000000000000000000000000, /* 3448 */
128'h00000000000000000000000000000000, /* 3449 */
128'h00000000000000000000000000000000, /* 3450 */
128'h00000000000000000000000000000000, /* 3451 */
128'h00000000000000000000000000000000, /* 3452 */
128'h00000000000000000000000000000000, /* 3453 */
128'h00000000000000000000000000000000, /* 3454 */
128'h00000000000000000000000000000000, /* 3455 */
128'h00000000000000000000000000000000, /* 3456 */
128'h00000000000000000000000000000000, /* 3457 */
128'h00000000000000000000000000000000, /* 3458 */
128'h00000000000000000000000000000000, /* 3459 */
128'h00000000000000000000000000000000, /* 3460 */
128'h00000000000000000000000000000000, /* 3461 */
128'h00000000000000000000000000000000, /* 3462 */
128'h00000000000000000000000000000000, /* 3463 */
128'h00000000000000000000000000000000, /* 3464 */
128'h00000000000000000000000000000000, /* 3465 */
128'h00000000000000000000000000000000, /* 3466 */
128'h00000000000000000000000000000000, /* 3467 */
128'h00000000000000000000000000000000, /* 3468 */
128'h00000000000000000000000000000000, /* 3469 */
128'h00000000000000000000000000000000, /* 3470 */
128'h00000000000000000000000000000000, /* 3471 */
128'h00000000000000000000000000000000, /* 3472 */
128'h00000000000000000000000000000000, /* 3473 */
128'h00000000000000000000000000000000, /* 3474 */
128'h00000000000000000000000000000000, /* 3475 */
128'h00000000000000000000000000000000, /* 3476 */
128'h00000000000000000000000000000000, /* 3477 */
128'h00000000000000000000000000000000, /* 3478 */
128'h00000000000000000000000000000000, /* 3479 */
128'h00000000000000000000000000000000, /* 3480 */
128'h00000000000000000000000000000000, /* 3481 */
128'h00000000000000000000000000000000, /* 3482 */
128'h00000000000000000000000000000000, /* 3483 */
128'h00000000000000000000000000000000, /* 3484 */
128'h00000000000000000000000000000000, /* 3485 */
128'h00000000000000000000000000000000, /* 3486 */
128'h00000000000000000000000000000000, /* 3487 */
128'h00000000000000000000000000000000, /* 3488 */
128'h00000000000000000000000000000000, /* 3489 */
128'h00000000000000000000000000000000, /* 3490 */
128'h00000000000000000000000000000000, /* 3491 */
128'h00000000000000000000000000000000, /* 3492 */
128'h00000000000000000000000000000000, /* 3493 */
128'h00000000000000000000000000000000, /* 3494 */
128'h00000000000000000000000000000000, /* 3495 */
128'h00000000000000000000000000000000, /* 3496 */
128'h00000000000000000000000000000000, /* 3497 */
128'h00000000000000000000000000000000, /* 3498 */
128'h00000000000000000000000000000000, /* 3499 */
128'h00000000000000000000000000000000, /* 3500 */
128'h00000000000000000000000000000000, /* 3501 */
128'h00000000000000000000000000000000, /* 3502 */
128'h00000000000000000000000000000000, /* 3503 */
128'h00000000000000000000000000000000, /* 3504 */
128'h00000000000000000000000000000000, /* 3505 */
128'h00000000000000000000000000000000, /* 3506 */
128'h00000000000000000000000000000000, /* 3507 */
128'h00000000000000000000000000000000, /* 3508 */
128'h00000000000000000000000000000000, /* 3509 */
128'h00000000000000000000000000000000, /* 3510 */
128'h00000000000000000000000000000000, /* 3511 */
128'h00000000000000000000000000000000, /* 3512 */
128'h00000000000000000000000000000000, /* 3513 */
128'h00000000000000000000000000000000, /* 3514 */
128'h00000000000000000000000000000000, /* 3515 */
128'h00000000000000000000000000000000, /* 3516 */
128'h00000000000000000000000000000000, /* 3517 */
128'h00000000000000000000000000000000, /* 3518 */
128'h00000000000000000000000000000000, /* 3519 */
128'h00000000000000000000000000000000, /* 3520 */
128'h00000000000000000000000000000000, /* 3521 */
128'h00000000000000000000000000000000, /* 3522 */
128'h00000000000000000000000000000000, /* 3523 */
128'h00000000000000000000000000000000, /* 3524 */
128'h00000000000000000000000000000000, /* 3525 */
128'h00000000000000000000000000000000, /* 3526 */
128'h00000000000000000000000000000000, /* 3527 */
128'h00000000000000000000000000000000, /* 3528 */
128'h00000000000000000000000000000000, /* 3529 */
128'h00000000000000000000000000000000, /* 3530 */
128'h00000000000000000000000000000000, /* 3531 */
128'h00000000000000000000000000000000, /* 3532 */
128'h00000000000000000000000000000000, /* 3533 */
128'h00000000000000000000000000000000, /* 3534 */
128'h00000000000000000000000000000000, /* 3535 */
128'h00000000000000000000000000000000, /* 3536 */
128'h00000000000000000000000000000000, /* 3537 */
128'h00000000000000000000000000000000, /* 3538 */
128'h00000000000000000000000000000000, /* 3539 */
128'h00000000000000000000000000000000, /* 3540 */
128'h00000000000000000000000000000000, /* 3541 */
128'h00000000000000000000000000000000, /* 3542 */
128'h00000000000000000000000000000000, /* 3543 */
128'h00000000000000000000000000000000, /* 3544 */
128'h00000000000000000000000000000000, /* 3545 */
128'h00000000000000000000000000000000, /* 3546 */
128'h00000000000000000000000000000000, /* 3547 */
128'h00000000000000000000000000000000, /* 3548 */
128'h00000000000000000000000000000000, /* 3549 */
128'h00000000000000000000000000000000, /* 3550 */
128'h00000000000000000000000000000000, /* 3551 */
128'h00000000000000000000000000000000, /* 3552 */
128'h00000000000000000000000000000000, /* 3553 */
128'h00000000000000000000000000000000, /* 3554 */
128'h00000000000000000000000000000000, /* 3555 */
128'h00000000000000000000000000000000, /* 3556 */
128'h00000000000000000000000000000000, /* 3557 */
128'h00000000000000000000000000000000, /* 3558 */
128'h00000000000000000000000000000000, /* 3559 */
128'h00000000000000000000000000000000, /* 3560 */
128'h00000000000000000000000000000000, /* 3561 */
128'h00000000000000000000000000000000, /* 3562 */
128'h00000000000000000000000000000000, /* 3563 */
128'h00000000000000000000000000000000, /* 3564 */
128'h00000000000000000000000000000000, /* 3565 */
128'h00000000000000000000000000000000, /* 3566 */
128'h00000000000000000000000000000000, /* 3567 */
128'h00000000000000000000000000000000, /* 3568 */
128'h00000000000000000000000000000000, /* 3569 */
128'h00000000000000000000000000000000, /* 3570 */
128'h00000000000000000000000000000000, /* 3571 */
128'h00000000000000000000000000000000, /* 3572 */
128'h00000000000000000000000000000000, /* 3573 */
128'h00000000000000000000000000000000, /* 3574 */
128'h00000000000000000000000000000000, /* 3575 */
128'h00000000000000000000000000000000, /* 3576 */
128'h00000000000000000000000000000000, /* 3577 */
128'h00000000000000000000000000000000, /* 3578 */
128'h00000000000000000000000000000000, /* 3579 */
128'h00000000000000000000000000000000, /* 3580 */
128'h00000000000000000000000000000000, /* 3581 */
128'h00000000000000000000000000000000, /* 3582 */
128'h00000000000000000000000000000000, /* 3583 */
128'h00000000000000000000000000000000, /* 3584 */
128'h00000000000000000000000000000000, /* 3585 */
128'h00000000000000000000000000000000, /* 3586 */
128'h00000000000000000000000000000000, /* 3587 */
128'h00000000000000000000000000000000, /* 3588 */
128'h00000000000000000000000000000000, /* 3589 */
128'h00000000000000000000000000000000, /* 3590 */
128'h00000000000000000000000000000000, /* 3591 */
128'h00000000000000000000000000000000, /* 3592 */
128'h00000000000000000000000000000000, /* 3593 */
128'h00000000000000000000000000000000, /* 3594 */
128'h00000000000000000000000000000000, /* 3595 */
128'h00000000000000000000000000000000, /* 3596 */
128'h00000000000000000000000000000000, /* 3597 */
128'h00000000000000000000000000000000, /* 3598 */
128'h00000000000000000000000000000000, /* 3599 */
128'h00000000000000000000000000000000, /* 3600 */
128'h00000000000000000000000000000000, /* 3601 */
128'h00000000000000000000000000000000, /* 3602 */
128'h00000000000000000000000000000000, /* 3603 */
128'h00000000000000000000000000000000, /* 3604 */
128'h00000000000000000000000000000000, /* 3605 */
128'h00000000000000000000000000000000, /* 3606 */
128'h00000000000000000000000000000000, /* 3607 */
128'h00000000000000000000000000000000, /* 3608 */
128'h00000000000000000000000000000000, /* 3609 */
128'h00000000000000000000000000000000, /* 3610 */
128'h00000000000000000000000000000000, /* 3611 */
128'h00000000000000000000000000000000, /* 3612 */
128'h00000000000000000000000000000000, /* 3613 */
128'h00000000000000000000000000000000, /* 3614 */
128'h00000000000000000000000000000000, /* 3615 */
128'h00000000000000000000000000000000, /* 3616 */
128'h00000000000000000000000000000000, /* 3617 */
128'h00000000000000000000000000000000, /* 3618 */
128'h00000000000000000000000000000000, /* 3619 */
128'h00000000000000000000000000000000, /* 3620 */
128'h00000000000000000000000000000000, /* 3621 */
128'h00000000000000000000000000000000, /* 3622 */
128'h00000000000000000000000000000000, /* 3623 */
128'h00000000000000000000000000000000, /* 3624 */
128'h00000000000000000000000000000000, /* 3625 */
128'h00000000000000000000000000000000, /* 3626 */
128'h00000000000000000000000000000000, /* 3627 */
128'h00000000000000000000000000000000, /* 3628 */
128'h00000000000000000000000000000000, /* 3629 */
128'h00000000000000000000000000000000, /* 3630 */
128'h00000000000000000000000000000000, /* 3631 */
128'h00000000000000000000000000000000, /* 3632 */
128'h00000000000000000000000000000000, /* 3633 */
128'h00000000000000000000000000000000, /* 3634 */
128'h00000000000000000000000000000000, /* 3635 */
128'h00000000000000000000000000000000, /* 3636 */
128'h00000000000000000000000000000000, /* 3637 */
128'h00000000000000000000000000000000, /* 3638 */
128'h00000000000000000000000000000000, /* 3639 */
128'h00000000000000000000000000000000, /* 3640 */
128'h00000000000000000000000000000000, /* 3641 */
128'h00000000000000000000000000000000, /* 3642 */
128'h00000000000000000000000000000000, /* 3643 */
128'h00000000000000000000000000000000, /* 3644 */
128'h00000000000000000000000000000000, /* 3645 */
128'h00000000000000000000000000000000, /* 3646 */
128'h00000000000000000000000000000000, /* 3647 */
128'h00000000000000000000000000000000, /* 3648 */
128'h00000000000000000000000000000000, /* 3649 */
128'h00000000000000000000000000000000, /* 3650 */
128'h00000000000000000000000000000000, /* 3651 */
128'h00000000000000000000000000000000, /* 3652 */
128'h00000000000000000000000000000000, /* 3653 */
128'h00000000000000000000000000000000, /* 3654 */
128'h00000000000000000000000000000000, /* 3655 */
128'h00000000000000000000000000000000, /* 3656 */
128'h00000000000000000000000000000000, /* 3657 */
128'h00000000000000000000000000000000, /* 3658 */
128'h00000000000000000000000000000000, /* 3659 */
128'h00000000000000000000000000000000, /* 3660 */
128'h00000000000000000000000000000000, /* 3661 */
128'h00000000000000000000000000000000, /* 3662 */
128'h00000000000000000000000000000000, /* 3663 */
128'h00000000000000000000000000000000, /* 3664 */
128'h00000000000000000000000000000000, /* 3665 */
128'h00000000000000000000000000000000, /* 3666 */
128'h00000000000000000000000000000000, /* 3667 */
128'h00000000000000000000000000000000, /* 3668 */
128'h00000000000000000000000000000000, /* 3669 */
128'h00000000000000000000000000000000, /* 3670 */
128'h00000000000000000000000000000000, /* 3671 */
128'h00000000000000000000000000000000, /* 3672 */
128'h00000000000000000000000000000000, /* 3673 */
128'h00000000000000000000000000000000, /* 3674 */
128'h00000000000000000000000000000000, /* 3675 */
128'h00000000000000000000000000000000, /* 3676 */
128'h00000000000000000000000000000000, /* 3677 */
128'h00000000000000000000000000000000, /* 3678 */
128'h00000000000000000000000000000000, /* 3679 */
128'h00000000000000000000000000000000, /* 3680 */
128'h00000000000000000000000000000000, /* 3681 */
128'h00000000000000000000000000000000, /* 3682 */
128'h00000000000000000000000000000000, /* 3683 */
128'h00000000000000000000000000000000, /* 3684 */
128'h00000000000000000000000000000000, /* 3685 */
128'h00000000000000000000000000000000, /* 3686 */
128'h00000000000000000000000000000000, /* 3687 */
128'h00000000000000000000000000000000, /* 3688 */
128'h00000000000000000000000000000000, /* 3689 */
128'h00000000000000000000000000000000, /* 3690 */
128'h00000000000000000000000000000000, /* 3691 */
128'h00000000000000000000000000000000, /* 3692 */
128'h00000000000000000000000000000000, /* 3693 */
128'h00000000000000000000000000000000, /* 3694 */
128'h00000000000000000000000000000000, /* 3695 */
128'h00000000000000000000000000000000, /* 3696 */
128'h00000000000000000000000000000000, /* 3697 */
128'h00000000000000000000000000000000, /* 3698 */
128'h00000000000000000000000000000000, /* 3699 */
128'h00000000000000000000000000000000, /* 3700 */
128'h00000000000000000000000000000000, /* 3701 */
128'h00000000000000000000000000000000, /* 3702 */
128'h00000000000000000000000000000000, /* 3703 */
128'h00000000000000000000000000000000, /* 3704 */
128'h00000000000000000000000000000000, /* 3705 */
128'h00000000000000000000000000000000, /* 3706 */
128'h00000000000000000000000000000000, /* 3707 */
128'h00000000000000000000000000000000, /* 3708 */
128'h00000000000000000000000000000000, /* 3709 */
128'h00000000000000000000000000000000, /* 3710 */
128'h00000000000000000000000000000000, /* 3711 */
128'h00000000000000000000000000000000, /* 3712 */
128'h00000000000000000000000000000000, /* 3713 */
128'h00000000000000000000000000000000, /* 3714 */
128'h00000000000000000000000000000000, /* 3715 */
128'h00000000000000000000000000000000, /* 3716 */
128'h00000000000000000000000000000000, /* 3717 */
128'h00000000000000000000000000000000, /* 3718 */
128'h00000000000000000000000000000000, /* 3719 */
128'h00000000000000000000000000000000, /* 3720 */
128'h00000000000000000000000000000000, /* 3721 */
128'h00000000000000000000000000000000, /* 3722 */
128'h00000000000000000000000000000000, /* 3723 */
128'h00000000000000000000000000000000, /* 3724 */
128'h00000000000000000000000000000000, /* 3725 */
128'h00000000000000000000000000000000, /* 3726 */
128'h00000000000000000000000000000000, /* 3727 */
128'h00000000000000000000000000000000, /* 3728 */
128'h00000000000000000000000000000000, /* 3729 */
128'h00000000000000000000000000000000, /* 3730 */
128'h00000000000000000000000000000000, /* 3731 */
128'h00000000000000000000000000000000, /* 3732 */
128'h00000000000000000000000000000000, /* 3733 */
128'h00000000000000000000000000000000, /* 3734 */
128'h00000000000000000000000000000000, /* 3735 */
128'h00000000000000000000000000000000, /* 3736 */
128'h00000000000000000000000000000000, /* 3737 */
128'h00000000000000000000000000000000, /* 3738 */
128'h00000000000000000000000000000000, /* 3739 */
128'h00000000000000000000000000000000, /* 3740 */
128'h00000000000000000000000000000000, /* 3741 */
128'h00000000000000000000000000000000, /* 3742 */
128'h00000000000000000000000000000000, /* 3743 */
128'h00000000000000000000000000000000, /* 3744 */
128'h00000000000000000000000000000000, /* 3745 */
128'h00000000000000000000000000000000, /* 3746 */
128'h00000000000000000000000000000000, /* 3747 */
128'h00000000000000000000000000000000, /* 3748 */
128'h00000000000000000000000000000000, /* 3749 */
128'h00000000000000000000000000000000, /* 3750 */
128'h00000000000000000000000000000000, /* 3751 */
128'h00000000000000000000000000000000, /* 3752 */
128'h00000000000000000000000000000000, /* 3753 */
128'h00000000000000000000000000000000, /* 3754 */
128'h00000000000000000000000000000000, /* 3755 */
128'h00000000000000000000000000000000, /* 3756 */
128'h00000000000000000000000000000000, /* 3757 */
128'h00000000000000000000000000000000, /* 3758 */
128'h00000000000000000000000000000000, /* 3759 */
128'h00000000000000000000000000000000, /* 3760 */
128'h00000000000000000000000000000000, /* 3761 */
128'h00000000000000000000000000000000, /* 3762 */
128'h00000000000000000000000000000000, /* 3763 */
128'h00000000000000000000000000000000, /* 3764 */
128'h00000000000000000000000000000000, /* 3765 */
128'h00000000000000000000000000000000, /* 3766 */
128'h00000000000000000000000000000000, /* 3767 */
128'h00000000000000000000000000000000, /* 3768 */
128'h00000000000000000000000000000000, /* 3769 */
128'h00000000000000000000000000000000, /* 3770 */
128'h00000000000000000000000000000000, /* 3771 */
128'h00000000000000000000000000000000, /* 3772 */
128'h00000000000000000000000000000000, /* 3773 */
128'h00000000000000000000000000000000, /* 3774 */
128'h00000000000000000000000000000000, /* 3775 */
128'h00000000000000000000000000000000, /* 3776 */
128'h00000000000000000000000000000000, /* 3777 */
128'h00000000000000000000000000000000, /* 3778 */
128'h00000000000000000000000000000000, /* 3779 */
128'h00000000000000000000000000000000, /* 3780 */
128'h00000000000000000000000000000000, /* 3781 */
128'h00000000000000000000000000000000, /* 3782 */
128'h00000000000000000000000000000000, /* 3783 */
128'h00000000000000000000000000000000, /* 3784 */
128'h00000000000000000000000000000000, /* 3785 */
128'h00000000000000000000000000000000, /* 3786 */
128'h00000000000000000000000000000000, /* 3787 */
128'h00000000000000000000000000000000, /* 3788 */
128'h00000000000000000000000000000000, /* 3789 */
128'h00000000000000000000000000000000, /* 3790 */
128'h00000000000000000000000000000000, /* 3791 */
128'h00000000000000000000000000000000, /* 3792 */
128'h00000000000000000000000000000000, /* 3793 */
128'h00000000000000000000000000000000, /* 3794 */
128'h00000000000000000000000000000000, /* 3795 */
128'h00000000000000000000000000000000, /* 3796 */
128'h00000000000000000000000000000000, /* 3797 */
128'h00000000000000000000000000000000, /* 3798 */
128'h00000000000000000000000000000000, /* 3799 */
128'h00000000000000000000000000000000, /* 3800 */
128'h00000000000000000000000000000000, /* 3801 */
128'h00000000000000000000000000000000, /* 3802 */
128'h00000000000000000000000000000000, /* 3803 */
128'h00000000000000000000000000000000, /* 3804 */
128'h00000000000000000000000000000000, /* 3805 */
128'h00000000000000000000000000000000, /* 3806 */
128'h00000000000000000000000000000000, /* 3807 */
128'h00000000000000000000000000000000, /* 3808 */
128'h00000000000000000000000000000000, /* 3809 */
128'h00000000000000000000000000000000, /* 3810 */
128'h00000000000000000000000000000000, /* 3811 */
128'h00000000000000000000000000000000, /* 3812 */
128'h00000000000000000000000000000000, /* 3813 */
128'h00000000000000000000000000000000, /* 3814 */
128'h00000000000000000000000000000000, /* 3815 */
128'h00000000000000000000000000000000, /* 3816 */
128'h00000000000000000000000000000000, /* 3817 */
128'h00000000000000000000000000000000, /* 3818 */
128'h00000000000000000000000000000000, /* 3819 */
128'h00000000000000000000000000000000, /* 3820 */
128'h00000000000000000000000000000000, /* 3821 */
128'h00000000000000000000000000000000, /* 3822 */
128'h00000000000000000000000000000000, /* 3823 */
128'h00000000000000000000000000000000, /* 3824 */
128'h00000000000000000000000000000000, /* 3825 */
128'h00000000000000000000000000000000, /* 3826 */
128'h00000000000000000000000000000000, /* 3827 */
128'h00000000000000000000000000000000, /* 3828 */
128'h00000000000000000000000000000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00000000000000000000000000000000, /* 3840 */
128'h00000000000000000000000000000000, /* 3841 */
128'h00000000000000000000000000000000, /* 3842 */
128'h00000000000000000000000000000000, /* 3843 */
128'h00000000000000000000000000000000, /* 3844 */
128'h00000000000000000000000000000000, /* 3845 */
128'h00000000000000000000000000000000, /* 3846 */
128'h00000000000000000000000000000000, /* 3847 */
128'h00000000000000000000000000000000, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule

