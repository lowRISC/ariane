/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'h00008297ff81011b2000913711249263, /*    1 */
128'h0402829300008297000280e701a28293, /*    2 */
128'h00000597000280e71305051300000517, /*    3 */
128'h000046b7a19606130000c617fc458593, /*    4 */
128'h240e8e9b000f4eb7011696933ff6869b, /*    5 */
128'hfe0e9ae30085b703fffe8e930005b703, /*    6 */
128'h0006b703ff81011301b111130110011b, /*    7 */
128'h00e6b4230085b70300e6b0230005b703, /*    8 */
128'h00e6bc230185b70300e6b8230105b703, /*    9 */
128'h00000797fcc5cce30206869302058593, /*   10 */
128'h0007806740b787b300d787b301478793, /*   11 */
128'h0000c597305790730907879300000797, /*   12 */
128'h0005b023f94606130010d617a3458593, /*   13 */
128'h020585930005bc230005b8230005b423, /*   14 */
128'h00100913020004b73fe090effec5c6e3, /*   15 */
128'h4009091b02000937004484930124a023, /*   16 */
128'h008979133440297310500073ff24c6e3, /*   17 */
128'h00291913f1402973020004b7fe090ae3, /*   18 */
128'hfe091ee30004a9030009202300990933, /*   19 */
128'hff24c6e34009091b0200093700448493, /*   20 */
128'hffdff06f1050007334102373342022f3, /*   21 */
128'h6e61697241206d6f7266206f6c6c6548, /*   22 */
128'h61207469617720657361656c50202165, /*   23 */
128'h00000000000a2e2e2e746e656d6f6d20, /*   24 */
128'h00000000000000000000000000000000, /*   25 */
128'h00000000000000000000000000000000, /*   26 */
128'h00000000000000000000000000000000, /*   27 */
128'h00000000000000000000000000000000, /*   28 */
128'h00000000000000000000000000000000, /*   29 */
128'h00000000000000000000000000000000, /*   30 */
128'h00000000000000000000000000000000, /*   31 */
128'hd963454c0005cc635735c28587ae6914, /*   32 */
128'he21c97b6470102a787b30a00051300b7, /*   33 */
128'h853e85b200030563018533038082853a, /*   34 */
128'h738686930000b697b7edfda007138302, /*   35 */
128'h87930000c7976294820707130000c717, /*   36 */
128'h87b30280069302d787bb878d8f998167, /*   37 */
128'h47148082853a470100e7956397ba02d7, /*   38 */
128'hf0efe4061141b7f502870713fea68de3, /*   39 */
128'hbfe545018082014160a26108c509fbbf, /*   40 */
128'hf0efe852ec4ef04af426f822fc067139, /*   41 */
128'h0000ba17440144814985892acd31f9bf, /*   42 */
128'hc091553500f44d6300c927832c4a0a13, /*   43 */
128'h61216a4269e2790274a2744270e24501, /*   44 */
128'h67a2ed19f29ff0ef854a85a200308082, /*   45 */
128'h50ef8552000995632485cb990087c783, /*   46 */
128'h0513bf65240511c080ef498165224960, /*   47 */
128'hf2dff0efe42ef406f0227179b7c1fda0, /*   48 */
128'h842aee7ff0ef083065a2c105fda00413, /*   49 */
128'h00f7096300c547030ff007936562e911, /*   50 */
128'h547980826145740270a285220e2080ef, /*   51 */
128'hf0efec4ef04af426f822fc067139bfd5, /*   52 */
128'h0000a9970ff00913440184aacd01eebf, /*   53 */
128'h74a2744270e200f4496344dc44498993, /*   54 */
128'hf0ef852685a200308082612169e27902, /*   55 */
128'h85a20127896300c7c78367a2ed09e83f, /*   56 */
128'hb7d9240507c080ef65223f2050ef854e, /*   57 */
128'he8dff0ef892eec26f406e84af0227179, /*   58 */
128'he45ff0ef84aa85ca0030c11dfda00413, /*   59 */
128'h3e8505130000a517864a608ced01842a, /*   60 */
128'h740270a2852203e080ef65223b4050ef, /*   61 */
128'hf406ec26f022717980826145694264e2, /*   62 */
128'h85a6842ac11dfda00413e47ff0ef84ae, /*   63 */
128'hcf63445c37c050ef3c0505130000a517, /*   64 */
128'h5435004080ef3be505130000a51700f4, /*   65 */
128'h003085228082614564e2740270a28522, /*   66 */
128'h7d9070ef6522f565842adcfff0ef85a6, /*   67 */
128'h5479fcf71be30ff0079300c7c70367a2, /*   68 */
128'he50965a2de1ff0eff406e42e7179bfc1, /*   69 */
128'hf96dd97ff0ef08308082614570a24501, /*   70 */
128'he42eec064108842ae8221101bfc56562, /*   71 */
128'h852200030e6302053303c919db9ff0ef, /*   72 */
128'h60e2fda005138302610560e265a26442, /*   73 */
128'h0000b7977139bfdd4501808261056442, /*   74 */
128'h04130000b417f426f822639c4c478793, /*   75 */
128'h043b840d8c0559e484930000b4975a64, /*   76 */
128'h892afc06e852ec4ef04a0280079302f4, /*   77 */
128'h942602f404332fea0a130000aa1789ae, /*   78 */
128'h69e2790274a2744270e2450100849b63, /*   79 */
128'h278050ef855285ca6090808261216a42, /*   80 */
128'hbfc902848493c501685060ef854a608c, /*   81 */
128'hb7e16522f569cdbff0ef852685ce0030, /*   82 */
128'h84b68432e42efc06f04af426f8227139, /*   83 */
128'hcb5ff0ef083065a2c115cf7ff0ef893a, /*   84 */
128'h70e2978285a2615c862686ca6562e519, /*   85 */
128'hbfc5fda0051380826121790274a27442, /*   86 */
128'h84b68432e42efc06f04af426f8227139, /*   87 */
128'hc75ff0ef083065a2c115cb7ff0ef893a, /*   88 */
128'h70e2978285a2655c862686ca6562e519, /*   89 */
128'hbfc5fda0051380826121790274a27442, /*   90 */
128'hc7dff0ef84b2e42ef822fc06f4267139, /*   91 */
128'h701ce509c39ff0ef842a083065a2c105, /*   92 */
128'h8082612174a2744270e2978285a66562, /*   93 */
128'h2785c3190017f713419cbfcdfda00513, /*   94 */
128'hd71b8e5927a106220086571b419cc19c, /*   95 */
128'h0ff77713c19c0087d7138ed906a20086, /*   96 */
128'h122300d5112300c510238fd90087979b, /*   97 */
128'hf022f4067179419c80820005132300f5, /*   98 */
128'h419c00f510230457879b6785c19c27d1, /*   99 */
128'h0087979b0ff777130087d713c632842a, /*  100 */
128'hc4360509084c57fd460900f11a238fd9, /*  101 */
128'h0513016105934609773060ef00f11b23, /*  102 */
128'h00041323082c462147c1765060ef0044, /*  103 */
128'h00f404a347c5751060efec3e00840513, /*  104 */
128'h73b060ef00c4051300041523006c4611, /*  105 */
128'h0144069372f060ef01040513002c4611, /*  106 */
128'hfed79ce39f31ffe7d6030789470187a2, /*  107 */
128'h9fb94107d71b9fb9934117424107579b, /*  108 */
128'h80826145740270a200f41523fff7c793, /*  109 */
128'h97ba46a167856398338787930000b797, /*  110 */
128'hc7bb27850077e793fff6079b8007bc23, /*  111 */
128'h3823973e678500f547636805450102d7, /*  112 */
128'h010686bb0035169b0005b883808280c7, /*  113 */
128'he0221141bff105a125050116b02396ba, /*  114 */
128'hfa5ff0efe406450185aa86220005841b, /*  115 */
128'hec26f022717980820141640260a28522, /*  116 */
128'h67b060efe436f4064619051984b2842a, /*  117 */
128'h162347a166f060ef85b64619852266a2, /*  118 */
128'h614564e200e4859b70a27402852200f4, /*  119 */
128'h3a8130236785737dc5010113fadff06f, /*  120 */
128'h3931342338913c233a11342339213823, /*  121 */
128'h377134233761382337513c2339413023, /*  122 */
128'h3507879335a1382335913c2337813023, /*  123 */
128'hce042023d00007b7943e747d978a911a, /*  124 */
128'hd0040023f0040023e0040023ca040b23, /*  125 */
128'ha51785aa00e7ea63892a5800073797aa, /*  126 */
128'h00054703a00178f040ef002505130000, /*  127 */
128'h970a3507871374fd678526f711634789, /*  128 */
128'hcb848b13970a350787139abacd848a93, /*  129 */
128'h9c3a9b3a49818a368cb28baed0048c13, /*  130 */
128'hc7830015cd03013907b395ca0f098593, /*  131 */
128'h869b01a989bb058902a0071329890f07, /*  132 */
128'h24e78163471904f76b6326e78d630007, /*  133 */
128'hcc848513470d2ae78963470502f76263, /*  134 */
128'h40ef0f2505130000a51785b622e78963, /*  135 */
128'hfee794e3473d22e785634731b77d7070, /*  136 */
128'h953e866ae0048513978a350787936785, /*  137 */
128'h03600713b759e00d0023535060ef9d22, /*  138 */
128'h22e780630330071300f76e6322e78363, /*  139 */
128'haad94605cb648513fae798e303500713, /*  140 */
128'hf8e79ce30ff0071324e7856303800713, /*  141 */
128'h24e781630007859b747d471500614783, /*  142 */
128'h000ca7833ae79063470936e784634719, /*  143 */
128'h05134985978a350a87936a8516079263, /*  144 */
128'h60ef013ca023953e461101090593ce44, /*  145 */
128'h01490593ce840513978a350a87934b90, /*  146 */
128'hed8505130000a5174a3060ef953e4611, /*  147 */
128'h978a350a879363f040efde0254e25a52, /*  148 */
128'h429060ef854a55fd4619993ecf840913, /*  149 */
128'h879346f115231350079300f103a3478d, /*  150 */
128'h85a6460594becb740493c2a6978a350a, /*  151 */
128'h06a303200793451060efc0d246c10513, /*  152 */
128'h4a1195becf040593978a350a879346f1, /*  153 */
128'h079342d060ef4741072346f105134611, /*  154 */
128'hcf440593978a350a879346f109a30360, /*  155 */
128'h40b060ef47410a2347510513461195be, /*  156 */
128'h03a346f10ca347b1051385a6460557fd, /*  157 */
128'h0613102007933f1060ef47310d230001, /*  158 */
128'h079338b060efde3e37a1051345810f00, /*  159 */
128'h3961051385de4799464136f11d231010, /*  160 */
128'h13232637879377e13c3060ef36f10e23, /*  161 */
128'h350a879346f1142335378793679946f1, /*  162 */
128'h0440061304300693943ecec40413978a, /*  163 */
128'h85a2460156fdba1ff0ef3721051385a2, /*  164 */
128'h0e8885de86ca5672bd5ff0ef35e10513, /*  165 */
128'h3a0134033a813083911a6305cebff0ef, /*  166 */
128'h38013a03388139833901390339813483, /*  167 */
128'h36013c0336813b8337013b0337813a83, /*  168 */
128'h851380823b01011335013d0335813c83, /*  169 */
128'ha00d953e978a3507879367854611cd04, /*  170 */
128'h953e866af0048513978a350787936785, /*  171 */
128'h85564611b39df00d0023315060ef9d22, /*  172 */
128'h87936785bfdd855a4611bbb1307060ef, /*  173 */
128'h2eb060ef4611953ece048513978a3507, /*  174 */
128'h00f40123ce14478300f401a3ce044783, /*  175 */
128'h00f40023ce34478300f400a3ce244783, /*  176 */
128'h866ab759cc048513bb29cef42023401c, /*  177 */
128'h2783b311d00d00232b3060ef9d228562, /*  178 */
128'h0000a51700fa2023478510079d63000a, /*  179 */
128'h0e88010905934611441040efcec50513, /*  180 */
128'hcb840513978a350487936485287060ef, /*  181 */
128'h3531470326f060ef014905934611953e, /*  182 */
128'h0000a517350145833511460335214683, /*  183 */
128'h00a1468335015783401040efcbc50513, /*  184 */
128'h35215783fcf71e230000b71700914603, /*  185 */
128'h0000b717cbc505130000a51700814583, /*  186 */
128'h01b147033cd040ef00b14703fcf71323, /*  187 */
128'h0000a517018145830191460301a14683, /*  188 */
128'h01214683013147033b1040efcbc50513, /*  189 */
128'hcc0505130000a5170101458301114603, /*  190 */
128'h05130000a51755c201015783395040ef, /*  191 */
128'hb71701215783f6f713230000b717cce5, /*  192 */
128'h978a3504879336f040eff4f71e230000, /*  193 */
128'h40efcba505130000a51795bee0040593, /*  194 */
128'ha51795be978af0040593350487933570, /*  195 */
128'h0000a517bd2933f040efcb2505130000, /*  196 */
128'h93e3000a2783b531331040efcb450513, /*  197 */
128'hca8505130000a51700fa20234785e007, /*  198 */
128'h309040efcac505130000a517315040ef, /*  199 */
128'ha51795be978ad0040593350787936785, /*  200 */
128'hcb8505130000a517bf45cb2505130000, /*  201 */
128'he4a6e8a2ec86711d737db3c12e5040ef, /*  202 */
128'h0000a517911a89aaf456f852fc4ee0ca, /*  203 */
128'h8793747d2bd040efca026a85ccc50513, /*  204 */
128'h852655fd461994beff840493978a020a, /*  205 */
128'h0913439cd1c787930000b7970a5060ef, /*  206 */
128'h879312f11d2313500793c83e4a05fef4, /*  207 */
128'h014107a31a68460585ca993e978a020a, /*  208 */
128'h0f23479112f10ea3037007930c7060ef, /*  209 */
128'h461195beff040593978a020a879312f1, /*  210 */
128'h0513460585ca57fd0a3060ef13f10513, /*  211 */
128'h60ef000107a31541022314f101a31451, /*  212 */
128'h04a1051345810f0006130fc007930890, /*  213 */
128'h85ce04f1152310100793023060efca3e, /*  214 */
128'h05b060ef04f106230661051346414799, /*  215 */
128'h35378793679912f11b232637879377e1, /*  216 */
128'h85a2943e1451978a020a879312f11c23, /*  217 */
128'h83bff0ef044006130430069304210513, /*  218 */
128'h465286fff0ef460156fd02e1051385a2, /*  219 */
128'h60e6911a6305985ff0ef85ce86a61008, /*  220 */
128'h61257aa27a4279e2690664a664464501, /*  221 */
128'h1990406fbbc505130000a51785aa8082, /*  222 */
128'h7c913c237e8130237e11342381010113, /*  223 */
128'h05a1051384aa71597d3134237d213823, /*  224 */
128'h60efd602e83eec3ae442893689b2e046, /*  225 */
128'h6762747d97ba81078793101867857b80, /*  226 */
128'h0521051385a2864a86ba943e7fc40413, /*  227 */
128'h863e86c285a267c26822fa4ff0efd64e, /*  228 */
128'h85a6180856326882fd4ff0ef03e10513, /*  229 */
128'h340345017e81308361658e9ff0ef86c6, /*  230 */
128'h01137c8139837d0139037d8134837e01, /*  231 */
128'h480300554883e222e606716d80827f01, /*  232 */
128'h46030015468300254703003547830045, /*  233 */
128'h0000a517b0c585930000a597842a0005, /*  234 */
128'h842adedff0ef85220d1040efb0c50513, /*  235 */
128'h0000a517aec585930000a597860ac10d, /*  236 */
128'h6151641260b285220b1040efb1450513, /*  237 */
128'hab230000b797b2e505130000a5178082, /*  238 */
128'he4ceeca6f0a27159b7cd093040efc007, /*  239 */
128'hf486e86aec66f062f45ef85afc56e0d2, /*  240 */
128'hba974401ff05049389ae8a2ae46ee8ca, /*  241 */
128'h0b93b02b0b130000ab17802a8a930000, /*  242 */
128'h8c930000ac97b0ec0c130000ac170600, /*  243 */
128'h64e6740670a603344163fff58d1bafec, /*  244 */
128'h6ce27c027ba27b427ae26a0669a66946, /*  245 */
128'he7a9c42900f47793808261656da26d42, /*  246 */
128'hc583012487b34dc14901013040ef855a, /*  247 */
128'h856602fbe2630ff7f793fe05879b0007, /*  248 */
128'h05130000a517ffb912e309057f4040ef, /*  249 */
128'h8562a0317dc040ef85567e2040ef5d65, /*  250 */
128'h0000a5170104c583dbe5b7c57d4040ef, /*  251 */
128'hfffd4913028d1d637c0040efa8c50513, /*  252 */
128'h2d857aa040ef8556a02900f979134d81, /*  253 */
128'h079bff04791379e040ef855aff2dcce3, /*  254 */
128'h40ef57a505130000a51700f45b630009, /*  255 */
128'h0007c583012a07b3b781048524057860, /*  256 */
128'h40ef856600fbe7630ff7f793fe05879b, /*  257 */
128'h7179bfdd75c040ef8562b7e909057660, /*  258 */
128'h893289ae84b6f022f406e44ee84aec26, /*  259 */
128'h86930000a697c5092a8686930000a697, /*  260 */
128'h06130000a617b167071300009717a066, /*  261 */
128'h00098f63842a6de040ef854a85a69fe6, /*  262 */
128'h06130000a61786ce40a485bb00955d63, /*  263 */
128'h4463ffe4879b9c296c0040ef954a9e66, /*  264 */
128'h85930000a59700890533ffd4841b00f4, /*  265 */
128'h694264e2854a740270a2278060ef9b65, /*  266 */
128'hf73ff06f4581862e86b28082614569a2, /*  267 */
128'hfebff0efed8645050c800613002c7115, /*  268 */
128'h60ee6aa040ef99e505130000a517002c, /*  269 */
128'h862e9ff787133b9ad7b78082612d4501, /*  270 */
128'h04a7676323f78713000f47b704a76963, /*  271 */
128'hb7173e80079346890ca7f7633e700793, /*  272 */
128'h00074903e04a97361101902707130000, /*  273 */
128'h64a260e2644202091663e426e822ec06, /*  274 */
128'h406f6105944505130000a51785aa6902, /*  275 */
128'h240787934685b7d9a007879346816460, /*  276 */
128'h3e800793c02102f555b302f57433bf7d, /*  277 */
128'h0713c70502f4773347a90287e6634729, /*  278 */
128'h743302f457b306400713028774630630, /*  279 */
128'h5433a039943e001444130324341302e4, /*  280 */
128'h05130000a517f86102f45433bfc102e4, /*  281 */
128'h0000a51785a2c8015e0040ef84b28ee5, /*  282 */
128'h85ca862660e264425d0040ef8e450513, /*  283 */
128'h406f61058d4505130000a517690264a2, /*  284 */
128'h862eb78d8a4505130000a51785aa5b60, /*  285 */
128'h55b303c6871b02f886bb481958d94781, /*  286 */
128'h810808130000b81793811782cd8500e5, /*  287 */
128'he04ae822ec060007c483e42697c21101, /*  288 */
128'h0000a51785aa690264a260e26442e495, /*  289 */
128'hfb079de3278555e0406f610588450513, /*  290 */
128'h97b357fdb7f586e505130000a51785aa, /*  291 */
128'h053347a9c10d44018d7dfff7c79300e7, /*  292 */
128'h942a47a500d41433440503b6869b02f5, /*  293 */
128'h0000a517058514590087f46300e45433, /*  294 */
128'ha51785a2c80150e040ef893281c50513, /*  295 */
128'h864a60e264424fe040ef812505130000, /*  296 */
128'h610581a505130000a51764a2690285a6, /*  297 */
128'hf1a202c7073b8cbaed6671514e40406f, /*  298 */
128'hf95afd56e1d2eda6f586e96ae5cee9ca, /*  299 */
128'h8d3289ae892a04000793e56ef162f55e, /*  300 */
128'h956302ccdcbb04000c9300e7f6638436, /*  301 */
128'h020d1a13001d179b03acdcbb4cc1000c, /*  302 */
128'h9b1703810a93020a5a130017849be03e, /*  303 */
128'h8c1772ab8b9300009b977c2b0b130000, /*  304 */
128'h64ee740e70ae4501e00d2f2c0c130000, /*  305 */
128'h6cea7c0a7baa7b4a7aea6a0e69ae694e, /*  306 */
128'h05130000951785ca8082616d6daa6d4a, /*  307 */
128'h8d9b008cf46300040d9b442040ef77e5, /*  308 */
128'h0007061b430948a14811470186ce000c, /*  309 */
128'h99ba034707339301020d971305b66c63, /*  310 */
128'h861b02e00813875603bd06bb0d9de663, /*  311 */
128'h85d6963e011c0ac5ed63415705bb0006, /*  312 */
128'h40effa060c23e4367385051300009517, /*  313 */
128'h60ef99369281168241b4043b66a23e60, /*  314 */
128'h15934290030d1b63b795557dd1357c70, /*  315 */
128'h855a658292011602c190260195d60027, /*  316 */
128'h66a23aa040efe436e83aec42f046f41a, /*  317 */
128'h1863bf8568627882070596d273226742, /*  318 */
128'h1c63bfc1e19095d6003715936290011d, /*  319 */
128'h9241164295d6001715930006d603006d, /*  320 */
128'h761300ea85b30006c603bf6500c59023, /*  321 */
128'h7f3060efe43a855eb75d00c580230ff6, /*  322 */
128'hbfdd4701bf1d3cfdfe976ae327056722, /*  323 */
128'h097575130005450300bc053300074583, /*  324 */
128'h00230005d4634185d59b0185959bc519, /*  325 */
128'hf4634501918187aa1582bf3907050107, /*  326 */
128'h04000793bfd58f8d25058082e21c00b7, /*  327 */
128'h57f70713464c47370005668312b7f463, /*  328 */
128'h10e6976347090045468310e69c634789, /*  329 */
128'hf0a202f7073371590380079303855703, /*  330 */
128'he4cee8caeca6f48602059a93fc567100, /*  331 */
128'hda93e46ee86aec66f062f45ef85ae0d2, /*  332 */
128'h942a84aa892e06eae663478d9722020a, /*  333 */
128'h00009c175ecb8b9300009b974b054a01, /*  334 */
128'h0384d78360cc8c9300009c9762cc0c13, /*  335 */
128'h741c09679b63401ca835478100fa6463, /*  336 */
128'h8d630204398326e040ef855e85d2cbc1, /*  337 */
128'hfa6395ce00b48db301843d03640c0409, /*  338 */
128'h248040ef5ac5051300009517864a02ba, /*  339 */
128'h7ae26a0669a6694664e6740670a6478d, /*  340 */
128'h6165853e6da26d426ce27c027ba27b42, /*  341 */
128'h864e21a040ef856686ce85ea866e8082, /*  342 */
128'hf163701c02843983062060ef856a85ee, /*  343 */
128'h85ea9d3e864e40f989b301843d030337, /*  344 */
128'h7e9050ef856a4581864e1f2040ef8562, /*  345 */
128'h45058082853e4785bf99038404132a05, /*  346 */
128'h07130000a7178082400005378082057e, /*  347 */
128'h95360017869300756513157d631c56e7, /*  348 */
128'h8082953e057e450597aa20000537e308, /*  349 */
128'h08a74463862a0ce50763820787136785, /*  350 */
128'h06e60b6354c505130000951780878713, /*  351 */
128'h52850513000095178006079b04c74963, /*  352 */
128'h5a8505130000951787f787936785c3ad, /*  353 */
128'h95979e3d11417c07879b77fd04c7c963, /*  354 */
128'he4064d2505130000a51759a585930000, /*  355 */
128'h01414c2505130000a51760a2120040ef, /*  356 */
128'h0a634fa5051300009517810787138082, /*  357 */
128'h12e34fa50513000095178187879300e6, /*  358 */
128'h5185051300009517830787138082faf6, /*  359 */
128'h000095178287879300c74963fee609e3, /*  360 */
128'h05130000951783878713bfe94f450513, /*  361 */
128'h05130000951784078793fce608e35065, /*  362 */
128'h717980824bc5051300009517bf755065, /*  363 */
128'h4463440184ae892af406e84aec26f022, /*  364 */
128'h01045513942a90411442010455130290, /*  365 */
128'h694264e21542fff54513740270a29522, /*  366 */
128'h6db050ef0068460985ca808261459141, /*  367 */
128'h00d1478300f107a334f9090900c14783, /*  368 */
128'h6785715dbf55943e00e1578300f10723, /*  369 */
128'h842e80678793f44ef84afc26e486e0a2, /*  370 */
128'h079b0af50e636dd7879367a13cf50563, /*  371 */
128'h50ef4611082884b205e944079a638005, /*  372 */
128'h05130000a517461985ca006409136890, /*  373 */
128'h896302e0079301744583675050ef3c65, /*  374 */
128'h04b7e5631cf5826347b108b7e76332f5, /*  375 */
128'h10f58463478502b7e3631af583634791, /*  376 */
128'h951702f5836344650513000095174789, /*  377 */
128'h82634799a41d7df030ef5e2505130000, /*  378 */
128'hfef591e344c505130000951747a118f5, /*  379 */
128'h00b7ed632cf5826347f5a4317c5030ef, /*  380 */
128'h468505130000951747d916f58a6347c5, /*  381 */
128'h07932af5866302100793bf6dfef580e3, /*  382 */
128'hb7c94825051300009517faf596e30290, /*  383 */
128'h0330079304b7e2632cf5826306200793, /*  384 */
128'h28f5876302f0079300b7ef632af58263, /*  385 */
128'hf8f58ae3484505130000951703200793, /*  386 */
128'h951705e0079328f5846305c00793b7bd, /*  387 */
128'h08400793bf91f6f58de349a505130000, /*  388 */
128'h26f58b630670079300b7ef6328f58663, /*  389 */
128'hf4f58ae34ac505130000951706c00793, /*  390 */
128'h89630ff0079326f5886308900793b73d, /*  391 */
128'h051300009517f0f59ce30880079326f5, /*  392 */
128'h2d87d7830000a79701e45703b73d4b65, /*  393 */
128'h0204570312f714632d0989930000a997, /*  394 */
128'h85ca461910f71c632c27d7830000a797, /*  395 */
128'h290585930000a5974619515050ef8522, /*  396 */
128'h12230204012301a45783505050ef854a, /*  397 */
128'h0513fde4859b01c4578300f41f230204, /*  398 */
128'hd78300f41d230009d78302f410230224, /*  399 */
128'h812100a10ea3db9ff0ef00f41e230029, /*  400 */
128'h85a202f41223862601c1578300a10e23, /*  401 */
128'h2b85051300009517a06ddbffe0ef4501, /*  402 */
128'h00009517b5592c65051300009517bd41, /*  403 */
128'h0ea30264470302444783bdb52d450513, /*  404 */
128'h0ea301c1178300f10e230254478300f1, /*  405 */
128'h0224470300e10e2327810274470300e1, /*  406 */
128'h00e10e230234470300e10ea301c11903, /*  407 */
128'h0000a79704e79b6301c1568304500713, /*  408 */
128'h188585930000a597461947e21ad79823, /*  409 */
128'h18f728230000a717190505130000a517, /*  410 */
128'h87930000a79766a24762425050efe436, /*  411 */
128'h4ca060ef450102a40593ff89061b1667, /*  412 */
128'h07138082616179a2794274e2640660a6, /*  413 */
128'h14f728230000a71747e204e694630430, /*  414 */
128'h0000a797c799439c154787930000a797, /*  415 */
128'h138686930000a697f7e9439c14478793, /*  416 */
128'h138585930000a597134606130000a617, /*  417 */
128'h98634d200713b765d61fe0ef02a40513, /*  418 */
128'h85a654b030ef1ee505130000951702e7, /*  419 */
128'h30ef1ea5051300009517cb6ff0ef8522, /*  420 */
128'h0713bf95ca0ff0ef02a4051385ca5370, /*  421 */
128'h01e317fd67c101e45703f6e787e35fe0, /*  422 */
128'h0000a5974611f4f70de302045703f6f7, /*  423 */
128'h00009517b799351050ef08680f458593, /*  424 */
128'hb30d1ca5051300009517b3351c450513, /*  425 */
128'h051300009517bb211e05051300009517, /*  426 */
128'h9517b3112045051300009517b3391ee5, /*  427 */
128'h2285051300009517b9ed20a505130000, /*  428 */
128'h00009517b1dd2365051300009517b9c5, /*  429 */
128'hb9c92725051300009517b9f124c50513, /*  430 */
128'ha7970265d703b1e12805051300009517, /*  431 */
128'h11e306a484930000a4970727d7830000, /*  432 */
128'h19e305c7d7830000a7970285d703ecf7, /*  433 */
128'h9a23016589930205891320000793eaf7, /*  434 */
128'ha597461929f050ef854a85ce461900f5, /*  435 */
128'ha597461928f050ef854e01a585930000, /*  436 */
128'h461927d050ef0064051300a585930000, /*  437 */
128'h02a0061301c45783273050ef852285ca, /*  438 */
128'h0004d78302f4142301e4578302f41323, /*  439 */
128'h6080079300f41f230024d78300f41e23, /*  440 */
128'h208505130000951785aab36900f41623, /*  441 */
128'h8307b603300017b7bba546013e5030ef, /*  442 */
128'h171b00f674132601608130239f010113, /*  443 */
128'h05379f2d8406871b0387759366850034, /*  444 */
128'h34235e913c23630c8387b783972a3000, /*  445 */
128'h696335b95f200813ffc5849b25816011, /*  446 */
128'hfff7c79300c5963b101005938a1d08b8, /*  447 */
128'h4390f42787930000a797cfb527818ff1, /*  448 */
128'h9ebd8006869b7007f7930084179bea25, /*  449 */
128'h0106969b00d100a3872646d496aa068e, /*  450 */
128'h0001550300d100230086d69b0106d69b, /*  451 */
128'h02d51a63806686936685c6918005069b, /*  452 */
128'h46a1007767139fad377d8005859b6585, /*  453 */
128'h08378f95868a83f502d7473b17822705, /*  454 */
128'haa1ff0ef862602e6446397c285b63000, /*  455 */
128'h3403608130838287b823300017b70405, /*  456 */
128'h88338082610101135f81348385266001, /*  457 */
128'hb7e1ff06bc2306a126050008380300d7, /*  458 */
128'h2401ec06e42643c0e8220c2007b71101, /*  459 */
128'hc163033716938304b703300014b74781, /*  460 */
128'h2a9030ef0e45051300009517e7990206, /*  461 */
128'h8082610564a2644260e2c3c00c2007b7, /*  462 */
128'h8432ec26f0227179bfc14785eb9ff0ef, /*  463 */
128'hf4060068e6c585930000a597461184ae, /*  464 */
128'h0007a803e24787930000a7970c7050ef, /*  465 */
128'ha717e0a888930000a89785a6862247b2, /*  466 */
128'h05130000a51704500693e0e757030000, /*  467 */
128'h614564e2740270a285228aeff0efe165, /*  468 */
128'h8082914115428d5d05220085579b8082, /*  469 */
128'hf00686938fd966c10185579b0185171b, /*  470 */
128'h00ff07370085151b8fd98f750085571b, /*  471 */
128'h051300009517715d808225018d5d8d79, /*  472 */
128'hec56f052f44ef84afc26e0a2e4860465, /*  473 */
128'h47e1da0785230000a7971e3030efe85a, /*  474 */
128'h0000a71703e00793daf700a30000a717, /*  475 */
128'h578dd8f706a30000a7174789d8f70b23, /*  476 */
128'ha59707f007934611d8f702230000a717, /*  477 */
128'hd68404130000a4170028d74585930000, /*  478 */
128'h85a246097de050efd6f702a30000a717, /*  479 */
128'h89930000a997448145227d4050ef0068, /*  480 */
128'hf00606130100063746b2f4fff0efd2e9, /*  481 */
128'h15028f558f710ff6f69382a10086971b, /*  482 */
128'hb423934180a7b02317429101300017b7, /*  483 */
128'h0513000095178087b7038007b70380e7, /*  484 */
128'h8087b5838007b60382e7b4234721f965, /*  485 */
128'h91c115c2cdca0a130000aa1700800737, /*  486 */
128'h47030000a71710f030ef80e7b4238f4d, /*  487 */
128'h48030000a817cd27c7830000a797cd97, /*  488 */
128'h46030000a617cc06c6830000a697ccb8, /*  489 */
128'h051300009517cae5c5830000a597cb76, /*  490 */
128'h00989b376a89000447830d3030eff465, /*  491 */
128'h3000193700144783c8f70c230000a717, /*  492 */
128'h0000a71700244783c8f704a30000a717, /*  493 */
128'hc6f709a30000a71700344783c6f70f23, /*  494 */
128'h00544783c6f704230000a71700444783, /*  495 */
128'hc2079a230000a797c4f70ea30000a717, /*  496 */
128'hc207a8230000a797c207a4230000a797, /*  497 */
128'hc007ac230000a797c207a2230000a797, /*  498 */
128'h0493f4bfe0ef8522e78d0009a783e4a9, /*  499 */
128'h3783020745630337971383093783680b, /*  500 */
128'hbfc5c4fff0effc075de3033797138309, /*  501 */
128'h8493781050ef4501dff154fd000a2783, /*  502 */
128'h17b7b7d914fdb7e9c35ff0efbfc1710a, /*  503 */
128'he40616fd1141ff8006b78087b7033000, /*  504 */
128'h82e7b823f0070713670580e7b4238f75, /*  505 */
128'h7d8030efe7c50513000095178307b583, /*  506 */
128'h300027f37cc030efe985051300009517, /*  507 */
128'h07fe4785300790738fd9880707136709, /*  508 */
128'h7a8030efe94505130000951734179073, /*  509 */
128'h47838082014160a2302000730000100f, /*  510 */
128'h4503002547838f5d07a2000547030015, /*  511 */
128'h57fd808225018d5d05628fd907c20035, /*  512 */
128'h058505050005c703808200f61363367d, /*  513 */
128'h808200f61363367d57fdb7f5fee50fa3, /*  514 */
128'hec06e8221101495cbfcd050500b50023, /*  515 */
128'h478101853903cfa500958413e04ae426, /*  516 */
128'h462d02e0031348a5481586ca02000513, /*  517 */
128'h07130107146300a70e6327850006c703, /*  518 */
128'h00e40023040500640023011795630e50, /*  519 */
128'h01c9051300b94783fcc79ee306850405, /*  520 */
128'h01994783c088f59ff0ef00f5842384ae, /*  521 */
128'h478300f492238fd90087979b01894703, /*  522 */
128'h00f493238fd90087979b016947030179, /*  523 */
128'h80826105690264a2644260e200040023, /*  524 */
128'h468303a0061302000593cf99873e611c, /*  525 */
128'h06630017869300c6986302d5fc630007, /*  526 */
128'h46050007c683b7dd0705a00d577d00d7, /*  527 */
128'h078900b666630ff6f593fd06869b577d, /*  528 */
128'h47030000a7178082853ae11c0006871b, /*  529 */
128'hc70d0007c703cb85611cc915bfd5a6e7, /*  530 */
128'he406114102e69063008557030067d683, /*  531 */
128'hc3914501001577932c8060ef0017c503, /*  532 */
128'h01b5c783808245258082014160a24525, /*  533 */
128'h0007079b8f5d0087979b468d01a5c703, /*  534 */
128'h0087979b0145c6830155c78300d51d63, /*  535 */
128'h71798082853e27818fd90107979b8fd5, /*  536 */
128'h0993e052e84af4065904e44eec26f022, /*  537 */
128'h60ef85ce8626468500154503842a0345, /*  538 */
128'h87bb000402234c58505ce13125012560, /*  539 */
128'h694264e2740270a2450100e7eb6340f4, /*  540 */
128'h74e34a0500344903808261456a0269a2, /*  541 */
128'h85ce86269cbd4685001445034c5cff2a, /*  542 */
128'h00454783b7f94505b7e5397d214060ef, /*  543 */
128'he8221101591c80824501f8dff06fc399, /*  544 */
128'h892e84aa02b787634401e04ae426ec06, /*  545 */
128'h46850014c503ec190005041bfddff0ef, /*  546 */
128'h4405c119250119c060ef03448593864a, /*  547 */
128'h690264a2644260e285220324a823597d, /*  548 */
128'h57fde04ae426ec06e822110180826105, /*  549 */
128'he52d2501fa3ff0ef842ad91c00050223, /*  550 */
128'h8fd90087979b45092324470323344783, /*  551 */
128'h1f63a55707134107d79b776d0107979b, /*  552 */
128'h05370005079bd59ff0ef06a4051302f7, /*  553 */
128'hf7b31465049300544537fff509130100, /*  554 */
128'hd33ff0ef0864051300978c6345010127, /*  555 */
128'h644260e200a035338d05012575332501, /*  556 */
128'hf84a715dbfcd450d80826105690264a2, /*  557 */
128'h3023e85aec56f052fc26e0a2e486f44e, /*  558 */
128'h4e6347addd9ff0ef8932852e89aa0005, /*  559 */
128'h97ba872787930000a797003517130205, /*  560 */
128'h000447830089b023c01547b184aa6380, /*  561 */
128'he38d001577930e6060ef00144503cb85, /*  562 */
128'h74e2640660a647a9c111891100090563, /*  563 */
128'h80826161853e6b426ae27a0279a27942, /*  564 */
128'h7f9050ef00a400a3000400230ff4f513, /*  565 */
128'hf569891100090463fb71478d00157713, /*  566 */
128'h848a04f51a634785ee1ff0ef85224581, /*  567 */
128'h4501ffc9478389a623a40a131fa40913, /*  568 */
128'h094100a9a0232501c5bff0ef854ac789, /*  569 */
128'h45090004aa8301048913ff2a14e30991, /*  570 */
128'h0491c10de9dff0ef852285d6000a8763, /*  571 */
128'h470db7bd00e519634785470dfe9915e3, /*  572 */
128'h4783bfb947b5c1194a81f6e504e34785, /*  573 */
128'h0107979b8fd90087979b03f447030404, /*  574 */
128'h04b44983fef711e3200007134107d79b, /*  575 */
128'h1a09866300f9e9b30089999b04a44783, /*  576 */
128'hfff9079b470501342e23044449032981, /*  577 */
128'h04144b03faf769e30ff7f793012401a3, /*  578 */
128'h00fb77b3fffb079bfa0b03e301640123, /*  579 */
128'h6a33008a1a1b0454478304644a03ffc9, /*  580 */
128'h04844503f3c100fa77930144142300fa, /*  581 */
128'h478314050e638d450085151b04744483, /*  582 */
128'hdfb18fd90087979b2501042447030434, /*  583 */
128'h00d7063b9f3d004a571b2781033906bb, /*  584 */
128'h84ae0364d5bb40c504bbf4c564e38732, /*  585 */
128'h0905165500b93933664119556905dd8d, /*  586 */
128'h015787bb248900ea873b490d00b67363, /*  587 */
128'h10e91263470dd05c03542023cc04d458, /*  588 */
128'h949bd408b17ff0ef06040513f00a15e3, /*  589 */
128'hee99e7e324810094d49b1ff4849b0024, /*  590 */
128'h478d00f402a3f8000793c45cc81c57fd, /*  591 */
128'h0087979b064447030654478308f91963, /*  592 */
128'h06f71b6347054107d79b0107979b8fd9, /*  593 */
128'h4783e13d2501ce5ff0ef8522001a859b, /*  594 */
128'h8fd90087979b000402a3232447032334, /*  595 */
128'h1263a55707134107d79b776d0107979b, /*  596 */
128'h2501416157b7a99ff0ef0344051304f7, /*  597 */
128'ha83ff0ef2184051302f5176325278793, /*  598 */
128'h051300f51c63272787932501614177b7, /*  599 */
128'ha63ff0ef22040513c808a6dff0ef21c4, /*  600 */
128'h93c117c227855f87d78300009797c448, /*  601 */
128'h0124002300f413235ef7152300009717, /*  602 */
128'ha33ff0ef05840513b351478100042a23, /*  603 */
128'hb545a25ff0ef05440513b5b90005099b, /*  604 */
128'h949b00f915634789d41c9fb5e00a05e3, /*  605 */
128'h0017d79b8885029787bb478db7010014, /*  606 */
128'hf0ef842ae426ec06e8221101bdc59cbd, /*  607 */
128'h0cf71063478d00044703ed692501bfff, /*  608 */
128'h0613034404930af71b63478500544703, /*  609 */
128'h092305500793a01ff0ef852645812000, /*  610 */
128'h0a230520079322f409a3faa0079322f4, /*  611 */
128'h0da302f40b230610079302f40aa302f4, /*  612 */
128'h20e40d2302e40ba304100713481c20f4, /*  613 */
128'h20f40e230087571b0107571b0107971b, /*  614 */
128'h20f40fa30187d79b0107d71b20e40ea3, /*  615 */
128'h0107571b0107971b501020e40f23445c, /*  616 */
128'h22f4002307200693001445030087571b, /*  617 */
128'h0c230187d79b0107d71b260522e400a3, /*  618 */
128'hd81022f401a322e4012320d40ca320d4, /*  619 */
128'h00144503000402a3541050ef85a64685, /*  620 */
128'h60e200a035332501535050ef45814601, /*  621 */
128'h37f9ffe5869b4d1c8082610564a26442, /*  622 */
128'h9d2d02d585bb55480025458300f6f963, /*  623 */
128'h71794d180eb7f7634785808245018082, /*  624 */
128'h02e5f963892ae44eec26f022f406e84a, /*  625 */
128'h0e63468d06d70c63842e468900054703, /*  626 */
128'hd59b9cad515c0015d49b00f71e6308d7, /*  627 */
128'h70a257fdc9112501ac7ff0ef9dbd0094, /*  628 */
128'h278380826145853e69a2694264e27402, /*  629 */
128'h94ca1ff4f4930099d59b0014899b0249, /*  630 */
128'hf5792501a93ff0ef0344c483854a9dbd, /*  631 */
128'h0087979b880503494783994e1ff9f993, /*  632 */
128'hbf458fe9157d6505bf658391c0198fc5, /*  633 */
128'hfd592501a63ff0ef9dbd0085d59b515c, /*  634 */
128'h45030359478399221fe474130014141b, /*  635 */
128'h0075d59b515cb7598fc90087979b0349, /*  636 */
128'h75130024151bf9352501a39ff0ef9dbd, /*  637 */
128'h100007b7807ff0ef954a034505131fc5, /*  638 */
128'hf82271398082853e4785b76517fd2501, /*  639 */
128'h1523e456e852ec4ef426fc06f04a4540, /*  640 */
128'h744270e2450900f41c63892a478500b5, /*  641 */
128'h611c808261216aa26a4269e2790274a2, /*  642 */
128'h470d0007c683e02184aefee474e34f98, /*  643 */
128'hfce4f7e30087d703eb15579800e69463, /*  644 */
128'h37839d3d0044d79bd171008928235788, /*  645 */
128'h00a92a2394be03478793049688bd0009, /*  646 */
128'h843a0027c9838722b75d450100993c23, /*  647 */
128'h0134f66385a2000935034a8509925a7d, /*  648 */
128'h0005041be6fff0efbf752501e59ff0ef, /*  649 */
128'h76e34f9c00093783f68afbe301440c63, /*  650 */
128'h00a55583b78d4505bfc1413484bbf6f4, /*  651 */
128'h049bf33ff0ef842aec06e426e8221101, /*  652 */
128'h0005049b933ff0ef6008484ce4950005, /*  653 */
128'h6c1cf3cff0ef4581020006136c08ec99, /*  654 */
128'h60e200e782234705601c00e780235715, /*  655 */
128'hfc06e85271398082610564a285266442, /*  656 */
128'h16ba75634a05e456ec4ef04af426f822, /*  657 */
128'h4709000547830af5f063498984aa4d1c, /*  658 */
128'h94630ee78863470d0ae78f63842e8932, /*  659 */
128'h009a559b00ba0a3b515c0015da1b1547, /*  660 */
128'h8805060996630005099b8b9ff0ef9dbd, /*  661 */
128'h87b3cc191ffa7a130ff97793001a0a9b, /*  662 */
128'h179b00f7f71316c166850347c7830144, /*  663 */
128'h02fa0a239a260ff7f7938fd98ff50049, /*  664 */
128'h9dbd8526009ad59b50dc00f482234785, /*  665 */
128'h1ffafa9300099f630005099b86bff0ef, /*  666 */
128'h032a8a239aa60ff979130049591bc40d, /*  667 */
128'h790274a2854e744270e200f482234785, /*  668 */
128'hc783015487b3808261216aa26a4269e2, /*  669 */
128'h0127e9339bc100f979130089591b0347, /*  670 */
128'h099b811ff0ef9dbd0085d59b515cb7e9, /*  671 */
128'h94261fe474130014141bfc0992e30005, /*  672 */
128'h0089591b0109591b0109191b03240a23, /*  673 */
128'h0075d59b515cbf790144822303240aa3, /*  674 */
128'h141bf80996e30005099bfd8ff0ef9dbd, /*  675 */
128'hf0ef85569aa603440a931fc474130024, /*  676 */
128'h179b012569338d71f00006372501da0f, /*  677 */
128'h0087d79b03240a230107d79b94260109, /*  678 */
128'h00fa81230189591b0109579b00fa80a3, /*  679 */
128'hec4ef4267139bf3d4989b745012a81a3, /*  680 */
128'he19d89ae84aae456e852f04af822fc06, /*  681 */
128'h844a04f977634d1c04090a6300c52903, /*  682 */
128'h052a606304f4636324054c9c5afd4a05, /*  683 */
128'hf86347850005041bc43ff0efa8214401, /*  684 */
128'h744270e28522547d00f41d6357fd0887, /*  685 */
128'h4c9c808261216aa26a4269e2790274a2, /*  686 */
128'h85a24409bf554905b7d5faf47ee3894e, /*  687 */
128'h0863fd5507e3c9012501c05ff0ef8526, /*  688 */
128'h85a2167d10000637b76dfb2411e30545, /*  689 */
128'h489c02099063e9052501de9ff0ef8526, /*  690 */
128'h0054c783c89c37fdfae783e3577dc4c0, /*  691 */
128'h852685ce8622bf4900f482a30017e793, /*  692 */
128'h4405f6f50fe34785dd612501dbbff0ef, /*  693 */
128'h2905f822fc0600a55903f04a7139bfad, /*  694 */
128'heb9993c1e456e852ec4ef42603091793, /*  695 */
128'h6aa26a4269e2790274a2744270e24511, /*  696 */
128'h842a8a2e00f97993d7ed495c80826121, /*  697 */
128'h5783e18dc85c61082785480c00099d63, /*  698 */
128'h15230996601cfcf775e30009071b0085, /*  699 */
128'h4783bf5d4501ec1c97ce034787930124, /*  700 */
128'hfc0a9fe30157fab337fd00495a9b0025, /*  701 */
128'h45090097e46347850005049bb27ff0ef, /*  702 */
128'h4d1c6008b761450500f4946357fdbf49, /*  703 */
128'h049be81ff0ef480cf60a0ee306f4e063, /*  704 */
128'h8de357fdfcf48be34785d4bd451d0005, /*  705 */
128'h06136008f5792501dd8ff0ef6008fcf4, /*  706 */
128'h00043a03beeff0ef0345051345812000, /*  707 */
128'h60084a0502aa2823aa5ff0ef855285a6, /*  708 */
128'hd91c415787bb591c00faed6300254783, /*  709 */
128'h0223b7b9c848a83ff0ef85a6c8046008, /*  710 */
128'h5b1c2a856018f1412501d1cff0ef0145, /*  711 */
128'hf04afc06f426f8227139b7e9db1c2785, /*  712 */
128'h02f007130005c783e05ae456e852ec4e, /*  713 */
128'h0ce7906305c0071300e78663842e84aa, /*  714 */
128'h0ae7fc6347fd000447030004a6230405, /*  715 */
128'h47834b2102e0099305c00a9302f00a13, /*  716 */
128'h462d0204b9030d5780630d4782630004, /*  717 */
128'h926300044783b40ff0ef854a02000593, /*  718 */
128'h07930b37906300144783013900230d37, /*  719 */
128'h470d1b378e630024478300f900a302e0, /*  720 */
128'h458100f905a302000793943a09479763, /*  721 */
128'h608848cc100510632501adbff0ef8526, /*  722 */
128'hc7e5000747836c98e96d2501cdaff0ef, /*  723 */
128'h8d6300b78593709cef918ba100b74783, /*  724 */
128'h08e3fff7c683fff74603078507050cb7, /*  725 */
128'h4bdc611cbf75dfdff0ef85264581fed6, /*  726 */
128'hbc232501a85ff0ef85264581b791c55c, /*  727 */
128'h6aa26a4269e2790274a2744270e20004, /*  728 */
128'h8be3bf954709bf1d0405808261216b02, /*  729 */
128'h02400793943a12f6e06302000693f757, /*  730 */
128'h486502000313478145a147014681b7ad, /*  731 */
128'h9101020695130027e793a8dd0505a0d1, /*  732 */
128'h4503c6ed4711a06d268500e50023954a, /*  733 */
128'h00d90023469500d515630e5006930009, /*  734 */
128'h0037f6930ff7f7930027979b01659663, /*  735 */
128'h946346918bb10107671300b694634585, /*  736 */
128'h00e905a39432920116020087671300d7, /*  737 */
128'hc50500b7c783709c4511bf654701bdfd, /*  738 */
128'hcb890207f7930047f713f4e518e34711, /*  739 */
128'hbf154501e80703e30004bc230004a623, /*  740 */
128'h00b5c7836c8cfbf58b91b73d4515fb0d, /*  741 */
128'hc4c8af2ff0ef0007c503609cdbe58bc1, /*  742 */
128'h46a10ff7f7930027979b05659a63bdb9, /*  743 */
128'h47039722930117020017061b873245ad, /*  744 */
128'h0ae3f95704e3f94706e3f4e374e30007, /*  745 */
128'h4c634185551b0187151b02b6f263fd37, /*  746 */
128'h866300054883fce50513000085170005, /*  747 */
128'h7513fbf7051bbd6d4519f11710e30008, /*  748 */
128'h66e30ff57513f9f7051beea87ae30ff5, /*  749 */
128'h7179bdf90ff777130017e7933701eea8, /*  750 */
128'h451184aef406842ae44ee84aec26f022, /*  751 */
128'h6008a0b1c90de199484c49bd0e500913, /*  752 */
128'hc3210007c7036c1ce1292501afaff0ef, /*  753 */
128'h033780630327026303f7f79300b7c783, /*  754 */
128'h70a2450100979a630017b79317e18bfd, /*  755 */
128'h852245818082614569a2694264e27402, /*  756 */
128'h4511b7cd00042a23d9452501c13ff0ef, /*  757 */
128'hf0ef842ae426ec06e82245811101bfe5, /*  758 */
128'hf0ef6008484c0e500493e50d250188ff, /*  759 */
128'h00978d630007c7836c1ced092501a8cf, /*  760 */
128'h4791dd792501bcdff0ef85224585cb99, /*  761 */
128'h8082610564a2644260e2451d00f51363, /*  762 */
128'h049bfa9ff0ef842aec06e426e8221101, /*  763 */
128'h0005049ba42ff0ef6008484ce49d0005, /*  764 */
128'h700c84cff0ef4581020006136c08e085, /*  765 */
128'h00e782234705601c82aff0ef462d6c08, /*  766 */
128'hed6347858082610564a28526644260e2, /*  767 */
128'h694264e2740270a245098082450900b7, /*  768 */
128'hec26f02271794d1c808261456a0269a2, /*  769 */
128'hfcf5fde384ae842ae052e44ee84af406, /*  770 */
128'hf0ef852285a600f4fa634c1c59fd4a05, /*  771 */
128'h0ce3bf754501000914630005091bec8f, /*  772 */
128'h8afff0ef852285a6460103390763fb49, /*  773 */
128'h4783c81c278501378a63481cf15d2501, /*  774 */
128'hbf5d0009049b00f402a30017e7930054, /*  775 */
128'he432e82efc061028ec2a7139b7594505, /*  776 */
128'h8793000097970405426383eff0eff42e, /*  777 */
128'h0023c3196622631800a78733050eade7, /*  778 */
128'h4501e39897aa00070023c31967620007, /*  779 */
128'hf0ef0828080c460100f618634785cb11, /*  780 */
128'h7175bfe5452d8082612170e22501a0ef, /*  781 */
128'he8daecd6f0d2f4cefca6e122e506f8ca, /*  782 */
128'h84aa89b20005302314050d634925e42e, /*  783 */
128'h10630005091b9d6ff0ef1028002c8a79, /*  784 */
128'h2501b6dff0efe4be1028083c65a21409, /*  785 */
128'h01f9fa1301c9f7934519e011e1196406, /*  786 */
128'he75ff0ef102800f516634791c54dc3e1, /*  787 */
128'hcfcd008a77936406e949008a6a132501, /*  788 */
128'h0ca300f408a302100713046007937aa2, /*  789 */
128'h0b2300e40823000407a30004072300f4, /*  790 */
128'h0e23000405a300e40c2300040ba30004, /*  791 */
128'hc50300040fa300040f2300040ea30004, /*  792 */
128'h0da300040d234785fc9fe0ef85a2000a, /*  793 */
128'h82230005099b00040aa300040a230004, /*  794 */
128'hf0ef030aab03855685ce04098b6300fa, /*  795 */
128'h0135262385da39fd7522e9112501e3ff, /*  796 */
128'h00b44783a895892ac90d250183aff0ef, /*  797 */
128'ha0854921f60981e30049f993e3d98bc5, /*  798 */
128'h0029f993e72d0107f71300b44783f565, /*  799 */
128'h6a13c399008a7793e3ad8b8500098463, /*  800 */
128'h01448523f4800309a78385a279a2020a, /*  801 */
128'hc8c8f33fe0ef0009c503000485a3d09c, /*  802 */
128'ha623c8880069d783dbbfe0ef01c40513, /*  803 */
128'h60aa00f494230134b0230004ae230004, /*  804 */
128'h6b466ae67a0679a6794674e6854a640a, /*  805 */
128'hf8a27119b7d5491db7e5491180826149, /*  806 */
128'hfc5ee0daf0caf4a6fc86e4d6e8d2ecce, /*  807 */
128'h8a2e842a0006a023ec6ef06af466f862, /*  808 */
128'h000998630005099be91fe0ef8ab6e432, /*  809 */
128'h744670e60007899bc39d662200b44783, /*  810 */
128'h7be26b066aa66a4669e6790674a6854e, /*  811 */
128'h00a44783808261096de27d027ca27c42, /*  812 */
128'h40f907bb445c01042903160789638b85, /*  813 */
128'h0b1320000b930006091b00f67463893e, /*  814 */
128'h90631ff777934458fa090ce35c7d0304, /*  815 */
128'hfcb337fd0025478300975c9b60081207, /*  816 */
128'h47854848eb11020c99630ffcfc930197, /*  817 */
128'h4c0cb741498900f405a3478900a7ec63, /*  818 */
128'h05a3478501851763b7e52501bd6ff0ef, /*  819 */
128'h856e4c0c00043d83cc08b7a5498500f4, /*  820 */
128'h0099579b000c861bd5792501b98ff0ef, /*  821 */
128'h002dc683c4b58d3a0007849b00a6073b, /*  822 */
128'h86a6001dc503419684bb00f6f4639fb1, /*  823 */
128'h00a44783f94d250104e050ef85d2863a, /*  824 */
128'h0097fc6341a507bb4c48c3850407f793, /*  825 */
128'h955285da20000613910115020097951b, /*  826 */
128'h9a3e9381020497930094949bc5ffe0ef, /*  827 */
128'h9fa5000aa783c45c9fa54099093b445c, /*  828 */
128'h00a4478304e601634c50b70500faa023, /*  829 */
128'he43a85da4685001dc503c38d0407f793, /*  830 */
128'hf793672200a44783f1392501014050ef, /*  831 */
128'h0017c503863a4685601c00f40523fbf7, /*  832 */
128'h444c01a42e23f11525017c1040ef85da, /*  833 */
128'h0127f46340bb87bb1ff5f5930009049b, /*  834 */
128'he0ef855295a28626030585930007849b, /*  835 */
128'he4cee8caf0a27159b59d499dbf9dbd1f, /*  836 */
128'hec66f062f45ef85aeca6f486fc56e0d2, /*  837 */
128'h8ab689328a2e842a0006a023e46ee86a, /*  838 */
128'h00b44783000997630005099bcb5fe0ef, /*  839 */
128'h694664e6854e740670a60007899bc39d, /*  840 */
128'h6d426ce27c027ba27b427ae26a0669a6, /*  841 */
128'h18078f638b8900a44783808261656da2, /*  842 */
128'h0b1320000b9304f76c630127873b445c, /*  843 */
128'h93631ff777930409046344585c7d0304, /*  844 */
128'hfcb337fd0025478300975c9b60081407, /*  845 */
128'h4581485cef01040c9a630ffcfc930197, /*  846 */
128'h498900f405a3478902e798634705cb91, /*  847 */
128'h445cf3fd0005079bd86ff0ef4c0cb759, /*  848 */
128'h05230207e79300a4478312f76a634818, /*  849 */
128'h498500f405a3478501879763b79500f4, /*  850 */
128'hf79300a44783c85ce311cc1c4858bf99, /*  851 */
128'h85da0017c50346854c50601cc38d0407, /*  852 */
128'hfbf7f79300a44783f96925016b5040ef, /*  853 */
128'h97cff0ef856e4c0c00043d8300f40523, /*  854 */
128'h00a6863b0099579b000c869bd1592501, /*  855 */
128'h74639fb5002dc703c4b58d320007849b, /*  856 */
128'h40ef85d286a6001dc503419704bb00f7, /*  857 */
128'h0297f26341a587bb4c4cf15125016670, /*  858 */
128'h855a95d220000613918115820097959b, /*  859 */
128'h00f40523fbf7f79300a44783a4ffe0ef, /*  860 */
128'h093b445c9a3e9381020497930094949b, /*  861 */
128'h00faa0239fa5000aa783c45c9fa54099, /*  862 */
128'h00e7fa63445c481800c78e634c5cbdd1, /*  863 */
128'hfd0925015cb040ef85da4685001dc503, /*  864 */
128'h87bb1ff575130009049b444801a42e23, /*  865 */
128'h8626030505130007849b0127f46340ab, /*  866 */
128'h0407e79300a447839dbfe0ef952285d2, /*  867 */
128'h1141bd2d499db5f9c81cbf4100f40523, /*  868 */
128'h4783e1752501acffe0ef842ae406e022, /*  869 */
128'h601cc3950407f793cf690207f71300a4, /*  870 */
128'h589040ef030405930017c50346854c50, /*  871 */
128'h00f40523fbf7f79300a44783ed552501, /*  872 */
128'hc703741ce15d2501b77fe0ef6008500c, /*  873 */
128'h0107169b481800e785a30207671300b7, /*  874 */
128'h00d78ea300e78e230086d69b0106d69b, /*  875 */
128'h00e78fa300d78f230187571b0107569b, /*  876 */
128'h169b00e78d2300078ba300078b234858, /*  877 */
128'h0107171b00e78a2327010107571b0107, /*  878 */
128'h0106d69b00e78aa30087571b0107571b, /*  879 */
128'h046007130086d69b00e78c2302100713, /*  880 */
128'h000789a30007892300e78ca300d78da3, /*  881 */
128'h478500f40523fdf7f793600800a44783, /*  882 */
128'h4505ebbfe06f014160a2640200f50223, /*  883 */
128'h842ae406e022114180820141640260a2, /*  884 */
128'h25019cbfe0ef8522e9012501effff0ef, /*  885 */
128'h110180820141640260a200043023e119, /*  886 */
128'h879700054a6395bfe0efec060028e42a, /*  887 */
128'h452d8082610560e2450140a785230000, /*  888 */
128'hf486f0a21028002c4601e42a7159bfe5, /*  889 */
128'h083c65a2ec190005041bb3bfe0efeca6, /*  890 */
128'h6586e41d0005041bcd2ff0efe4be1028, /*  891 */
128'h64e6740670a68522cbd8575277a2e991, /*  892 */
128'hc50374a2cb998bc100b5c78380826165, /*  893 */
128'hfcf41ee34791b7c5c8c897bfe0ef0004, /*  894 */
128'hf8cae122e506e42afca67175bfd94415, /*  895 */
128'h1828002c460184ae00050023f0d2f4ce, /*  896 */
128'h842677e2ecbe081ce5292501acdfe0ef, /*  897 */
128'h040a12634a16c2be02f009934bdc597d, /*  898 */
128'h071b3527470300008717e50567a24501, /*  899 */
128'h186300e780a303a0071300e780230307, /*  900 */
128'h00078023078d00e7812302f007130e94, /*  901 */
128'h808261497a0679a6794674e6640a60aa, /*  902 */
128'h18284581fd452501f89fe0ef18284585, /*  903 */
128'h0007c50365c677e2f5552501e6eff0ef, /*  904 */
128'h2501f63fe0ef18284581c2aa8cdfe0ef, /*  905 */
128'h77e2e1052501e48ff0ef18284581f949, /*  906 */
128'h01450e6325018a7fe0ef0007c50365c6, /*  907 */
128'h67a24711dd612501a9eff0ef18284581, /*  908 */
128'hf5cfe0ef1828100cb7594509f8e516e3, /*  909 */
128'hfc974703973610949301020797134781, /*  910 */
128'h05bbfff7871b04e462630037871beb05, /*  911 */
128'h96b2920166a20206961300e586bb40f4, /*  912 */
128'hb7319c3d01368023fff7c79301271a63, /*  913 */
128'h4603962a1088920102071613b7c12785, /*  914 */
128'h0789bddd4545b7e900c68023377dfc96, /*  915 */
128'h07850007470397369281020416936722, /*  916 */
128'hf8227139b709fe9465e3fee78fa32405, /*  917 */
128'h84ae842ae456e852ec4efc06f04af426, /*  918 */
128'h00b44783000917630005091bfb4fe0ef, /*  919 */
128'h790274a2854a744270e20007891bcf89, /*  920 */
128'h009777634818808261216aa26a4269e2, /*  921 */
128'h00042623445884bae3918b8900a44783, /*  922 */
128'h00a44783c81cfcf778e34818445ce4bd, /*  923 */
128'hf793445c4481bf7d00f405230207e793, /*  924 */
128'h099300a44783fc960ee34c50d3e51ff7, /*  925 */
128'hc50385ce4685601cc3850407f7930304, /*  926 */
128'hf79300a44783ed512501213040ef0017, /*  927 */
128'h0017c50386264685601c00f40523fbf7, /*  928 */
128'h6008bf59cc44ed3525011c1040ef85ce, /*  929 */
128'hfff4869b377dc7290097999b00254783, /*  930 */
128'h413007bb02c6ed630337563b0336d6bb, /*  931 */
128'h4a855a7dd1c19c9dc45c27814c0c8ff9, /*  932 */
128'hd7b51ff4f793c45c9fa5445c0499ea63, /*  933 */
128'h9ca90094d49bcd112501c87fe0ef6008, /*  934 */
128'h47850005059b814ff0efe595484cbfb1, /*  935 */
128'h57fdbded490900f405a3478900f59763, /*  936 */
128'hc84cb5ed490500f405a3478500f59763, /*  937 */
128'he0efcb818b89600800a44783b765cc0c, /*  938 */
128'hc4bfe0efbf6984cee5990005059bfddf, /*  939 */
128'h4f9c601cfabafee3fd4588e30005059b, /*  940 */
128'h013787bb413484bbcc0c445cfaf5fae3, /*  941 */
128'h842ac52de42ef822fc067139b7bdc45c, /*  942 */
128'h67e2e1152501fe6fe0ef0828002c4601, /*  943 */
128'h250197cff0eff01c101ce01c852265a2, /*  944 */
128'h4515e7898bc100b5c783cd996c0ce529, /*  945 */
128'he30fe0ef0007c50367e2a02d00043023, /*  946 */
128'h00f414230067d7838522458167e2c448, /*  947 */
128'h70e2f971fcf50be347912501cbdfe0ef, /*  948 */
128'hfcf501e34791bfdd4525808261217442, /*  949 */
128'h2501dbafe0ef842ae406e0221141b7c1, /*  950 */
128'h717980820141640260a200043023e119, /*  951 */
128'hd98fe0ef892e842af406e84aec26f022, /*  952 */
128'he0ef8522458100091f63e8890005049b, /*  953 */
128'h64e269428526740270a20005049bc5ff, /*  954 */
128'hb32ff0ef852245810224302380826145, /*  955 */
128'h852285ca00042a2302f5136347912501, /*  956 */
128'h47912501f8bfe0ef85224581c68fe0ef, /*  957 */
128'hbf6584aad16dbf7d00042a2300f51663, /*  958 */
128'hf0a21028002c460184aee42aeca67159, /*  959 */
128'h083c65a2e00d0005041bedafe0eff486, /*  960 */
128'h6786e8010005041b872ff0efe4be1028, /*  961 */
128'h70a68522c10fe0ef102885a6c489cf81, /*  962 */
128'hf0a27159bfcd44198082616564e67406, /*  963 */
128'he0d28522002c46018b2ee42af85a8432, /*  964 */
128'hec66f062f45efc56e4cee8caeca6f486, /*  965 */
128'h2c836000000a1c6300050a1be7cfe0ef, /*  966 */
128'h00fb202302f76263ffec871b481c0184, /*  967 */
128'h7ae26a0669a6694664e68552740670a6, /*  968 */
128'h00044b83808261656ce27c027ba27b42, /*  969 */
128'h85ca4a8559fd4481490902fb9f634785, /*  970 */
128'h09550863093508632501a55fe0ef8522, /*  971 */
128'h00544783fef963e329054c1c2485e111, /*  972 */
128'hb74d009b202300f402a30017e793c804, /*  973 */
128'h1afd4c0944814981490110000ab7504c, /*  974 */
128'h2501d10fe0ef0015899b852200099e63, /*  975 */
128'h038b9163200009930344091385cee921, /*  976 */
128'he3918fd90087979b0009470300194783, /*  977 */
128'h854ab745fc0c94e33cfd39f909092485, /*  978 */
128'he1116582015575332501abcfe0efe02e, /*  979 */
128'hbfbd4a09b7494a05b7c539f109112485, /*  980 */
128'h842ae04aec06e426e8221101bfad8a2a, /*  981 */
128'hcb9100b44783e4910005049bbc4fe0ef, /*  982 */
128'h610564a269028526644260e20007849b, /*  983 */
128'h48144458cf390027f71300a447838082, /*  984 */
128'h600800f40523c8180207e793fed772e3, /*  985 */
128'hc53900042a232501a58ff0ef484cef01, /*  986 */
128'h091b94dfe0ef4c0cbf7d84aa00a405a3, /*  987 */
128'h06374c0cb7dd450502f9146357fd0005, /*  988 */
128'h85ca6008f9792501b37fe0ef167d1000, /*  989 */
128'h45094785b769449db7e12501a1cff0ef, /*  990 */
128'h00a44783fcf96ae34d1c6008fcf900e3, /*  991 */
128'h0017c50346854c50601cdba50407f793, /*  992 */
128'h00a44783f55d25015f0040ef03040593, /*  993 */
128'h4605e42a7175b7b100f40523fbf7f793, /*  994 */
128'hca0fe0eff8cafca6e122e5061008002c, /*  995 */
128'he3bfe0efe0be1008081c65a2e9052501, /*  996 */
128'h0207f79300b7c78345196786e1052501, /*  997 */
128'hcb810014f79300b5c483c59975e2eb89, /*  998 */
128'h790280826149794674e6640a60aa451d, /*  999 */
128'h88c1cc0d0005041bad8fe0ef00094503, /* 1000 */
128'h100c02800613fc878de301492783c89d, /* 1001 */
128'h951fe0efcaa200a8458996cfe0ef00a8, /* 1002 */
128'hd94d2501836ff0ef00a84581f1612501, /* 1003 */
128'hf15525019f5fe0ef1008faf518e34791, /* 1004 */
128'h85a27502bf612501f20fe0ef7502e411, /* 1005 */
128'h4605e42a7171b769d575250191cff0ef, /* 1006 */
128'he152e54ee94aed26f506f1221028002c, /* 1007 */
128'hbd0fe0efe8eaece6f0e2f4def8dafcd6, /* 1008 */
128'he4be1028083c65a21c0414630005041b, /* 1009 */
128'h176347911c0409630005041bd67fe0ef, /* 1010 */
128'h9f630207f79300b7c783441967a61af4, /* 1011 */
128'h02630005091bb45fe0ef458175221807, /* 1012 */
128'h0b63440557fd16f90f63440947851809, /* 1013 */
128'h160414630005041ba98fe0ef752216f9, /* 1014 */
128'h0a13f6efe0ef85220109549b85ca7422, /* 1015 */
128'he0ef855200050c1b4581200006130344, /* 1016 */
128'h248188cfe0ef855202000593462d898f, /* 1017 */
128'h0fa30104949b0109199b0ff4fb1347c1, /* 1018 */
128'h0b930104d49b021007930109d99b02f4, /* 1019 */
128'hd99b046007930ff97a9304f4062302e0, /* 1020 */
128'h0a230200061304f406a30084d49b0089, /* 1021 */
128'h07a305540723040405a3040405230374, /* 1022 */
128'h0544051385d2049404a3056404230534, /* 1023 */
128'h00074603468d05740aa3772280efe0ef, /* 1024 */
128'h0723478100f69363571400d6166357d2, /* 1025 */
128'h06f4042327810107d79b0107969b06f4, /* 1026 */
128'h0086d69b0107d79b0106d69b0107979b, /* 1027 */
128'h00274b8306f404a306d407a30087d79b, /* 1028 */
128'h0005041bf59fe0ef1028040b99634c85, /* 1029 */
128'h0210071300e785a3752247416786e835, /* 1030 */
128'h00078ba300078b230460071300e78c23, /* 1031 */
128'h01678a2301378da301578d2300e78ca3, /* 1032 */
128'h041bd5afe0ef00f50223478500978aa3, /* 1033 */
128'h022303852823001c0d1b7522a82d0005, /* 1034 */
128'h20000613ec090005041b8dcfe0ef0195, /* 1035 */
128'h8c6a0ffbfb93f61fd0ef3bfd85524581, /* 1036 */
128'h70aa8522f25fe0ef85ca7522441db749, /* 1037 */
128'h7ba67b467ae66a0a69aa694a64ea740a, /* 1038 */
128'h7159b7c544218082614d6d466ce67c06, /* 1039 */
128'h10284605002c843284aee42aeca6f0a2, /* 1040 */
128'h1028083c65a2e13125019cafe0eff486, /* 1041 */
128'hc783451967a6e9152501b65fe0efe4be, /* 1042 */
128'h00b74783c30d6706e39d0207f79300b7, /* 1043 */
128'h008705a38c3d027474138c658cbd7522, /* 1044 */
128'h740670a62501c9efe0ef00f502234785, /* 1045 */
128'h002c4605e02ee42a71718082616564e6, /* 1046 */
128'h0005079b964fe0efed26f122f5060088, /* 1047 */
128'hf0be083cf4be008865a2678612079663, /* 1048 */
128'hc703778610079a630005079baf7fe0ef, /* 1049 */
128'h479165e61007126302077713479900b7, /* 1050 */
128'h0613e55fd0ef102805ad46550e058e63, /* 1051 */
128'hf05fd0ef850ae49fd0ef10a8008c0280, /* 1052 */
128'h079baadfe0ef10a865820c054d6347ad, /* 1053 */
128'hdc5fe0ef10a80ce793634711cbf90005, /* 1054 */
128'h851302a10593464d648aefc50005079b, /* 1055 */
128'h0207e793640602814783e0dfd0ef00d4, /* 1056 */
128'h8bc100b4c78300f40223478500f485a3, /* 1057 */
128'h85a60004450306f7086357d64736cbbd, /* 1058 */
128'h059bcaefe0ef85220005059bf2dfd0ef, /* 1059 */
128'h0005079bfc3fd0ef8522c5a547890005, /* 1060 */
128'h02f69d630557468302e007936706efb1, /* 1061 */
128'h27810107d79b06f707230107969b57d6, /* 1062 */
128'h0087d79b0107d79b0107979b06f70423, /* 1063 */
128'h07a3478506f704a30086d69b0106d69b, /* 1064 */
128'h0005079be24fe0ef008800f7022306d7, /* 1065 */
128'h740a70aa0005079bb50fe0ef6506e791, /* 1066 */
128'he8a2711dbfcd47a18082614d853e64ea, /* 1067 */
128'h810fe0efec861028002c4605842ee42a, /* 1068 */
128'h9abfe0efe4be1028083c65a2e9292501, /* 1069 */
128'h0207f79300b7c783451967a6e1292501, /* 1070 */
128'h00e78b23752200645703cb856786eb95, /* 1071 */
128'h00e78c230044570300e78ba30087571b, /* 1072 */
128'he0ef00f50223478500e78ca30087571b, /* 1073 */
128'he4a6711d80826125644660e62501ad6f, /* 1074 */
128'he8a208284601002c893284aee42ae0ca, /* 1075 */
128'h4581c4b9e0510005041bf9bfd0efec86, /* 1076 */
128'h08284585e5592501ca8fe0efd2020828, /* 1077 */
128'hd0ef8526462d75c2e93d2501b8ffe0ef, /* 1078 */
128'h000700230200061346ad00b48713ca1f, /* 1079 */
128'h97a6938117820007869bfff6879bce89, /* 1080 */
128'h656202090a63fec783e3177d0007c783, /* 1081 */
128'h470d6562e0150005041be69fd0ef510c, /* 1082 */
128'h0270079300e684630005468304300793, /* 1083 */
128'h852200a92023c29fd0ef953e03478793, /* 1084 */
128'h1563479180826125690664a6644660e6, /* 1085 */
128'he42a711db7d5842abf550004802300f5, /* 1086 */
128'h041bee3fd0efec86e8a21028002c4605, /* 1087 */
128'h02061793460100010c2366a2ec550005, /* 1088 */
128'hea2902000593eba10007c78397b69381, /* 1089 */
128'he8410005041bbd6fe0efda0210284581, /* 1090 */
128'h01814783e1792501abbfe0ef10284585, /* 1091 */
128'h07136786bc7fd0ef082c462dc3dd6506, /* 1092 */
128'h8ba300078b230460071300e78c230210, /* 1093 */
128'hbf45863eb74d2605a06100e78ca30007, /* 1094 */
128'h000747039736930102079713fff6079b, /* 1095 */
128'h07f00e9343658e2e4781082cfeb706e3, /* 1096 */
128'h91411542f9f7051b27850006c70348b1, /* 1097 */
128'h05130000751793411742370100a36c63, /* 1098 */
128'h8522441900eef863a82100070f1b9e65, /* 1099 */
128'h48030505bfcdf36d80826125644660e6, /* 1100 */
128'h00fe06b3b7cdffe81be3060805630005, /* 1101 */
128'h752200f500235795a885078500c68023, /* 1102 */
128'hb7c10005041b8fefe0ef00f502234785, /* 1103 */
128'he0ef1028dbd50181478302f51b634791, /* 1104 */
128'h4581020006136506f4450005041ba55f, /* 1105 */
128'h6786ae5fd0ef082c462d6506b07fd0ef, /* 1106 */
128'hf91780e3b751842abf1900e785a34721, /* 1107 */
128'h93811782f4c7e5e30585068500e58023, /* 1108 */
128'h4703f8d771e30007869b020006134729, /* 1109 */
128'h05052e83bf89eaf71de30e5007930181, /* 1110 */
128'hec22110105c528830585230305452e03, /* 1111 */
128'h87f2869a8646040502938f2ae44ae826, /* 1112 */
128'h8dfd00c6c5b316ef8f9300005f978876, /* 1113 */
128'h008fa403000f2583000fa38300b64733, /* 1114 */
128'h004f2703ff4fa3839db9007585bb0fc1, /* 1115 */
128'h0105e8330198581b0078159b0105883b, /* 1116 */
128'h8e6d00f6c6339f3100f805bb0077073b, /* 1117 */
128'h0146561b00c6171b9e39008f23838e35, /* 1118 */
128'hc6b300d383bb00c5873b008383bb8e59, /* 1119 */
128'hd39b007686bb8ebd00cf24038ef900b7, /* 1120 */
128'hffcfa4039fa100d3e6b30116969b00f6, /* 1121 */
128'h9fa1007777338f2d0007061b00d703bb, /* 1122 */
128'h0f418f5d0167171b00a7579b9f3d8f2d, /* 1123 */
128'hf45f17e300e387bb0003869b0005881b, /* 1124 */
128'h0e8f8f9300005f971b05859300005597, /* 1125 */
128'h00cf7f3300d7cf331b02829300005297, /* 1126 */
128'h0025c4030015c383000faf0301e6c733, /* 1127 */
128'h972a070a93aa038a0005c70300ef0f3b, /* 1128 */
128'h083b004fa70300ef0f3b942a040a4318, /* 1129 */
128'h0003a70301b8581b9e3900581f1b010f, /* 1130 */
128'h8e7501e7c6339f3100f80f3b010f6833, /* 1131 */
128'h0176561b0096139b008fa7039e398e3d, /* 1132 */
128'h05919f3500cf03bb00c3e63340189eb9, /* 1133 */
128'h0fc101e6c6b3fff5c4838efd007f46b3, /* 1134 */
128'h9fb900e6941b94aa048affcfa7039eb9, /* 1135 */
128'hc7339fb900d3843b8ec140980126d69b, /* 1136 */
128'h00c7579b9f3d0077473301e777330083, /* 1137 */
128'h069b0003861b000f081b8f5d0147171b, /* 1138 */
128'h0f1300005f17f25599e300e407bb0004, /* 1139 */
128'h010fc40303c38393000053978ffa0c6f, /* 1140 */
128'h00c2c4b3942a040a00d7c2b30003a703, /* 1141 */
128'h048a0043a4039f21011fc4839f254000, /* 1142 */
128'h171b012fc4830107083b40809e2194aa, /* 1143 */
128'h0083a4039e210107683301c8581b0048, /* 1144 */
128'h863b9ea194aa00e2c2b3048a00f8073b, /* 1145 */
128'h0156561b013fc90300b6129b408000c2, /* 1146 */
128'hffc3a4839c3500c702bb03c100c2e633, /* 1147 */
128'h941b992a9ea1090a0056c6b300e7c6b3, /* 1148 */
128'h843b8ec1000924830106d69b9fa50106, /* 1149 */
128'h9f3d8f219fa5005747330007081b00d2, /* 1150 */
128'h0002861b0f918f5d0177171b0097579b, /* 1151 */
128'h00005297f5f592e300e407bb0004069b, /* 1152 */
128'ha70300d745b38f5dfff64713fb428293, /* 1153 */
128'h020f45839f2d022f4403021f43830002, /* 1154 */
128'h9f2d942a040a418c95aa058a93aa038a, /* 1155 */
128'ha5839e2d0068171b0107083b0042a583, /* 1156 */
128'h9db100f8073b0107683301a8581b0003, /* 1157 */
128'h139b0082a5839e2d8e3d8e59fff6c613, /* 1158 */
128'h03bb00c3e633400c9ead0166561b00a6, /* 1159 */
128'h0075e5b3fff7c593023f44839ead00c7, /* 1160 */
128'h00f5969b048a9db5ffc2a4038db902c1, /* 1161 */
128'h00b385bb40809fa18dd50115d59b94aa, /* 1162 */
128'h007747339fa18f4dfff747130007081b, /* 1163 */
128'h861b0f118f5d0157171b00b7579b9f3d, /* 1164 */
128'h6462f3ef9de300e587bb0005869b0003, /* 1165 */
128'h00c8863b00d306bb00fe07bb010e883b, /* 1166 */
128'h6105692264c2cd70cd34c97c05052823, /* 1167 */
128'he85af44ef84afc26e0a2715d653c8082, /* 1168 */
128'h84aa97b203f7f413ec56f052e486e45e, /* 1169 */
128'h07bb04000b9304000b13e53c893289ae, /* 1170 */
128'h0a1b00f974639381178200078a1b408b, /* 1171 */
128'h0084853385ce020ada93020a1a930009, /* 1172 */
128'h99d641590933481020ef0144043b8656, /* 1173 */
128'h60a6b7c997824401852660bc01741763, /* 1174 */
128'h6ba26b426ae27a0279a2794274e26406, /* 1175 */
128'h842a03f7f793f0227179653c80826161, /* 1176 */
128'hf800071300178513e84af406e44eec26, /* 1177 */
128'h40a9863b449d0400099300e7802397a2, /* 1178 */
128'h3c9020ef95224581920116020006091b, /* 1179 */
128'h97828522603cfc1c078e643c0124f563, /* 1180 */
128'h69a2694264e2740270a2fd24fde34501, /* 1181 */
128'h3423639cf94787930000779780826145, /* 1182 */
128'hed3c639cf8c7879300007797e93c0405, /* 1183 */
128'h059311018082e13cb6c7879300000797, /* 1184 */
128'h769747013bf020efec06850a46410505, /* 1185 */
128'h454147a5859300006597172686930000, /* 1186 */
128'h0047d613070506890007c78300e107b3, /* 1187 */
128'h8f230007c78397ae000646038bbd962e, /* 1188 */
128'h0000751760e2fca71de3fef68fa3fec6, /* 1189 */
128'h0808842ae12271758082610513450513, /* 1190 */
128'hf0ef080885a26622f71ff0efe42ee506, /* 1191 */
128'h60aaf83ff0ef0808f01ff0ef0808e85f, /* 1192 */
128'h00d70d63711c46a1595880826149640a, /* 1193 */
128'h80824501cf980200071300d717634691, /* 1194 */
128'he426e82211018082556dbfe50007ac23, /* 1195 */
128'h569702f5026384ae842a200007b7ec06, /* 1196 */
128'h85930000659708800613d62686930000, /* 1197 */
128'hfc2409f030ef3ee50513000065173de5, /* 1198 */
128'h6100e82211018082610564a2644260e2, /* 1199 */
128'h569702f4026384ae200007b7ec06e426, /* 1200 */
128'h85930000659702f00613d3a686930000, /* 1201 */
128'he00405f030ef3ae505130000651739e5, /* 1202 */
128'h6100e82211018082610564a2644260e2, /* 1203 */
128'h569702f4026384ae200007b7ec06e426, /* 1204 */
128'h85930000659703600613d0a686930000, /* 1205 */
128'he40401f030ef36e505130000651735e5, /* 1206 */
128'h6104e42611018082610564a2644260e2, /* 1207 */
128'h769702f48263842e200007b7ec06e822, /* 1208 */
128'h85930000659703e00613eb2686930000, /* 1209 */
128'h14027de030ef32e505130000651731e5, /* 1210 */
128'h11018082610564a2644260e2e8809001, /* 1211 */
128'h8263842e200007b7ec06e8226104e426, /* 1212 */
128'h659704500613e66686930000769702f4, /* 1213 */
128'h30ef2ea50513000065172da585930000, /* 1214 */
128'h610564a2644260e2ec809001140279a0, /* 1215 */
128'h200007b7ec06e4266100e82211018082, /* 1216 */
128'h0613c52686930000569702f4026384ae, /* 1217 */
128'h051300006517296585930000659704c0, /* 1218 */
128'h610564a2644260e2f004756030ef2a65, /* 1219 */
128'h200007b7ec06e4266100e82211018082, /* 1220 */
128'h0613c22686930000569702f4026384ae, /* 1221 */
128'h05130000651725658593000065970530, /* 1222 */
128'h610564a2644260e2f404716030ef2665, /* 1223 */
128'hf04af426f82200053983ec4e71398082, /* 1224 */
128'h02f984638436893284ae200007b7fc06, /* 1225 */
128'h0000659705a00613be86869300005697, /* 1226 */
128'h30efe43a21c505130000651720c58593, /* 1227 */
128'h0029191b8b0589890014159b67226ca0, /* 1228 */
128'h88a10125e5b30034949b8dd900497913, /* 1229 */
128'h69e2790274a202b9b8238dc5744270e2, /* 1230 */
128'h4605468147057100e022114180826121, /* 1231 */
128'hf0ef45818522f7dff0efe40645818522, /* 1232 */
128'hf67ff0ef45814605468547058522f35f, /* 1233 */
128'h01414501640260a2d97ff0ef45816008, /* 1234 */
128'h3c23460546814705e022e40611418082, /* 1235 */
128'h8522f39ff0ef842a4581040530230205, /* 1236 */
128'h46054685470545818522ef1ff0ef4581, /* 1237 */
128'hf06f0141458160a264026008f23ff0ef, /* 1238 */
128'h200007b7ec06e8226104e4261101d4df, /* 1239 */
128'h0613b12686930000569702f48263842e, /* 1240 */
128'h05130000651712658593000065970610, /* 1241 */
128'h644260e2fc80904114425e6030ef1365, /* 1242 */
128'hec06e8226104e42611018082610564a2, /* 1243 */
128'h86930000569702f48263842e200007b7, /* 1244 */
128'h65170e2585930000659706800613ade6, /* 1245 */
128'h8c7d17fd67855a2030ef0f2505130000, /* 1246 */
128'he82211018082610564a2644260e2e0a0, /* 1247 */
128'h02f4026384ae200007b7ec06e4266100, /* 1248 */
128'h0000659706f00613aa86869300005697, /* 1249 */
128'h55c030ef0ac505130000651709c58593, /* 1250 */
128'he04a11018082610564a2644260e2e424, /* 1251 */
128'h842a200007b7ec06e426e82200053903, /* 1252 */
128'h0613a72686930000569702f9026384ae, /* 1253 */
128'h05130000651705658593000065970760, /* 1254 */
128'h644260e2c84404993c23516030ef0665, /* 1255 */
128'heca67100f0a2715980826105690264a2, /* 1256 */
128'hf062f45ef85afc56e0d2e4cef486e8ca, /* 1257 */
128'he03084b2892e0005d783020408a3ec66, /* 1258 */
128'h9c636ca020ef00c9051345814611d01c, /* 1259 */
128'h07b700043983bf5ff0ef458560080e04, /* 1260 */
128'h44810049278316f99a6304043a032000, /* 1261 */
128'h4c1c4485e391448d8b89c7090017f713, /* 1262 */
128'h8b85008a2783000a09638cdd03243c23, /* 1263 */
128'h45814605468147050144e49316078663, /* 1264 */
128'h2583be1ff0ef85224581d71ff0ef8522, /* 1265 */
128'hc4fff0ef9ecc0c1300005c1785220089, /* 1266 */
128'hf0eff82a0a1300006a17852200095583, /* 1267 */
128'hf0ef85224581cbdff0ef852285a6c81f, /* 1268 */
128'hd27ff0ef85224581460546854705cf5f, /* 1269 */
128'h4585e93ff0ef852224058593000f45b7, /* 1270 */
128'h009899b785220d89b583cd1ff0ef8522, /* 1271 */
128'h6a9768198993eb7ff0ef25810015e593, /* 1272 */
128'h64e6740670a6efe9485cf42a8a930000, /* 1273 */
128'h6ce27c027ba27b427ae26a0669a66946, /* 1274 */
128'hdb7ff0efe024852244cc808261654501, /* 1275 */
128'hee079be38b85449cdf3ff0ef8522488c, /* 1276 */
128'h458163900107e683654100043883603c, /* 1277 */
128'h6e89f005051300ff0e37431147014781, /* 1278 */
128'h183b070500371f1b00064803ec0689e3, /* 1279 */
128'h0067036316fd060527810107e7b301e8, /* 1280 */
128'h981b010767330187971b0187d81bf2e5, /* 1281 */
128'h8fe9010767330087d79b01c878330087, /* 1282 */
128'h9746938183751782170200be873b8fd9, /* 1283 */
128'h869300005697b765470147812585e31c, /* 1284 */
128'h6517e6258593000065971490061388e6, /* 1285 */
128'h00c4e493bd85322030efe72505130000, /* 1286 */
128'h5597000b1d633b7d20000bb78b4ebd61, /* 1287 */
128'h00efe625051300006517872585930000, /* 1288 */
128'h061386e20179096300043903b7116f60, /* 1289 */
128'h485c070934832e2030ef855685d20f20, /* 1290 */
128'h37830209370312048e6324818cfd4c81, /* 1291 */
128'hcc5cf9200793c7817c1c00f76f630c89, /* 1292 */
128'hb27ff0ef85224581b6fff0ef85224581, /* 1293 */
128'hff397913852201442903c3950044f793, /* 1294 */
128'h0000651785cad47ff0ef85ca00896913, /* 1295 */
128'h2903c3950084f793680000efe0450513, /* 1296 */
128'hf0ef85ca00496913ff39791385220144, /* 1297 */
128'h658000efe04505130000651785cad1ff, /* 1298 */
128'h8c630384390300043c83cfb50014f793, /* 1299 */
128'h85d209c006137de6869300004697017c, /* 1300 */
128'h3c2300492783cba97c1c236030ef8556, /* 1301 */
128'h018c871308e69f630037f693470d0204, /* 1302 */
128'hff87051363104591480d468100c90793, /* 1303 */
128'h8361ff87370301068763c3900086161b, /* 1304 */
128'h603cfeb690e30791872a2685c3988f51, /* 1305 */
128'hc85c9bf9485cc85c0027e793485ccbb5, /* 1306 */
128'h01748c63040439036004cc9d4c858889, /* 1307 */
128'h855685d20ca006137786869300004697, /* 1308 */
128'h0089278300090963040430231b8030ef, /* 1309 */
128'h9bf54c85485cb4dff0ef8522ef8d8b85, /* 1310 */
128'h4505d80c8ee3c47ff0ef8522484cc85c, /* 1311 */
128'h2623000cb783dbd98b85bd955d5020ef, /* 1312 */
128'h97a667a1bf41b1dff0ef8522b77100f9, /* 1313 */
128'h8913fa978de394be00093c8301096483, /* 1314 */
128'h39a020efe43e002c46218566639c0087, /* 1315 */
128'h0513717908b041635535b7dd87ca0ca1, /* 1316 */
128'h892e84b2e44ef406e84aec26f0220480, /* 1317 */
128'h0000451785a2cc1d5551842a0a8030ef, /* 1318 */
128'h6517862285aa89aa785010ef6e450513, /* 1319 */
128'h07b702098b634fe000efcd2505130000, /* 1320 */
128'hcb990024f793f40401242423e01c2000, /* 1321 */
128'h69a2694264e2740270a24501c45c4789, /* 1322 */
128'hb7e5c45c4785d4fd4501888580826145, /* 1323 */
128'h458146098082bff9557d090030ef8522, /* 1324 */
128'h953e050e200007b7f73ff06f20000537, /* 1325 */
128'he4066380e0221141711c808225016108, /* 1326 */
128'h680686930000469702f40263200007b7, /* 1327 */
128'h00006517bb4585930000659734c00613, /* 1328 */
128'h557de3914505703c074030efbc450513, /* 1329 */
128'h4501842ae822110180820141640260a2, /* 1330 */
128'h60e26622644285a24d3010efe42eec06, /* 1331 */
128'hf4062000051371797940006f61054685, /* 1332 */
128'h84aa7af020efe052e44ee84aec26f022, /* 1333 */
128'h0001b5030b6030efc285051300006517, /* 1334 */
128'h206010ef842a491010ef450144b010ef, /* 1335 */
128'h3f8000ef638cc0e5051300006517681c, /* 1336 */
128'h3e8000efc0c505130000651706f44583, /* 1337 */
128'h15c20085d59bc165051300006517546c, /* 1338 */
128'h0000651706c44583583c3d2000ef91c1, /* 1339 */
128'h0187d61b0107d69b0087d71bc0c50513, /* 1340 */
128'h00ef26010ff6f6930ff7f7930ff77713, /* 1341 */
128'h398000efbfc50513000065175c0c3a60, /* 1342 */
128'h00006597c789b865859300006597545c, /* 1343 */
128'h378000efbec5051300006517b7458593, /* 1344 */
128'h65977448006030efbf85051300006517, /* 1345 */
128'h584c19c42783db9fb0ef152585930000, /* 1346 */
128'h061300006617e789b506061300006617, /* 1347 */
128'h852633a000efbd65051300006517eae6, /* 1348 */
128'h0a1300006a174481ed5ff0ef84264581, /* 1349 */
128'hf79320000913bd69899300006997bd6a, /* 1350 */
128'h0004458330c000ef855285a6e78901f4, /* 1351 */
128'h04052fa000ef819100f5f6132485854e, /* 1352 */
128'h2e8000ef0dc5051300006517fd249fe3, /* 1353 */
128'h614545016a0269a2694264e2740270a2, /* 1354 */
128'h07b30003b6830083b7830103b7038082, /* 1355 */
128'h0017079300d7fe6393811782278540f7, /* 1356 */
128'h802345050103b78300a7002300f3b823, /* 1357 */
128'h0103b7830083b7038082450180820007, /* 1358 */
128'hfff706930003b7038f99920102059613, /* 1359 */
128'h86bb87aa9d9dfff7059b00c6f5638e9d, /* 1360 */
128'h852e0007002300b6e6630103b70340a7, /* 1361 */
128'h07850007c68300d3b823001706938082, /* 1362 */
128'h053be681000556634881bfe900d70023, /* 1363 */
128'hf81304100693c21906100693488540a0, /* 1364 */
128'h02b6733b0005061b385986ba4e250ff6, /* 1365 */
128'h02b6563b0305051b046e67630ff37513, /* 1366 */
128'h85bbfe718532fea68fa306850ff57513, /* 1367 */
128'h07930008876302f5e9630300051340e6, /* 1368 */
128'h0015559b40e6853b068500f6802302d0, /* 1369 */
128'h00b61b63fff5081b86ba258100068023, /* 1370 */
128'h2585fea68fa30685bf5d00a8053b8082, /* 1371 */
128'h0007c30397ba9381178240c807bbb7d9, /* 1372 */
128'h0685011780230066802326050006c883, /* 1373 */
128'heccef4a6f8a2597d011cf0ca7119b7f1, /* 1374 */
128'hf42afc3e843684b2e0dafc86e4d6e8d2, /* 1375 */
128'h03000a9306c00a1302500993f82af02e, /* 1376 */
128'hc52d8f1d0004c50377a2774202095913, /* 1377 */
128'h086304d7ff639381178276820017079b, /* 1378 */
128'hc503bfe1e7bff0ef0201039304850135, /* 1379 */
128'hc783035510634781048905450f630014, /* 1380 */
128'hf36346a50ff7f793fd07879bcb9d0004, /* 1381 */
128'h0f630640069304890014c503478100f6, /* 1382 */
128'h079304d50f630580069302a6eb6306d5, /* 1383 */
128'h790674a6744670e6f55d08f509630630, /* 1384 */
128'h808261090007051b6b066aa66a4669e6, /* 1385 */
128'h06e50e6307300713b74d048d0024c503, /* 1386 */
128'h00840b13f6e51ee30700071300a76c63, /* 1387 */
128'h02e5006307500713a00d460146850038, /* 1388 */
128'h00840b13fa850613f6e510e307800713, /* 1389 */
128'hf8b50693a81145c10016361346850038, /* 1390 */
128'h400845a946010016b693003800840b13, /* 1391 */
128'hf0ef0028020103930005059be37ff0ef, /* 1392 */
128'h00840b130201039300044503a809ddbf, /* 1393 */
128'h7433600000840b13b5fd845ad93ff0ef, /* 1394 */
128'h020103930005059b4db010ef85220124, /* 1395 */
128'hfc3ef83aec061034f436715db7f18522, /* 1396 */
128'h8082616160e2e8dff0efe436e4c6e0c2, /* 1397 */
128'hec06100005931014862ef436f032715d, /* 1398 */
128'h60e2e69ff0efe436e4c6e0c2fc3ef83a, /* 1399 */
128'h1234862afe36fa32f62e710d80826161, /* 1400 */
128'heac2e6bee2baea22ee06080810000593, /* 1401 */
128'h0bd020ef0808842ae3fff0efe436eec6, /* 1402 */
128'hb303679c691c80826135645260f28522, /* 1403 */
128'hee63479d808245018302000303630087, /* 1404 */
128'h83f91da70713000047170205979304b7, /* 1405 */
128'h878297bae426e822ec061101439c97ba, /* 1406 */
128'h97930c5010ef7540f55c08c52483795c, /* 1407 */
128'he91c64a2644260e202f457b393810204, /* 1408 */
128'h35f1bfd9617cbfe97d5c808261054501, /* 1409 */
128'h557d8082557db7e9659c95aa058e05e1, /* 1410 */
128'h5e63ff5ff0ef842ae406e02211418082, /* 1411 */
128'h8522000307630207b303679c681c0005, /* 1412 */
128'h0141640260a245018302014160a26402, /* 1413 */
128'h4797150200a7eb6347ad8082557d8082, /* 1414 */
128'h551780826108953e8175162787930000, /* 1415 */
128'h0007b303679c691c80827d2505130000, /* 1416 */
128'h4785d23e47d502f1102347a1715d8302, /* 1417 */
128'h100c200007930030e83ee42e07851782, /* 1418 */
128'h8082616160a6fd3ff0efcc3ed402e486, /* 1419 */
128'h45018082450100e6fe63400407374d14, /* 1420 */
128'h24010113228134832301340323813083, /* 1421 */
128'h980101f1041322813823dc0101138082, /* 1422 */
128'hf0ef1a05348322113c232291342385a2, /* 1423 */
128'h02f71c630a0447830a04c703f579f95f, /* 1424 */
128'h0c04c70302f716630dd447830dd4c703, /* 1425 */
128'h0e0447830e04c70302f710630c044783, /* 1426 */
128'h10ef0d4485130d440593461100f71a63, /* 1427 */
128'h842af0227179b761fb600513d55156f0, /* 1428 */
128'h858a4601852267e020eff4063e800513, /* 1429 */
128'he509842af21ff0efc202c40200011023, /* 1430 */
128'h6145740270a28522660020ef7d000513, /* 1431 */
128'hf406f022478500f11023478571798082, /* 1432 */
128'h008007b745386914c195842ac402c23e, /* 1433 */
128'h8f75600006b78ff58ff9f80787934ad4, /* 1434 */
128'h8522858a4601c43e8fd98f55400006b7, /* 1435 */
128'h6145740270a2c43c47b2e119ec9ff0ef, /* 1436 */
128'h5783c23e47d500f1102347b5711d8082, /* 1437 */
128'hfdf949370107979bf852fc4ee0ca07c5, /* 1438 */
128'h842e8aaaec86f456e4a6e8a26a056989, /* 1439 */
128'he00a0a13e0098993080909134495c43e, /* 1440 */
128'hf79345b2ed0de73ff0ef8556858a4601, /* 1441 */
128'h0125f7b3054793630135f7b3c7891005, /* 1442 */
128'h0513d4bff0ef62e5051300005517c78d, /* 1443 */
128'h7aa27a4279e2690664a6644660e6fba0, /* 1444 */
128'h0014079b347dfe04c6e334fd80826125, /* 1445 */
128'h4501b75556c020ef3e80051300f05763, /* 1446 */
128'hd09ff0ef6045051300005517fc8049e3, /* 1447 */
128'h47c17139e7a919c52783bf7df9200513, /* 1448 */
128'hfc06f822858a460147d5c42e00f11023, /* 1449 */
128'h1b842783c11dde3ff0efc23e842af426, /* 1450 */
128'hdcdff0ef8522858a46014495cb918b89, /* 1451 */
128'h8082612174a2744270e2f8ed34fdc901, /* 1452 */
128'hec86e0cae4a6711d80824501bfd54501, /* 1453 */
128'h270347c906d7f66384b6892a4785e8a2, /* 1454 */
128'hd432cf3108c92783260102f1102302c9, /* 1455 */
128'hd23a854a100c47850030cc3ee42e4755, /* 1456 */
128'hf0634785e529842ad75ff0efc83eca26, /* 1457 */
128'h854a100c47f5460102f1102347b10497, /* 1458 */
128'h051300005517c11dd55ff0efd23ed402, /* 1459 */
128'h690664a6644660e68522c43ff0ef55e5, /* 1460 */
128'h841bb74d02f6063bbf6147c580826125, /* 1461 */
128'hf426f822fc067139b7c54401b7d50004, /* 1462 */
128'h8a2e4148842ace05e456e852ec4ef04a, /* 1463 */
128'h00b44583c11d892a482010ef8ab684b2, /* 1464 */
128'h014485b3681000054d638e3fa0ef8522, /* 1465 */
128'hbd9ff0ef514505130000551700b67a63, /* 1466 */
128'hf96decdff0ef854a08c92583a0894481, /* 1467 */
128'h844e0089f3630207e4030109378389a6, /* 1468 */
128'hfc851ae3f01ff0ef854a85d6865286a2, /* 1469 */
128'h9aa2028784339a22408989b308c96783, /* 1470 */
128'h69e274a279028526744270e2fc0999e3, /* 1471 */
128'h00f1102347997139808261216aa26a42, /* 1472 */
128'h161b8edd030007b70086969bc23e47f5, /* 1473 */
128'h440dc43684aafc06f426f8228ed10106, /* 1474 */
128'h3e800593e919c53ff0ef8526858a4601, /* 1475 */
128'h8082612174a2744270e2d91ff0ef8526, /* 1476 */
128'hbffc07b7db0101134d18bfcdfc79347d, /* 1477 */
128'h3c2324813023241134239fb923213823, /* 1478 */
128'h1ce7f56349013ffc0737233134232291, /* 1479 */
128'h892ac09ff0ef84aa85a2980101f10413, /* 1480 */
128'h20ef20000513e7991a04b7831e051863, /* 1481 */
128'h06131e0503631a04b5031aa4b02366a0, /* 1482 */
128'h6b6347210c044783123010ef85a22000, /* 1483 */
128'h53b897ba078ad0e70713000047171cf7, /* 1484 */
128'h278300e7fd63cc981ff78793400407b7, /* 1485 */
128'h73630147d69307a68007071367050d44, /* 1486 */
128'h06f48f2309b449830a044783f8dc00d7, /* 1487 */
128'h4783c7890e244783e7810019f9938b85, /* 1488 */
128'h8b890a04478300098a6308f480a30b34, /* 1489 */
128'h07130e24478306f48fa309c44783c789, /* 1490 */
128'h05130a844783fcdc07c60c8486130914, /* 1491 */
128'h00074583fff74783e0fc07c6468109d4, /* 1492 */
128'h97aeffe745839fad0105959b0087979b, /* 1493 */
128'h02f585b30e04458300098c634685c391, /* 1494 */
128'h0621070de21c07ce02b787b30dd44783, /* 1495 */
128'h08d4470308e4478304098f63fca714e3, /* 1496 */
128'h08c447039fb90087171b0107979b4685, /* 1497 */
128'h87b30dd4478302f707330e04470397ba, /* 1498 */
128'h979b08a4470308b44783f8fc07ce02e7, /* 1499 */
128'h0087171b089447039fb90107171b0187, /* 1500 */
128'h07a6c319f4fc54d89fb9088447039fb9, /* 1501 */
128'h8bfd09c44783c7898b850a044783f4fc, /* 1502 */
128'hf0ef852645850af006134685ce81e391, /* 1503 */
128'h46830af447830af407a34785ed35e0bf, /* 1504 */
128'h54dc08f4aa2300a6979bc7b98b850e04, /* 1505 */
128'h4783f8dc07a60d44278300098663c799, /* 1506 */
128'h478308d4ac2302f686bb00a6969b0dd4, /* 1507 */
128'h854a240134032481308308f480230a74, /* 1508 */
128'h25010113228139832301390323813483, /* 1509 */
128'h8bfd8b7d0057d79b00a7d71b50fc8082, /* 1510 */
128'h892abf4d08f4aa2302f707bb27852705, /* 1511 */
128'hbf651a04b0234cc020efd1691a04b503, /* 1512 */
128'h22113c23dc010113bf455929bf555951, /* 1513 */
128'h88634789232130232291342322813823, /* 1514 */
128'h2381308354a9c585468102b7e16302f5, /* 1515 */
128'h01132281348322013903852623013403, /* 1516 */
128'h4685fef760e34705ffc5879b80822401, /* 1517 */
128'h84aad1fff0ef892a45850b900613842e, /* 1518 */
128'h01f10413f1e9258199f5ffe4059bf571, /* 1519 */
128'h0b944783e51998dff0ef854a85a29801, /* 1520 */
128'hec267179b74d84aab75ddf400493f7d5, /* 1521 */
128'h0ff5f99308154783f022f406e44ee84a, /* 1522 */
128'h45850b3006138edd892e9be10079f693, /* 1523 */
128'h00f51e63842a57b5c519cc7ff0ef84aa, /* 1524 */
128'h8526842a875ff0ef852685ca00091c63, /* 1525 */
128'h64e2740270a28522013505a315e010ef, /* 1526 */
128'h28113c23d60101138082614569a26942, /* 1527 */
128'h27313c23292130232891342328813823, /* 1528 */
128'h25713c23276130232751342327413823, /* 1529 */
128'h23b13c2325a130232591342325813823, /* 1530 */
128'hbff7879bbffc07b74d180ac7e9634789, /* 1531 */
128'h84ae8b32892abfe787933ffc07b79f3d, /* 1532 */
128'h07e9460300e7eb631185051300005517, /* 1533 */
128'hf0ef13a5051300005517e7b900167793, /* 1534 */
128'h29013403298130838522f8400413f96f, /* 1535 */
128'h27013a03278139832801390328813483, /* 1536 */
128'h25013c0325813b8326013b0326813a83, /* 1537 */
128'h2a01011323813d8324013d0324813c83, /* 1538 */
128'hdb451125051300005517098927038082, /* 1539 */
128'hac83e79102eaf7bb060a81630045aa83, /* 1540 */
128'h1185051300005517cb8902ecf7bb0005, /* 1541 */
128'h02eadabb02c92783bf415429f24ff0ef, /* 1542 */
128'h856200c488138c0a009c9c9be3994b85, /* 1543 */
128'h0017859b000828834e114e85478189d6, /* 1544 */
128'h110505130000551700030d6302e8f33b, /* 1545 */
128'hd33bb7f14b814a814c81b7c1ee4ff0ef, /* 1546 */
128'hc78397a6078e020880630065202302e8, /* 1547 */
128'hfb9300dbebb300be96bbcb898b850107, /* 1548 */
128'hfbc596e387ae05110821013309bb0ffb, /* 1549 */
128'h00e30f250513000055178a09000b8963, /* 1550 */
128'hf0ef854a85d2fe0a7a1302f10a13f006, /* 1551 */
128'h09ea478309fa4603ee0519e3842af94f, /* 1552 */
128'h963e09da47839e3d0087979b0106161b, /* 1553 */
128'hf0ef0e2505130000551785ce01367a63, /* 1554 */
128'h0017f7130a7a46830084c783b5c1e56f, /* 1555 */
128'h0016e993c3990fe6f9938b89c71989b6, /* 1556 */
128'h4b189726070e0017059b461145054701, /* 1557 */
128'h00b517bb02080463001878130017581b, /* 1558 */
128'hd79b8b050189999b0187979b0027571b, /* 1559 */
128'h0ff9f99300f9e9b3c70d4189d99b4187, /* 1560 */
128'h8b850a6a478302d98263fcc592e3872e, /* 1561 */
128'hb591274020ef0965051300005517ef89, /* 1562 */
128'h8b8509ba4783bfd100f9f9b3fff7c793, /* 1563 */
128'h547ddbaff0ef0c65051300005517cb89, /* 1564 */
128'h4685e3958b850afa4783e20b02e3b51d, /* 1565 */
128'h4785e569a21ff0ef854a45850af00613, /* 1566 */
128'h08f92a2300a7979b0e0a47830afa07a3, /* 1567 */
128'hf69301acd6bb08c00d934d0108800493, /* 1568 */
128'h2485ed499f1ff0ef854a458586260ff6, /* 1569 */
128'h08f00d134c81ffb492e32d210ff4f493, /* 1570 */
128'hf0ef854a458586260ff6f693019ad6bb, /* 1571 */
128'hffa492e32ca10ff4f4932485e9359cbf, /* 1572 */
128'h8656000c26834c818aa609b00d934d61, /* 1573 */
128'h99dff0ef854a0ff6f6930196d6bb4585, /* 1574 */
128'h248dffac90e30ffafa932ca12a85e139, /* 1575 */
128'h09c0061386defdb498e30c110ff4f493, /* 1576 */
128'hd4fb0de34785ed19975ff0ef854a4585, /* 1577 */
128'h458509b00613468501379b630a7a4783, /* 1578 */
128'h0a70061386cebb3d842a957ff0ef854a, /* 1579 */
128'h1141b32ddd79842a945ff0ef854a4585, /* 1580 */
128'h681c00055e63810ff0ef842ae406e022, /* 1581 */
128'h60a264028522000307630187b303679c, /* 1582 */
128'h713980820141640260a2450583020141, /* 1583 */
128'h00f5866384aa4791f04af822fc06f426, /* 1584 */
128'h00f110230370079304f5926355294785, /* 1585 */
128'h858a46010107979b4955842e07c4d783, /* 1586 */
128'h10234799ed19d52ff0efc43ec24a8526, /* 1587 */
128'h4601c43e478900f41f634791c24a00f1, /* 1588 */
128'h790274a2744270e2d34ff0ef8526858a, /* 1589 */
128'hee09b7cdc402fef414e3478580826121, /* 1590 */
128'h85be27814f1887ae00f5f3634f5c6918, /* 1591 */
128'hf06f02c50823dd0c0007059b00e7f463, /* 1592 */
128'h4b9c711910000737691c80828082c2cf, /* 1593 */
128'he4d6e8d2eccef0caf4a6fc86f8a2070d, /* 1594 */
128'hf0ef842ac17c8fd9f466f862fc5ee0da, /* 1595 */
128'h02042423eb8d6b9c679c681cc509f11f, /* 1596 */
128'hf8500493bacff0efed85051300005517, /* 1597 */
128'h6aa66a4669e674a679068526744670e6, /* 1598 */
128'h4481541c808261097ca27c427be26b06, /* 1599 */
128'h082347851af42c23478df93ff0eff3e5, /* 1600 */
128'h7d000513ba2ff0ef852202042c2302f4, /* 1601 */
128'h84aa97826b9c679c8522681c3b5010ef, /* 1602 */
128'h22231a04282318042e2308842783f945, /* 1603 */
128'h45814601b72ff0ef8522d85c478508f4, /* 1604 */
128'hf14984aacf2ff0ef8522f1dff0ef8522, /* 1605 */
128'h00f1102347a1000505a345d000ef8522, /* 1606 */
128'he3991aa007138ff94bdc00ff8737681c, /* 1607 */
128'hc23ec43a8522858a460147d50aa00713, /* 1608 */
128'h15630aa0079300c14703e911bf8ff0ef, /* 1609 */
128'h037009933e900913cc1c800207b700f7, /* 1610 */
128'h80020c3700ff8bb74b0502900a934a55, /* 1611 */
128'hc252013110238522858a460140000cb7, /* 1612 */
128'h015110234c18681ce13dbb6ff0efc402, /* 1613 */
128'he7b301871563c43e0177f7b3c25a4bdc, /* 1614 */
128'hed1db8eff0ef8522858a4601c43e0197, /* 1615 */
128'h3e80051306090863397d0007ca6347b2, /* 1616 */
128'h00e68563800207374c14bf452c5010ef, /* 1617 */
128'hd45c8b8541e7d79bc43ccc1880010737, /* 1618 */
128'hf9200793b55d18f40ca3478506041e23, /* 1619 */
128'hf0ef85224581c04ff0ef852202f51f63, /* 1620 */
128'h18f40c2347850007d663443ced09c34f, /* 1621 */
128'h00005517d965c1cff0ef85224585bfd1, /* 1622 */
128'h84aab595fa100493a10ff0efd5450513, /* 1623 */
128'he74eeb4aef26f706f3227161551cb585, /* 1624 */
128'he6eeeaeaeee6f2e2f6defadafed6e352, /* 1625 */
128'h199bc783193010ef45018baae3b54401, /* 1626 */
128'h10234789e7b5180b8ca3198bc783c7b1, /* 1627 */
128'hf0efc482c2be855e008c479d460104f1, /* 1628 */
128'hcf818b851b8ba783120500e3842aabaf, /* 1629 */
128'h03e3842aaa0ff0ef855e008c46014495, /* 1630 */
128'hf0ef855ea031020ba423f4fd34fd1005, /* 1631 */
128'h695a64fa741a70ba8522d55d842ad99f, /* 1632 */
128'h6d566cf67c167bb67b567af66a1a69ba, /* 1633 */
128'hc163180b8c23048ba7838082615d6db6, /* 1634 */
128'h1493101010ef4501b16ff0ef855e0407, /* 1635 */
128'hb36ff0ef855e45853e80091390810205, /* 1636 */
128'h10ef85260007cc63048ba783f155842a, /* 1637 */
128'hbfe916b010ef0640051312a96ee30dd0, /* 1638 */
128'h41e7d79b048ba78300fbac23400007b7, /* 1639 */
128'h450dbf0506fb9e23478502fba6238b85, /* 1640 */
128'ha029400406370ea61ee345111aa60f63, /* 1641 */
128'h0036d61b00cbac234006061b40010637, /* 1642 */
128'h964e068a8a3d31e98993000039978a9d, /* 1643 */
128'h018ba88345051086a6830f86460396ce, /* 1644 */
128'hae231a0ba8238a0500c7d61b02d606bb, /* 1645 */
128'hd69b08dba22308dba42304cba823180b, /* 1646 */
128'h1408dc63090ba62300d5183b8abd0107, /* 1647 */
128'h0107979b14068e6302cba683090ba823, /* 1648 */
128'h938117828fd98ff50107571b003f06b7, /* 1649 */
128'hbc23030787b300e797b3070907854721, /* 1650 */
128'hbc230c0bb8230c0bb4230c0bb0230a0b, /* 1651 */
128'hd463200007930afbb8230e0bb0230c0b, /* 1652 */
128'hf46320000793090ba70308fba6230107, /* 1653 */
128'h8e63577d04cba783c21508fba82300e7, /* 1654 */
128'h1023855e008c46010107979b471100e7, /* 1655 */
128'h04f11023479d902ff0efc282c4be04e1, /* 1656 */
128'h855e008c0107979b4601495507cbd783, /* 1657 */
128'h4785e40516e3842a8e4ff0efc4bec2ca, /* 1658 */
128'hc9aff0ef855e08fb80a357fd08fbaa23, /* 1659 */
128'h00b545830f7000ef855ee2051ae3842a, /* 1660 */
128'h018ba703e0051fe3842affbfe0ef855e, /* 1661 */
128'h079304fba0232789100007b754075a63, /* 1662 */
128'h979b108c460107cbd78306f110230370, /* 1663 */
128'hd2caed05880ff0efd4bed2ca855e0107, /* 1664 */
128'h988102091a93033007930bf104934905, /* 1665 */
128'h108c08104b210a854a11d48206f11023, /* 1666 */
128'h3a7dc131850ff0efd05aec56e826855e, /* 1667 */
128'h0637a7a940020637bb45842afe0a16e3, /* 1668 */
128'ha82300b515bb89bd0165d59bbd994003, /* 1669 */
128'h569b8ff50027979b16f16685b54d08bb, /* 1670 */
128'hb5558b1d938100f7571b17828fd501e7, /* 1671 */
128'h161b0187179b0187569b00ff05374098, /* 1672 */
128'h06138fd167410087569b8e698fd50087, /* 1673 */
128'h559b40d804fbaa2327818fd58ef1f007, /* 1674 */
128'h571b8de90087159b8ecd0187169b0187, /* 1675 */
128'h0187d71b04ebac238f558f718ecd0087, /* 1676 */
128'h8001073720d702634689212700638b3d, /* 1677 */
128'h040ba7830007596302d7971300ebac23, /* 1678 */
128'h07b7018ba70304fba0238fd920000737, /* 1679 */
128'h639c08278793000057971ef718638001, /* 1680 */
128'h020d1a13044ba783f0be4d05040ba903, /* 1681 */
128'h0ff1079300f979331384849300003497, /* 1682 */
128'h97bb478540980a05fe07fc1383f97913, /* 1683 */
128'h017d8b3716078563278100f977b300e7, /* 1684 */
128'h40dc0007ac8397d6109c840b0b1b4a81, /* 1685 */
128'h400007b7140781630197f7b300f977b3, /* 1686 */
128'h00fc88634591200007b700fc8d6345a1, /* 1687 */
128'hf0ef855e0015b59340bc85b3100005b7, /* 1688 */
128'h8d6347a1400007370e051c638daa971f, /* 1689 */
128'h100007b700ec886347912000073700ec, /* 1690 */
128'he0ef855e02fbaa23001cb79340fc8cb3, /* 1691 */
128'h4d850ce79163470d01a78663409cdfdf, /* 1692 */
128'h2d81810007b7d33e47d50af110234799, /* 1693 */
128'h110c040007930110d53e00fde7b317c1, /* 1694 */
128'h4783e941e91fe0efc93ee552e162855e, /* 1695 */
128'h9a631afba823409c09b794638bbd010c, /* 1696 */
128'h08bba2230017b79317ed088ba5831407, /* 1697 */
128'h0ff10793947ff0ef855e460118fbae23, /* 1698 */
128'h07cbd7830af1102303700793fe07fd93, /* 1699 */
128'hd33a8cee855e110c0107979b46014755, /* 1700 */
128'h102347b56702e915e35fe0efd53ee03a, /* 1701 */
128'h110c0110040007134791d502d33a0af1, /* 1702 */
128'he0dfe0efe03ac93ae552e16ee43e855e, /* 1703 */
128'h85b74785f3ed37fd670267a20e050c63, /* 1704 */
128'h4601180bae23096ba2231afba823017d, /* 1705 */
128'h94e347a10a918c9ff0ef855e84058593, /* 1706 */
128'he6f49fe3fb4787930000379704a1eafa, /* 1707 */
128'hdf400413cbdfe0ef8305051300005517, /* 1708 */
128'h80020737b519a007071b80011737b61d, /* 1709 */
128'h80030737de075ee30307971300ebac23, /* 1710 */
128'h9881190201000ab70ff104934905bbc5, /* 1711 */
128'h10234799020a08633a7d09053ac54a15, /* 1712 */
128'h855e010c040007931030c33e47d508f1, /* 1713 */
128'hd0051ce3d61fe0efdc3ef84af426c556, /* 1714 */
128'hf006869366c144dcfbe18b8583a54cdc, /* 1715 */
128'h02e796938fd18ff50087d79b0087961b, /* 1716 */
128'h04fba02300876793da06d9e3040ba703, /* 1717 */
128'h837902079713eaf768e34581472db35d, /* 1718 */
128'h0537040d859366c1b54511872583974e, /* 1719 */
128'h0187d61b0d91000da783f006869300ff, /* 1720 */
128'h0087d79b8e690087961b8f510187971b, /* 1721 */
128'ha703fdb59ee3fefdae238fd98ff58f51, /* 1722 */
128'ha60300f6f8638bbd00c7579b46a5008c, /* 1723 */
128'h86930000369704d61c63800306b7018b, /* 1724 */
128'hae230087171b1487a78397b6078ae066, /* 1725 */
128'h0186d61b8ff917fd67c100cca68308fb, /* 1726 */
128'hc305c38d03f7771327810126d71b8fd1, /* 1727 */
128'h57bb8a8d0106d69b02e6073b3e800613, /* 1728 */
128'ha7830adba2230afba02302d606bb02f7, /* 1729 */
128'h20000793c79919cba7831afbaa231b0b, /* 1730 */
128'h1523484000ef855e08fba82308fba623, /* 1731 */
128'hd6b7aaaab7b708cba703000506230005, /* 1732 */
128'h27818ef98ff9ccc68693aaa78793cccc, /* 1733 */
128'hf0f0f6b79fb500f037b3068600d036b3, /* 1734 */
128'h06b79fb5068a00d036b38ef90f068693, /* 1735 */
128'h9fb5068e00d036b38ef9f0068693ff01, /* 1736 */
128'h9fb9071200e037338f750207161376c1, /* 1737 */
128'hd70302c7d7b3ed1092010a8bb783d11c, /* 1738 */
128'h0000459784aa06fbc603074bd68307ab, /* 1739 */
128'ha95fe0effef536230245051366c58593, /* 1740 */
128'h0088579b06cbc603077bc883070ba803, /* 1741 */
128'h0ff878130ff7f7930188569b0108571b, /* 1742 */
128'h851364a585930000459726810ff77713, /* 1743 */
128'h859300004597074ba603a5ffe0ef04d4, /* 1744 */
128'h8abd0146561b0106569b062485136465, /* 1745 */
128'ha42347856e8010ef8526a3ffe0ef8a3d, /* 1746 */
128'h07b704fba0232785100007b7b8d102fb, /* 1747 */
128'h00004517e691ecf76ce31a0bb6834004, /* 1748 */
128'ha0230017079b70000737bb955c450513, /* 1749 */
128'hf6931adba42303f7f6930c46c78304fb, /* 1750 */
128'ha0230217071bc68900c7f693ce910027, /* 1751 */
128'h8b8504eba02301076713040ba70304eb, /* 1752 */
128'haa0304fba02300c7e793040ba783c799, /* 1753 */
128'h7a33855e4601088ba583044ba783040b, /* 1754 */
128'h4a85db4ff0efcb6484930000349700fa, /* 1755 */
128'h8c9300003c974c2dcc8b0b1300003b17, /* 1756 */
128'hcbb5278100fa77b300fa97bb409ccfac, /* 1757 */
128'h10000db720000d37ca89091300003917, /* 1758 */
128'h04f718630017b79317ed00494703409c, /* 1759 */
128'h4683c3a18ff900fa77b30009270340dc, /* 1760 */
128'he0ef855e0fb6f69345850b7006130089, /* 1761 */
128'he0ef855e45850b7006134681c131debf, /* 1762 */
128'ha223180bae231a0ba823088ba783ddbf, /* 1763 */
128'h11e30931973fe0ef855e035baa2308fb, /* 1764 */
128'h4985051300004517f7649fe304a1fb99, /* 1765 */
128'h4721400006b700092783bb6d925fe0ef, /* 1766 */
128'hb71341b787b301a78663471100d78963, /* 1767 */
128'h855e408c933fe0ef855e02ebaa230017, /* 1768 */
128'he79d0046f79300892683f941808ff0ef, /* 1769 */
128'hb79317ed088ba583ef8d1afba823409c, /* 1770 */
128'hf0ef855e460118fbae2308bba2230017, /* 1771 */
128'h0ff6f693bb91fd319fdfe0ef855ecb0f, /* 1772 */
128'hb7c9f521d31fe0ef855e45850b700613, /* 1773 */
128'h2583974e837902079713fcfc65e34581, /* 1774 */
128'h6da000ef06cb851300ec4641bf6d1187, /* 1775 */
128'h979b008c460107cbd78304f11023478d, /* 1776 */
128'h842a96ffe0efc2be47d5855ec4be0107, /* 1777 */
128'h04e157830007d663018ba783ec051b63, /* 1778 */
128'hd783c2be479d04f1102347a506fb9e23, /* 1779 */
128'he0efc4be855e0107979b008c460107cb, /* 1780 */
128'h45e6475647c646b6ea051163842a93bf, /* 1781 */
128'h06eba22306fba02304dbae23018ba503, /* 1782 */
128'h01a6d61bf2c51a634000063706bba423, /* 1783 */
128'h09634505f0c543638ca602e345098a3d, /* 1784 */
128'h0413f0eff06f2006061b40010637f0a6, /* 1785 */
128'h8082557d80824501c56ce54ff06ffa10, /* 1786 */
128'h879300005797808218b50d238082557d, /* 1787 */
128'h842ae406e02247851141ef9d439cbfa7, /* 1788 */
128'he0ef852212a000efbef7222300005717, /* 1789 */
128'h02c00513fc5ff0ef852200055563aeef, /* 1790 */
128'h01414501640260a20dc000ef13e000ef, /* 1791 */
128'h631cbb27071300005717808245018082, /* 1792 */
128'h05130000451785aa114102e790636394, /* 1793 */
128'h0141853e478160a2f60fe0efe4064465, /* 1794 */
128'h853ebfd187b600a604630fc7a6038082, /* 1795 */
128'hc105fbdff0efe42eec06110141488082, /* 1796 */
128'h07930815470302b7006365a210354703, /* 1797 */
128'h5535eb3fe06f610560e200f70c630ff0, /* 1798 */
128'hbfcdf8400513bfe545018082610560e2, /* 1799 */
128'hcd09f7dff0ef84aee822ec06e4261101, /* 1800 */
128'h60e2e0800f840413e501cf0ff0ef842a, /* 1801 */
128'h00005797bfd555358082610564a26442, /* 1802 */
128'h05138082c3980015071b438899c78793, /* 1803 */
128'h80824388984787930000579780820f85, /* 1804 */
128'he4266380e822ae678793000057971101, /* 1805 */
128'h610564a2644260e20094176384beec06, /* 1806 */
128'h6000a9cff0ef8522c78119a447838082, /* 1807 */
128'h5797e79ce39cab67879300005797b7d5, /* 1808 */
128'h879300005797e50880829207ad230000, /* 1809 */
128'h711d8082e308e518e11ce7886798a9e7, /* 1810 */
128'hfc4e6080e8a2a864849300005497e4a6, /* 1811 */
128'hec86e06ae466e862ec5ef05af456f852, /* 1812 */
128'h00004a97334a0a1300004a1789aae0ca, /* 1813 */
128'h00004b9732cb0b1300004b17324a8a93, /* 1814 */
128'h8c0c8c9300004c9700050c1b32cb8b93, /* 1815 */
128'h79e2690664a660e66446029415634d29, /* 1816 */
128'h45176d026ca26c426be27b027aa27a42, /* 1817 */
128'h4901541cddcfe06f61253d2505130000, /* 1818 */
128'h2603681c89560007c36389524c1cc791, /* 1819 */
128'h85ca00090663dbefe0ef638c855a0fc4, /* 1820 */
128'h856685e200978e63601cdb2fe0ef855e, /* 1821 */
128'h848505130000451701a98863da4fe0ef, /* 1822 */
128'he426ec06e8221101b771600022e010ef, /* 1823 */
128'hcbbd4d5ccfad44014d1cc1414401e04a, /* 1824 */
128'h84aa892ec7ad639cc7bd651ccbad511c, /* 1825 */
128'h57fdcd21842a104010ef45051c000593, /* 1826 */
128'he90410f502a347850ef52c234799c57c, /* 1827 */
128'hfffff797e65ff0ef0405282303253023, /* 1828 */
128'h1c2787930000179716f43c2391c78793, /* 1829 */
128'h18f434231b2787930000179718f43023, /* 1830 */
128'h10f400230247c78385220ea42e23681c, /* 1831 */
128'h6105690264a2644260e28522e99ff0ef, /* 1832 */
128'h611c6fa68693000046970c00106f8082, /* 1833 */
128'he11897360017671302d786b365186294, /* 1834 */
128'h07b300f7553b93ed836d8f3d0127d713, /* 1835 */
128'h00005517808225018d5d00f717bb40f0, /* 1836 */
128'hf0efe022e4061141fc3ff06f8fc50513, /* 1837 */
128'h60a28d410105151bfe9ff0ef842afeff, /* 1838 */
128'hf0efe022e40611418082014125016402, /* 1839 */
128'h15029001fd1ff0ef14020005041bfdbf, /* 1840 */
128'hc703058587aa80820141640260a28d41, /* 1841 */
128'h87aa962a8082fb75fee78fa30785fff5, /* 1842 */
128'hfee78fa30785fff5c703058500c78963, /* 1843 */
128'heb09001786930007c70387aa8082fb65, /* 1844 */
128'h8082fb75fee78fa30785fff5c7030585, /* 1845 */
128'h0007c70387b68082e21987aab7d587b6, /* 1846 */
128'h8713fff5c6830585963efb7d00178693, /* 1847 */
128'h80a300c715638082e291fed70fa30017, /* 1848 */
128'hc783000547030585b7cd87ba80820007, /* 1849 */
128'he3994187d79b0187979b40f707bbfff5, /* 1850 */
128'h478100c59463962e8082853ef37d0505, /* 1851 */
128'h40f707bbfff5c783000547030585a839, /* 1852 */
128'h853eff790505e3994187d79b0187979b, /* 1853 */
128'h808200b79363000547830ff5f5938082, /* 1854 */
128'h47830ff5f59380824501bfcd0505c399, /* 1855 */
128'h87aabfcd0505dffd808200b793630005, /* 1856 */
128'hbfcd0785808240a78533e7010007c703, /* 1857 */
128'h65a2fe5ff0efec06842ae42ee8221101, /* 1858 */
128'h157d00b78663000547830ff5f5939522, /* 1859 */
128'h95aa80826105644260e24501fe857be3, /* 1860 */
128'h40a78533e7010007c70300b7856387aa, /* 1861 */
128'h85330007c68387aa862ab7fd07858082, /* 1862 */
128'h000748030705fed80fe38082ea9940c7, /* 1863 */
128'h87aa86aabfcd872eb7d50785fe081be3, /* 1864 */
128'h00c80a638082ea1140d785330007c603, /* 1865 */
128'hbfd5872e8082fe081be3000748030705, /* 1866 */
128'h8fe380824501eb1900054703bff90785, /* 1867 */
128'h87aeb7e50505fafd0007c6830785fee6, /* 1868 */
128'he519842a84aeec06e426e8221101bfd5, /* 1869 */
128'h85a68522cc1163806f87879300004797, /* 1870 */
128'h00004797ef8100044783942af9dff0ef, /* 1871 */
128'h610564a2644260e2852244016c07be23, /* 1872 */
128'h00054783c519f9fff0ef852285a68082, /* 1873 */
128'h6aa7b82300004797050500050023c781, /* 1874 */
128'h842ac891e822ec066104e4261101bfd9, /* 1875 */
128'he008050500050023c501f73ff0ef8526, /* 1876 */
128'h4783c11d8082610564a28526644260e2, /* 1877 */
128'h0017c703ce810007c68387aacf990005, /* 1878 */
128'hb7e5078900d780a300e780238082e311, /* 1879 */
128'h9063963e87aacb9d0075779380824501, /* 1880 */
128'h08b3872aff6d377d8fd507a2808204c7, /* 1881 */
128'h003657930106ef6340e88833469d00c5, /* 1882 */
128'h4725bfc1963a97aa078e02e787335761, /* 1883 */
128'h0785bfe1fef73c230721bfd10ff5f693, /* 1884 */
128'h8b9d00a5e7b300b50a63bf6dfeb78fa3, /* 1885 */
128'h38030721808202c79e63963e87aacb9d, /* 1886 */
128'hff06e8e340f88833ff07bc2307a1ff87, /* 1887 */
128'h963e95ba070e02f707b357e100365713, /* 1888 */
128'h469d00c508b387aa872ebfc100e507b3, /* 1889 */
128'hbf65fee78fa30785fff5c7030585bfe1, /* 1890 */
128'he84af406e432ec26852e842af0227179, /* 1891 */
128'h6582892ace1184aa6622dcdff0efe02e, /* 1892 */
128'hf0ef944a864a8522fff6091300c56463, /* 1893 */
128'h64e269428526740270a200040023f79f, /* 1894 */
128'h00a5e963842ae406e022114180826145, /* 1895 */
128'h95b280820141640260a28522f57ff0ef, /* 1896 */
128'h15fdd7e500e587b340b6073300c506b3, /* 1897 */
128'h1563962ab7fd00f6802316fd0005c783, /* 1898 */
128'h0005c703000547838082853e478100c5, /* 1899 */
128'h00c51363962ab7dd05850505fbed9f99, /* 1900 */
128'h7179bfc50505feb78de3000547838082, /* 1901 */
128'h89aee84af406e44eec26852e842af022, /* 1902 */
128'hd13ff0ef8522c8890005049bd1fff0ef, /* 1903 */
128'h740270a28522440100995b630005091b, /* 1904 */
128'h852285ce86268082614569a2694264e2, /* 1905 */
128'hf593962abfe90405d175f8bff0ef397d, /* 1906 */
128'h0793000547038082450100c514630ff5, /* 1907 */
128'h0ff5f59347c1b7ed853efeb70be30015, /* 1908 */
128'h8082853e4781e60187aa260100c7ef63, /* 1909 */
128'h7713b7f5367d0785feb71ce30007c703, /* 1910 */
128'h87aa0007069b40e7873b47a1c31d0075, /* 1911 */
128'h1793faf5078536fdfcb81ce30007c803, /* 1912 */
128'h00b7e733008597938e1d953e93810207, /* 1913 */
128'h8edd00365713020796938fd901071793, /* 1914 */
128'h1fe30007c703d24d8a1deb1187aa2701, /* 1915 */
128'h008785130007b803bfcd367d0785f8b7, /* 1916 */
128'h1be30785f8b712e30007c70300d80a63, /* 1917 */
128'h4703e7a9419cb7f1377d87aabfa5fef5, /* 1918 */
128'h27970015470308f71163030007930005, /* 1919 */
128'h8a850006c68300e786b3e02787930000, /* 1920 */
128'h1b63078006930ff777130207071bc689, /* 1921 */
128'h0447f7930007c78397ba0025470304d7, /* 1922 */
128'h470302f71c6347c14198c19c47c1c3b1, /* 1923 */
128'h27170015478302f71663030007930005, /* 1924 */
128'hc7098b0500074703973edb2707130000, /* 1925 */
128'h00e79363078007130ff7f7930207879b, /* 1926 */
128'he8221101bf6d47a9bf7d47a180820509, /* 1927 */
128'h00c16583f63ff0efc632ec06006c842e, /* 1928 */
128'h079b00054703d6e80813000028174681, /* 1929 */
128'h9863044678930006460300f806330007, /* 1930 */
128'h7893808261058536644260e2ec050008, /* 1931 */
128'h86b3feb7f4e3fd07879b00088b630046, /* 1932 */
128'hfe07079bc6098a09b7d196be050502d5, /* 1933 */
128'h7139b7e1e008b7cdfc97879b0ff7f793, /* 1934 */
128'h842ae42e00063023f04afc06f426f822, /* 1935 */
128'h744270e25529e90165a2b0dff0ef84b2, /* 1936 */
128'h8522082c892a862e80826121790274a2, /* 1937 */
128'hcb010007c703fe8782e367e2f5dff0ef, /* 1938 */
128'he088fcf718e347a9fd279be307858f81, /* 1939 */
128'h00e6846302d0071300054683b7e94501, /* 1940 */
128'h60a2f23ff0efe40605051141f2dff06f, /* 1941 */
128'h842ee406e02211418082014140a00533, /* 1942 */
128'h04630007c70304b00693601cf0dff0ef, /* 1943 */
128'h60a202d70e630470069300e6ea6302d7, /* 1944 */
128'h069302d7076304d00693808201416402, /* 1945 */
128'h052a069007130017c683fed716e306b0, /* 1946 */
128'h00e69863042007130027c683fce69fe3, /* 1947 */
128'hbfd50789bff1052a052ab7e9e01c078d, /* 1948 */
128'he0fff0efc632ec06006c842ee8221101, /* 1949 */
128'h4703c1a8081300002817468100c16583, /* 1950 */
128'h78930006460300f806330007079b0005, /* 1951 */
128'h61058536644260e2ec05000898630446, /* 1952 */
128'hf4e3fd07879b00088b63004678938082, /* 1953 */
128'hc6098a09b7d196be050502d586b3feb7, /* 1954 */
128'he008b7cdfc97879b0ff7f793fe07079b, /* 1955 */
128'h601cf87ff0ef842ee406e0221141b7e1, /* 1956 */
128'h00e6ea6302d704630007c70304b00693, /* 1957 */
128'h80820141640260a202d70e6304700693, /* 1958 */
128'hfed716e306b0069302d7076304d00693, /* 1959 */
128'hc683fce69fe3052a069007130017c683, /* 1960 */
128'hb7e9e01c078d00e69863042007130027, /* 1961 */
128'he406e0221141bfd50789bff1052a052a, /* 1962 */
128'hfff5c70300a405b395bff0efe589842a, /* 1963 */
128'h4703973efff58513b407879300002797, /* 1964 */
128'h80820141557d640260a2e7198b110007, /* 1965 */
128'h00074703973e00054703fea47ae3157d, /* 1966 */
128'h014105054581462960a26402f77d8b11, /* 1967 */
128'h00a107a31141fa5ff06f4581d7dff06f, /* 1968 */
128'h47818082014100e1550300a107238121, /* 1969 */
128'h069b8082853ee3190005470345a94625, /* 1970 */
128'h9fb902f587bb00d667630ff6f693fd07, /* 1971 */
128'h842ee406e0221141bff90505fd07879b, /* 1972 */
128'h02b455bb45a900b7f86347a500a04563, /* 1973 */
128'h60a2640202a4753b4529fe7ff0ef357d, /* 1974 */
128'h471707fe47854ac0006f030505130141, /* 1975 */
128'h808226f739230000471726f739230000, /* 1976 */
128'h862ee4262644041300004417e8221101, /* 1977 */
128'h60e2600ca2fff0efec06600885aa84ae, /* 1978 */
128'h479711418082610564a26442e00c95a6, /* 1979 */
128'h8793000047976380e022232787930000, /* 1980 */
128'h9d81e4068d45051300004517638c22e7, /* 1981 */
128'h014160a2640283220000100fba5fd0ef, /* 1982 */
128'h03638fefa0ef8432e406e02211418302, /* 1983 */
128'h8082450180820141640260a2557d0085, /* 1984 */
128'hf606852289aae64e01258413f2227169, /* 1985 */
128'h00a404b30505fe8ff0ef892eea4aee26, /* 1986 */
128'h071bee5ff0ef95260505fdcff0ef8526, /* 1987 */
128'haf230000479704e7ee631ff00793fff5, /* 1988 */
128'h05130000351784aafbaff0ef852218a7, /* 1989 */
128'h04a7f2630ff007939526facff0ef68e5, /* 1990 */
128'h6705051300003517842af9cff0ef8522, /* 1991 */
128'h838505130000451700a405b3f8eff0ef, /* 1992 */
128'h615569b2695264f2741270b2af5fd0ef, /* 1993 */
128'hb75514f7212300004717200007938082, /* 1994 */
128'h000035978cdff0ef850a458110000613, /* 1995 */
128'h079301294703e54ff0ef850a62c58593, /* 1996 */
128'h850a80a585930000459700f7096302f0, /* 1997 */
128'h00004797e5cff0ef850a85a2e64ff0ef, /* 1998 */
128'h7f05051300003517858a43900fc78793, /* 1999 */
128'h00004717451101f417934405a85fd0ef, /* 2000 */
128'hdefff0ef0ef73223000047170ef73223, /* 2001 */
128'h4797de1ff0ef4501eca7902300004797, /* 2002 */
128'hea858593000045974611eaa79a230000, /* 2003 */
128'hb7990a87932300004797eb1ff0ef854e, /* 2004 */
128'hdf638432478de04ae426ec06e8221101, /* 2005 */
128'h0004d783da3ff0ef84ae450d892a08c7, /* 2006 */
128'hf0ef076555030000451708a795632501, /* 2007 */
128'hffc4059b06a79a6325010024d783d8df, /* 2008 */
128'h4797d71ff0ef4511dfdff0ef00448513, /* 2009 */
128'hf0ef0465550300004517e4a791230000, /* 2010 */
128'h00004597e2a79723000047974611d5df, /* 2011 */
128'h256000ef4535e2dff0ef854ae2458593, /* 2012 */
128'h0513d6fff0ef451501c5d58300004597, /* 2013 */
128'hd7830067879300004797240000ef0200, /* 2014 */
128'h00004797fef71c230000471727850007, /* 2015 */
128'h000035170087cf63278d439cfec78793, /* 2016 */
128'h690264a260e26442971fd0ef6fc50513, /* 2017 */
128'h6105690264a2644260e2d9bff06f6105, /* 2018 */
128'h0fa347090105c783f022f40671798082, /* 2019 */
128'h8e6301e1578300f10f230115c78300f1, /* 2020 */
128'h0000351770a2740202e78a63470d00e7, /* 2021 */
128'h00003517842a91ffd06f61456dc50513, /* 2022 */
128'h65a27402852290ffd0efe42e6b450513, /* 2023 */
128'h05c170a241907402d8dff06f614570a2, /* 2024 */
128'h342322813823dc010113ebfff06f6145, /* 2025 */
128'h06134581893284ae842a232130232291, /* 2026 */
128'h061385a6eccff0ef22113c2300282180, /* 2027 */
128'h8522002cf0eff0efe802c44a08282040, /* 2028 */
128'h228134832301340323813083f63ff0ef, /* 2029 */
128'hd7830000479780822401011322013903, /* 2030 */
128'hf06fcea58593000045974611cb81f027, /* 2031 */
128'h1041e703474000efe40611418082cf5f, /* 2032 */
128'h10e1a02327051001a70300e57763878e, /* 2033 */
128'h91011782150260a21007e78310a7a223, /* 2034 */
128'he822ec06110180824501808201418d5d, /* 2035 */
128'h07933b0000ef842afc1ff0ef84aae426, /* 2036 */
128'hd533644260e29101150202f407b33e80, /* 2037 */
128'he022e40611418082610564a28d0502a7, /* 2038 */
128'h8793000f47b7384000ef842af95ff0ef, /* 2039 */
128'h014191011502640260a202f407b32407, /* 2040 */
128'he04ae426e822ec061101808202a7d533, /* 2041 */
128'h02a48533352000ef892af63ff0ef84aa, /* 2042 */
128'h0405944a0285543324040413000f4437, /* 2043 */
128'h690264a2644260e2fe856ee3f45ff0ef, /* 2044 */
128'hec06e822009894b7e426110180826105, /* 2045 */
128'h89260084f363892268048493842ae04a, /* 2046 */
128'h644260e2f47dfa1ff0ef41240433854a, /* 2047 */
128'h4503808200b5002380826105690264a2, /* 2048 */
128'h020575130147c503100007b780820005, /* 2049 */
128'hdfe50207f79301474783100007378082, /* 2050 */
128'h071300078223100007b7808200a70023, /* 2051 */
128'h0007822300e78023476d00e78623f800, /* 2052 */
128'h071300e78423fc70071300e78623470d, /* 2053 */
128'h842ae406e0221141808200e788230200, /* 2054 */
128'hf0ef80820141640260a2e50900044503, /* 2055 */
128'h7713ad27879300002797b7f50405fa5f, /* 2056 */
128'h0007c7830007470397aa973e811100f5, /* 2057 */
128'h002ce8221101808200f5802300e580a3, /* 2058 */
128'hf0ef00814503fd1ff0efec068121842a, /* 2059 */
128'h0ff47513002cf5dff0ef00914503f65f, /* 2060 */
128'h00914503f4bff0ef00814503fb7ff0ef, /* 2061 */
128'hf022717980826105644260e2f43ff0ef, /* 2062 */
128'h0089553b54e14461892af406e84aec26, /* 2063 */
128'h346100814503f81ff0ef0ff57513002c, /* 2064 */
128'hfe9410e3f0bff0ef00914503f13ff0ef, /* 2065 */
128'hf022717980826145694264e2740270a2, /* 2066 */
128'h553354e103800413892af406e84aec26, /* 2067 */
128'h00814503f3fff0ef0ff57513002c0089, /* 2068 */
128'h10e3ec9ff0ef00914503ed1ff0ef3461, /* 2069 */
128'h110180826145694264e2740270a2fe94, /* 2070 */
128'hea7ff0ef00814503f13ff0efec06002c, /* 2071 */
128'h100f8082610560e2e9fff0ef00914503, /* 2072 */
128'h9f858593000025974305f14025730000, /* 2073 */
128'h8593000035974605da0101138302037e, /* 2074 */
128'h382324113c23c56505130000451713e5, /* 2075 */
128'h2501ebbfa0ef25213023249134232481, /* 2076 */
128'h3083daafd0ef3865051300003517c115, /* 2077 */
128'h01132401390324813483250134032581, /* 2078 */
128'hd88fd0ef384505130000351780822601, /* 2079 */
128'hed3fa0ef080839658593000035974605, /* 2080 */
128'h0000391704e20bf00493ed2144012501, /* 2081 */
128'h95a66605007491810204159345490913, /* 2082 */
128'hde7ff0ef4521ed19250183afb0ef0808, /* 2083 */
128'hdd7ff0ef0007c50397ca8b8d00c4579b, /* 2084 */
128'h2501ceefb0ef54020808fbe19c3d47b2, /* 2085 */
128'h00003517bf8535e5051300003517c919, /* 2086 */
128'h07058593000035974605b79d33c50513, /* 2087 */
128'h051300003517c5112501e03fa0ef4501, /* 2088 */
128'h85a20184961386a20bf00493b7a134e5, /* 2089 */
128'h00003517cdcfd0ef3505051300003517, /* 2090 */
128'h90ef0184951385a2cd0fd0ef38c50513, /* 2091 */
128'h051300003517c981c62e0005059b9bef, /* 2092 */
128'hb705051300003517b721cb2fd0ef3865, /* 2093 */
128'h1141900200000023eabff0efca4fd0ef, /* 2094 */
128'h0513000f4537a001df9ff0efe4062501, /* 2095 */
128'haf870713000047178082450180822405, /* 2096 */
128'he30895360017869300756513157d631c, /* 2097 */
128'h110102b506338082953e055e10d00513, /* 2098 */
128'hc509842afd1ff0efe4328532ec06e822, /* 2099 */
128'h6105644260e28522a40ff0ef45816622, /* 2100 */
128'he4063225051300003517114180828082, /* 2101 */
128'h450160a2fe1fc0ef20000537c24fd0ef, /* 2102 */
128'hb0002573808245018082450180820141, /* 2103 */
128'h862e86b287361141808202f5553347a9, /* 2104 */
128'hbe8fd0efe40630e505130000351785aa, /* 2105 */
128'h952e842ae0221141a001d4bff0ef4505, /* 2106 */
128'h640260a29522408007b3f57ff0efe406, /* 2107 */
128'h45058082450580824505808201418d7d, /* 2108 */
128'h00c684bb842ef406ec26f02271798082, /* 2109 */
128'h80826145450164e2740270a200961863, /* 2110 */
128'h200404136622f33fc0efe432852285b2, /* 2111 */
128'h808245098082450980824509bff92605, /* 2112 */
128'hf06f8082450180824501808280828082, /* 2113 */
128'h003796934781e426e822ec061101c4bf, /* 2114 */
128'h644260e200c7986300d5043300d584b3, /* 2115 */
128'h036360980004380380826105450164a2, /* 2116 */
128'hd0ef28250513000035176090600c02e8, /* 2117 */
128'hd0ef29a505130000351785a28626b26f, /* 2118 */
128'h3517892ae0ca711dbf5d0785a001b16f, /* 2119 */
128'hf05af456f852fc4ee8a229a505130000, /* 2120 */
128'hd0ef44018b2ee466e4a6ec86e862ec5e, /* 2121 */
128'h8b9300003b97286a0a1300003a17ae6f, /* 2122 */
128'h4ac1292c0c1300003c17fff9499328eb, /* 2123 */
128'hd0ef855e85e600040c9bac2fd0ef8552, /* 2124 */
128'haa8fd0ef855203649863448187caab6f, /* 2125 */
128'h02b49b63458187caaa0fd0ef856285e6, /* 2126 */
128'hd0ef2ba5051300003517fd5417e30405, /* 2127 */
128'hc689873e8a85008486b3a8894501a86f, /* 2128 */
128'h07a104856398e39840e9873300349713, /* 2129 */
128'h9713c689873e8a856390008586b3bf5d, /* 2130 */
128'h00003517058e02e60d6340e987330035, /* 2131 */
128'h2485051300003517a40fd0ef21c50513, /* 2132 */
128'h79e2690664a6644660e6557da34fd0ef, /* 2133 */
128'h808261256ca26c426be27b027aa27a42, /* 2134 */
128'h8aaa6a05fc56e0d27159bfa507a10585, /* 2135 */
128'hf486f062f45ef85ae4ceeca602000513, /* 2136 */
128'h44818bb28b2ee46ee86aec66e8caf0a2, /* 2137 */
128'h0c1300003c179c4a0a134981bcfff0ef, /* 2138 */
128'h9b6300fb0cb300fa8db3003497934aec, /* 2139 */
128'h74069bafd0ef21650513000035170374, /* 2140 */
128'h6d426ce27c027ba26a0669a6694670a6, /* 2141 */
128'h61657ae285567b4264e685da86266da2, /* 2142 */
128'h8d2acd3fe0ef842acd9fe0efe33ff06f, /* 2143 */
128'h151b0344f7b3cc7fe0ef892accdfe0ef, /* 2144 */
128'h150201a4643300a96533010d1d1b0105, /* 2145 */
128'hef8100adb02300acb0238d4191011402, /* 2146 */
128'hc50397e20039f7930985b3dff0ef4521, /* 2147 */
128'he032e42e7139b7ad0485b2dff0ef0007, /* 2148 */
128'hc71fe0ef89aaec4ef04af426f822fc06, /* 2149 */
128'he0ef84aac65fe0ef892ac6bfe0ef842a, /* 2150 */
128'h15028fc18d450109179b0105151bc5ff, /* 2151 */
128'h0037971347818d5d9101178265a26602, /* 2152 */
128'h74a270e2744200c79c63974e00e58833, /* 2153 */
128'h6314d79ff06f6121863e69e2854e7902, /* 2154 */
128'h00e830238f2900083703e3148ea90785, /* 2155 */
128'hf04af426f822fc06e032e42e7139b7f1, /* 2156 */
128'h892abf3fe0ef842abf9fe0ef89aaec4e, /* 2157 */
128'h179b0105151bbe7fe0ef84aabedfe0ef, /* 2158 */
128'h9101178265a2660215028fc18d450109, /* 2159 */
128'h9c63974e00e588330037971347818d5d, /* 2160 */
128'h863e69e2854e790274a270e2744200c7, /* 2161 */
128'h3703e3148e8907856314d01ff06f6121, /* 2162 */
128'he032e42e7139b7f100e830238f090008, /* 2163 */
128'hb81fe0ef89aaec4ef04af426f822fc06, /* 2164 */
128'he0ef84aab75fe0ef892ab7bfe0ef842a, /* 2165 */
128'h15028fc18d450109179b0105151bb6ff, /* 2166 */
128'h0037971347818d5d9101178265a26602, /* 2167 */
128'h74a270e2744200c79c63974e00e58833, /* 2168 */
128'h6314c89ff06f6121863e69e2854e7902, /* 2169 */
128'h02a7073300083703e31402a686b30785, /* 2170 */
128'hf822fc06e032e42e7139b7e100e83023, /* 2171 */
128'he0ef842ab05fe0ef89aaec4ef04af426, /* 2172 */
128'h151baf3fe0ef84aaaf9fe0ef892aafff, /* 2173 */
128'h65a2660215028fc18d450109179b0105, /* 2174 */
128'h00e588330037971347818d5d91011782, /* 2175 */
128'h854e790274a270e2744200c79c63974e, /* 2176 */
128'h63144505e111c0dff06f6121863e69e2, /* 2177 */
128'h02a7573300083703e31402a6d6b30785, /* 2178 */
128'hf822fc06e032e42e7139b7d100e83023, /* 2179 */
128'he0ef842aa85fe0ef89aaec4ef04af426, /* 2180 */
128'h151ba73fe0ef84aaa79fe0ef892aa7ff, /* 2181 */
128'h65a2660215028fc18d450109179b0105, /* 2182 */
128'h00e588330037971347818d5d91011782, /* 2183 */
128'h854e790274a270e2744200c79c63974e, /* 2184 */
128'h8ec907856314b8dff06f6121863e69e2, /* 2185 */
128'h7139b7f100e830238f4900083703e314, /* 2186 */
128'h89aaec4ef04af426f822fc06e032e42e, /* 2187 */
128'ha01fe0ef892aa07fe0ef842aa0dfe0ef, /* 2188 */
128'h8d450109179b0105151b9fbfe0ef84aa, /* 2189 */
128'h47818d5d9101178265a2660215028fc1, /* 2190 */
128'h744200c79c63974e00e5883300379713, /* 2191 */
128'hf06f6121863e69e2854e790274a270e2, /* 2192 */
128'h8f6900083703e3148ee907856314b15f, /* 2193 */
128'hf822fc06e032e42e7139b7f100e83023, /* 2194 */
128'he0ef842a995fe0ef89aaec4ef04af426, /* 2195 */
128'h151b983fe0ef84aa989fe0ef892a98ff, /* 2196 */
128'h65a2660214828fc18cc90109179b0105, /* 2197 */
128'h00d988330037169347018fc590811782, /* 2198 */
128'h854e790274a270e2744200c71c6396ae, /* 2199 */
128'he28800f70533a9dff06f6121863a69e2, /* 2200 */
128'h3517892ae8ca7159bfc9070500a83023, /* 2201 */
128'hf85afc56e0d2e4cef0a2d7a505130000, /* 2202 */
128'h44018b3289aeec66eca6f486f062f45e, /* 2203 */
128'h00003b97d64a0a1300003a17dc5fc0ef, /* 2204 */
128'h04000a93d74c0c1300003c17d6cb8b93, /* 2205 */
128'h8885855e85a2fff44493da3fc0ef8552, /* 2206 */
128'h0036179314fd460140900cb3d95fc0ef, /* 2207 */
128'hc0efe43285520566186397ce00f905b3, /* 2208 */
128'h854a85ce6622d6ffc0ef856285a2d77f, /* 2209 */
128'h3517fb541be32405e12984aaa03ff0ef, /* 2210 */
128'h8526740670a6d4ffc0efd82505130000, /* 2211 */
128'h7c027ba27b427ae26a0669a664e66946, /* 2212 */
128'h8726c291876600167693808261656ce2, /* 2213 */
128'heca67159bfc154fdbf590605e198e398, /* 2214 */
128'he4cee8caf0a2ca6505130000351784aa, /* 2215 */
128'he86af486ec66f062f45ef85afc56e0d2, /* 2216 */
128'h899300003997ceffc0ef44018ab2892e, /* 2217 */
128'h8b9300003b97ef6b0b1300003b17c8e9, /* 2218 */
128'h8c9300003c97c86c0c1300003c17ef6b, /* 2219 */
128'h00147793cbdfc0ef854e04000a13c8ec, /* 2220 */
128'h4601cabfc0ef856285a2000bbd03cba5, /* 2221 */
128'h1c6397ca00f485b300361793fffd4513, /* 2222 */
128'hc0ef856685a2c8ffc0efe432854e0556, /* 2223 */
128'he5298d2a91bff0ef852685ca6622c87f, /* 2224 */
128'hc0efc9a5051300003517fb441ae32405, /* 2225 */
128'h6a0669a6694664e6856a740670a6c67f, /* 2226 */
128'h808261656d426ce27c027ba27b427ae2, /* 2227 */
128'h872ac291876a00167693bf49000b3d03, /* 2228 */
128'he8a2711db7e15d7db7790605e198e398, /* 2229 */
128'hf852e0cae4a6bb65051300003517842a, /* 2230 */
128'h8ab284aefc4eec86e862ec5ef05af456, /* 2231 */
128'h3b17ba29091300003917c03fc0ef4c01, /* 2232 */
128'h0a13bb2b8b9300003b97baab0b130000, /* 2233 */
128'h855a85ce000c099bbe1fc0ef854a1000, /* 2234 */
128'he7b38fd9010c1793008c1713bd5fc0ef, /* 2235 */
128'h17138fd9020c17138fd9018c17130187, /* 2236 */
128'h8fd9038c17138fd9030c17138fd9028c, /* 2237 */
128'h05561763972600e406b3003617134601, /* 2238 */
128'hb89fc0ef855e85ceb91fc0efe432854a, /* 2239 */
128'h0c05e91d89aa81dff0ef852285a66622, /* 2240 */
128'hb69fc0efb9c5051300003517f94c19e3, /* 2241 */
128'h7aa27a4279e2690664a6854e644660e6, /* 2242 */
128'h0605e29ce31c808261256c426be27b02, /* 2243 */
128'h0000351784aaf4a67119bff159fdb74d, /* 2244 */
128'he0dae4d6e8d2eccef0caf8a2acc50513, /* 2245 */
128'h8b32892eec6efc86f06af466f862fc5e, /* 2246 */
128'h3c97ab2a0a1300003a17b13fc0ef4401, /* 2247 */
128'h03f00c13498507f00b93abac8c930000, /* 2248 */
128'hc0ef855208000a93ab8d0d1300003d17, /* 2249 */
128'h9733408b873badffc0ef856685a2ae7f, /* 2250 */
128'h00f486b3003617934601008995b300e9, /* 2251 */
128'h85a2abbfc0efe432855205661a6397ca, /* 2252 */
128'hf46ff0ef852685ca6622ab3fc0ef856a, /* 2253 */
128'h051300003517fb541be32405e1398daa, /* 2254 */
128'h790674a6856e744670e6a93fc0efac65, /* 2255 */
128'h7d027ca27c427be26b066aa66a4669e6, /* 2256 */
128'h0605e28ce38c008c6663808261096de2, /* 2257 */
128'hf4a67119b7f15dfdbfe5e298e398bf61, /* 2258 */
128'heccef0caf8a29e6505130000351784aa, /* 2259 */
128'hfc86f06af466f862fc5ee0dae4d6e8d2, /* 2260 */
128'h00003a17a2dfc0ef44018b32892eec6e, /* 2261 */
128'h07f00b939d4c8c9300003c979cca0a13, /* 2262 */
128'h0a939d2d0d1300003d1703f00c134985, /* 2263 */
128'h9f9fc0ef856685a2a01fc0ef85520800, /* 2264 */
128'hfff7c793008996b300f997b3408b87bb, /* 2265 */
128'h974a00e485b3003617134601fff6c693, /* 2266 */
128'h856a85a29cdfc0efe432855205661a63, /* 2267 */
128'h8daae58ff0ef852685ca66229c5fc0ef, /* 2268 */
128'h9d85051300003517fb5417e32405e139, /* 2269 */
128'h69e6790674a6856e744670e69a5fc0ef, /* 2270 */
128'h6de27d027ca27c427be26b066aa66a46, /* 2271 */
128'hbf610605e194e314008c666380826109, /* 2272 */
128'h84aaf4a67119b7f15dfdbfe5e19ce31c, /* 2273 */
128'he8d2eccef0caf8a28f85051300003517, /* 2274 */
128'hec6efc86f06af466f862fc5ee0dae4d6, /* 2275 */
128'h89930000399793ffc0ef44018a32892e, /* 2276 */
128'h4d0507f00a938e6c0c1300003c178de9, /* 2277 */
128'h8e0c8c9300003c9703f00b9308100b13, /* 2278 */
128'h873b90bfc0ef856285a2913fc0ef854e, /* 2279 */
128'h8f5d00ed173300fd17b3408b07bb408a, /* 2280 */
128'h48938fd5008d16b300fd17b30024079b, /* 2281 */
128'h00d48533003616934601fff7c313fff7, /* 2282 */
128'h85a28cbfc0efe432854e05461c6396ca, /* 2283 */
128'hd56ff0ef852685ca66228c3fc0ef8566, /* 2284 */
128'h3517f8f41be3080007932405ed298daa, /* 2285 */
128'h856e744670e689ffc0ef8d2505130000, /* 2286 */
128'h7c427be26b066aa66a4669e6790674a6, /* 2287 */
128'hea6300167813808261096de27d027ca2, /* 2288 */
128'h0605e10ce28c85be00081363859a008b, /* 2289 */
128'hbf755dfdbfc585bafe081be385c6b761, /* 2290 */
128'hecce7e25051300002517892af0ca7119, /* 2291 */
128'hf4a6f8a2fc86ec6ef06af466fc5ee8d2, /* 2292 */
128'h829fc0ef4b81e03289aef862e0dae4d6, /* 2293 */
128'h7d0c8c9300002c977c8a0a1300002a17, /* 2294 */
128'h01779c3347854da17d8d0d1300002d17, /* 2295 */
128'h00848b3bffcfc0ef85524401003b949b, /* 2296 */
128'h67824601fffc4a93ff0fc0ef856685da, /* 2297 */
128'h855206f61063974e00e9083300361713, /* 2298 */
128'h6622fcafc0ef856a85dafd2fc0efe432, /* 2299 */
128'h8c562405e9318b2ac5eff0ef854a85ce, /* 2300 */
128'h2517fafb90e3040007932b85fbb41be3, /* 2301 */
128'h855a744670e6f9efc0ef7d2505130000, /* 2302 */
128'h7c427be26b066aa66a4669e6790674a6, /* 2303 */
128'h85e200167513808261096de27d027ca2, /* 2304 */
128'h5b7db749060500b83023e30c85d6e111, /* 2305 */
128'h0513892e84aaf4cef8cafca67175b7e9, /* 2306 */
128'hfc66e0e2e4dee8daecd6f0d269850200, /* 2307 */
128'h922ff0ef4a81e032f46ef86ae122e506, /* 2308 */
128'h3c979c498993006c0c1300004c174a01, /* 2309 */
128'h67824d214d818bca8b269fac8c930000, /* 2310 */
128'h852685ca866e04fd956396da003d9693, /* 2311 */
128'h00002517020a0863ed45842aba2ff0ef, /* 2312 */
128'h74e6640a60aa8522ef0fc0ef74c50513, /* 2313 */
128'h7ce26c066ba66b466ae67a0679a67946, /* 2314 */
128'hb7758ba68b4a4a05808261497da27d42, /* 2315 */
128'he0efe82aa04fe0ef842aa0afe0efec36, /* 2316 */
128'h0105151b664267a29f8fe0efe42a9fef, /* 2317 */
128'h66e29101140215028c510106161b8d5d, /* 2318 */
128'h86b34781e288f6a7b323000047978d41, /* 2319 */
128'h0ff6f693078500fb86330006c6830187, /* 2320 */
128'hef910ba1033df7b3ffa795e300d60023, /* 2321 */
128'h8b8d00078a9b001a879b84cff0ef4521, /* 2322 */
128'h547dbf0d0d85838ff0ef0007c50397e6, /* 2323 */
128'h051389ae892af0d2f4cef8ca7175bfa1, /* 2324 */
128'hfc66e0e2e4dee8daecd6fca66a050200, /* 2325 */
128'h802ff0ef4b018cb2f46ee122e506f86a, /* 2326 */
128'h3d179c4a0a13eee48493000044974a81, /* 2327 */
128'h003d97934d818c4e8bca8dad0d130000, /* 2328 */
128'h854a85ce866e059d956397de00fc06b3, /* 2329 */
128'h00002517020a8863e579842aa82ff0ef, /* 2330 */
128'h74e6640a60aa8522dd0fc0ef62c50513, /* 2331 */
128'h7ce26c066ba66b466ae67a0679a67946, /* 2332 */
128'hb7758c4a8bce4a85808261497da27d42, /* 2333 */
128'he42a8e2fe0ef842a8e8fe0efe836ec3e, /* 2334 */
128'h151b670266228d6fe0efe02a8dcfe0ef, /* 2335 */
128'h9101140215028c518d590106161b0105, /* 2336 */
128'he38866c267e2e4a7b723000047978d41, /* 2337 */
128'h0024d78300f6902393c117c20004d783, /* 2338 */
128'h93c117c20044d78300f6912393c117c2, /* 2339 */
128'h00f6932393c117c20064d78300f69223, /* 2340 */
128'h001b079bf17fe0ef4521ef91034df7b3, /* 2341 */
128'hf03fe0ef0007c50397ea8b8d00078b1b, /* 2342 */
128'hf8ca717580826505b789547dbf290d85, /* 2343 */
128'h962a84ae842afca6e122fff586138932, /* 2344 */
128'hecd6f0d2f4ce54e505130000251785aa, /* 2345 */
128'hec36e506f46ef86afc66e0e2e4dee8da, /* 2346 */
128'hd793e83e0014d9930044d793cd4fc0ef, /* 2347 */
128'h0b1300002b1744854a81e43e99a20034, /* 2348 */
128'h0c1300002c17536b8b9300002b97536b, /* 2349 */
128'h0d1300002d17536c8c9300002c97536c, /* 2350 */
128'h0a1300004a1753ed8d9300002d9753ed, /* 2351 */
128'hc0ef532505130000251702997863d46a, /* 2352 */
128'h7a0679a6794674e68556640a60aac76f, /* 2353 */
128'h61497da27d427ce26c066ba66b466ae6, /* 2354 */
128'h85ca00090663c4efc0ef855a85a68082, /* 2355 */
128'h856a85e6c3cfc0ef8562c42fc0ef855e, /* 2356 */
128'h856eed15920ff0ef852265a2c34fc0ef, /* 2357 */
128'h358302f749636762010a2783c24fc0ef, /* 2358 */
128'hc08fc0ef4b45051300002517c58d000a, /* 2359 */
128'h000025179782852285ce6642008a3783, /* 2360 */
128'h00002517b7e94a89bf0fc0ef4a450513, /* 2361 */
128'h25177179bfa10485be0fc0ef1d450513, /* 2362 */
128'he44ee84aec26f022f406492505130000, /* 2363 */
128'h490505130000251704000593ca9fe0ef, /* 2364 */
128'hba8fc0ef4ac5051300002517bb4fc0ef, /* 2365 */
128'h00002517b9cfc0ef4d05051300002517, /* 2366 */
128'h01f499934441b8efc0ef448518450513, /* 2367 */
128'h24050135853346054685008495b34979, /* 2368 */
128'h694264e2740270a2ff2417e3e6dff0ef, /* 2369 */
128'h00c51f1b02a3033b430d8082614569a2, /* 2370 */
128'h462946814e8147010015181b0025189b, /* 2371 */
128'h802340000e13c2678793000047974585, /* 2372 */
128'h802301078fb3000f802300a78fb30007, /* 2373 */
128'h10e397c63e7d000f802300678fb3000f, /* 2374 */
128'h26f38e15c020267302c71d632705fe0e, /* 2375 */
128'h059302a6873341d686b33e800513c000, /* 2376 */
128'h473302a767b302bf45bb02c747334000, /* 2377 */
128'h1ae3adafc06f456505130000251702a7, /* 2378 */
128'he4061141b761c0002ef3c02026f3f8b7, /* 2379 */
128'hf0ef4509f5fff0ef4505f65ff0ef4501, /* 2380 */
128'h4541f4dff0ef4521f53ff0ef4511f59f, /* 2381 */
128'he06f4825051300002517bff1f47ff0ef, /* 2382 */
128'he0efe4064780e022400007b71141b7bf, /* 2383 */
128'h2401b5ffe0ef43e5051300002517b39f, /* 2384 */
128'h579ba6afc0ef43e505130000251785a2, /* 2385 */
128'h8e634709cb8100e78e63470527810064, /* 2386 */
128'hc69fe0ef8522a00100e78f63470d00e7, /* 2387 */
128'h83df80ef8522bfc5e69ff0ef8522bfe5, /* 2388 */
128'h000000000000b7c5f69ff0ef8522b7e5, /* 2389 */
128'h00000000000000000000000000000000, /* 2390 */
128'h00000000000000000000000000000000, /* 2391 */
128'h00000000000000000000000000000000, /* 2392 */
128'h00000000000000000000000000000000, /* 2393 */
128'h00000000000000000000000000000000, /* 2394 */
128'h00000000000000000000000000000000, /* 2395 */
128'h00000000000000000000000000000000, /* 2396 */
128'h00000000000000000000000000000000, /* 2397 */
128'h00000000000000000000000000000000, /* 2398 */
128'h00000000000000000000000000000000, /* 2399 */
128'h08082828282828080808080808080808, /* 2400 */
128'h08080808080808080808080808080808, /* 2401 */
128'h101010101010101010101010101010a0, /* 2402 */
128'h10101010101004040404040404040404, /* 2403 */
128'h01010101010101010141414141414110, /* 2404 */
128'h10101010100101010101010101010101, /* 2405 */
128'h02020202020202020242424242424210, /* 2406 */
128'h08101010100202020202020202020202, /* 2407 */
128'h00000000000000000000000000000000, /* 2408 */
128'h00000000000000000000000000000000, /* 2409 */
128'h101010101010101010101010101010a0, /* 2410 */
128'h10101010101010101010101010101010, /* 2411 */
128'h01010101010101010101010101010101, /* 2412 */
128'h02010101010101011001010101010101, /* 2413 */
128'h02020202020202020202020202020202, /* 2414 */
128'h02020202020202021002020202020202, /* 2415 */
128'hc1bdceee242070dbe8c7b756d76aa478, /* 2416 */
128'hfd469501a83046134787c62af57c0faf, /* 2417 */
128'h895cd7beffff5bb18b44f7af698098d8, /* 2418 */
128'h49b40821a679438efd9871936b901122, /* 2419 */
128'he9b6c7aa265e5a51c040b340f61e2562, /* 2420 */
128'he7d3fbc8d8a1e68102441453d62f105d, /* 2421 */
128'h455a14edf4d50d87c33707d621e1cde6, /* 2422 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /* 2423 */
128'hfde5380c6d9d61228771f681fffa3942, /* 2424 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /* 2425 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /* 2426 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /* 2427 */
128'hfc93a039ab9423a7432aff97f4292244, /* 2428 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /* 2429 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /* 2430 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /* 2431 */
128'h0c07020d08030e09040f0a05000b0601, /* 2432 */
128'h020f0c090603000d0a0704010e0b0805, /* 2433 */
128'h09020b040d060f08010a030c050e0700, /* 2434 */
128'h6c5f7465735f64735f63736972776f6c, /* 2435 */
128'h6e67696c615f64730000000000006465, /* 2436 */
128'h645f6b6c635f64730000000000000000, /* 2437 */
128'h69747465735f64730000000000007669, /* 2438 */
128'h735f646d635f6473000000000000676e, /* 2439 */
128'h74657365725f64730000000074726174, /* 2440 */
128'h6e636b6c625f64730000000000000000, /* 2441 */
128'h69736b6c625f64730000000000000074, /* 2442 */
128'h6f656d69745f6473000000000000657a, /* 2443 */
128'h655f7172695f64730000000000007475, /* 2444 */
128'h5f63736972776f6c000000000000006e, /* 2445 */
128'h00000000646d635f74726174735f6473, /* 2446 */
128'h746e695f746961775f63736972776f6c, /* 2447 */
128'h000000000067616c665f747075727265, /* 2448 */
128'h00007172695f64735f63736972776f6c, /* 2449 */
128'h695f646d635f64735f63736972776f6c, /* 2450 */
128'h5f63736972776f6c0000000000007172, /* 2451 */
128'h007172695f646e655f617461645f6473, /* 2452 */
128'h0000000087fe99880000000087feb040, /* 2453 */
128'h004c4b40004c4b400030000020000000, /* 2454 */
128'h6d6d5f6472616f62000000020000ffff, /* 2455 */
128'h0000000087fe4e880064637465675f63, /* 2456 */
128'h0000000087fe4cf40000000087fe4a96, /* 2457 */
128'h00000000000000000000000000000000, /* 2458 */
128'hffffbe6affffbe66ffffbe66ffffbe40, /* 2459 */
128'hffffbe6effffbe6effffbe6effffbe6e, /* 2460 */
128'h0000000087feb3680000000087feb358, /* 2461 */
128'h0000000087feb3900000000087feb378, /* 2462 */
128'h0000000087feb3c00000000087feb3a8, /* 2463 */
128'h0000000087feb3f00000000087feb3d8, /* 2464 */
128'h0000000087feb4200000000087feb408, /* 2465 */
128'h0000000087feb4500000000087feb438, /* 2466 */
128'h40040300400402004004010040040000, /* 2467 */
128'h40050000400405004004040140040400, /* 2468 */
128'h30000000000000030000000040050100, /* 2469 */
128'h60000000000000053000000000000001, /* 2470 */
128'h70000000000000027000000000000004, /* 2471 */
128'h00000001400000007000000000000000, /* 2472 */
128'h00000005000000012000000000000006, /* 2473 */
128'h20000000000000020000000040000000, /* 2474 */
128'h00000000100000000000000100000000, /* 2475 */
128'h1e19140f0d0c0a000000000000000000, /* 2476 */
128'h000186a00000271050463c37322d2823, /* 2477 */
128'h017d7840017d784000989680000f4240, /* 2478 */
128'h031975000319750002faf080018cba80, /* 2479 */
128'h02faf08005f5e10002faf080017d7840, /* 2480 */
128'h00000020000000000bebc2000c65d400, /* 2481 */
128'h00000200000001000000008000000040, /* 2482 */
128'h00002000000010000000080000000400, /* 2483 */
128'h0000c000000080000000600000004000, /* 2484 */
128'h37363534333231300002000000010000, /* 2485 */
128'h2043534952776f4c4645444342413938, /* 2486 */
128'h746f6f622d7520646573696d696e696d, /* 2487 */
128'h00000000647261432d445320726f6620, /* 2488 */
128'h3809000038000000100c0000edfe0dd0, /* 2489 */
128'h00000000100000001100000028000000, /* 2490 */
128'h000000000000000000090000d8020000, /* 2491 */
128'h00000000010000000000000000000000, /* 2492 */
128'h02000000000000000400000003000000, /* 2493 */
128'h020000000f0000000400000003000000, /* 2494 */
128'h2c6874651b0000001400000003000000, /* 2495 */
128'h007665642d657261622d656e61697261, /* 2496 */
128'h2c687465260000001000000003000000, /* 2497 */
128'h0100000000657261622d656e61697261, /* 2498 */
128'h1a0000000300000000006e65736f6863, /* 2499 */
128'h303140747261752f636f732f2c000000, /* 2500 */
128'h0000003030323531313a303030303030, /* 2501 */
128'h00000000737570630100000002000000, /* 2502 */
128'h01000000000000000400000003000000, /* 2503 */
128'h000000000f0000000400000003000000, /* 2504 */
128'h40787d01380000000400000003000000, /* 2505 */
128'h03000000000000304075706301000000, /* 2506 */
128'h0300000080f0fa024b00000004000000, /* 2507 */
128'h03000000007570635b00000004000000, /* 2508 */
128'h03000000000000006700000004000000, /* 2509 */
128'h0000000079616b6f6b00000005000000, /* 2510 */
128'h7a6874651b0000001300000003000000, /* 2511 */
128'h0000766373697200656e61697261202c, /* 2512 */
128'h34367672720000000b00000003000000, /* 2513 */
128'h0b000000030000000000636466616d69, /* 2514 */
128'h0000393376732c76637369727c000000, /* 2515 */
128'h01000000850000000000000003000000, /* 2516 */
128'h6f72746e6f632d747075727265746e69, /* 2517 */
128'h04000000030000000000000072656c6c, /* 2518 */
128'h0000000003000000010000008f000000, /* 2519 */
128'h1b0000000f00000003000000a0000000, /* 2520 */
128'h000063746e692d7570632c7663736972, /* 2521 */
128'h02000000b50000000400000003000000, /* 2522 */
128'h02000000bb0000000400000003000000, /* 2523 */
128'h01000000020000000200000002000000, /* 2524 */
128'h0030303030303030384079726f6d656d, /* 2525 */
128'h6f6d656d5b0000000700000003000000, /* 2526 */
128'h67000000100000000300000000007972, /* 2527 */
128'h00000040000000000000008000000000, /* 2528 */
128'h000000007364656c0100000002000000, /* 2529 */
128'h6f6970671b0000000a00000003000000, /* 2530 */
128'h72616568010000000000007364656c2d, /* 2531 */
128'h0300000000000064656c2d7461656274, /* 2532 */
128'h0100000001000000c30000000c000000, /* 2533 */
128'hc90000000a0000000300000000000000, /* 2534 */
128'h03000000000000746165627472616568, /* 2535 */
128'h0200000002000000df00000000000000, /* 2536 */
128'h040000000300000000636f7301000000, /* 2537 */
128'h04000000030000000200000000000000, /* 2538 */
128'h1f00000003000000020000000f000000, /* 2539 */
128'h622d656e616972612c6874651b000000, /* 2540 */
128'h622d656c706d697300636f732d657261, /* 2541 */
128'hf6000000000000000300000000007375, /* 2542 */
128'h30303030303240746e696c6301000000, /* 2543 */
128'h1b0000000d0000000300000000000030, /* 2544 */
128'h0000000030746e696c632c7663736972, /* 2545 */
128'h02000000fd0000001000000003000000, /* 2546 */
128'h03000000070000000200000003000000, /* 2547 */
128'h00000002000000006700000010000000, /* 2548 */
128'h080000000300000000000c0000000000, /* 2549 */
128'h02000000006c6f72746e6f6311010000, /* 2550 */
128'h6f632d747075727265746e6901000000, /* 2551 */
128'h303030303030634072656c6c6f72746e, /* 2552 */
128'h00000000040000000300000000000000, /* 2553 */
128'h8f000000040000000300000000000000, /* 2554 */
128'h1b0000000c0000000300000001000000, /* 2555 */
128'h03000000003063696c702c7663736972, /* 2556 */
128'h1000000003000000a000000000000000, /* 2557 */
128'h020000000b00000002000000fd000000, /* 2558 */
128'h67000000100000000300000009000000, /* 2559 */
128'h00000004000000000000000c00000000, /* 2560 */
128'h070000001b0100000400000003000000, /* 2561 */
128'h030000002e0100000400000003000000, /* 2562 */
128'h03000000b50000000400000003000000, /* 2563 */
128'h03000000bb0000000400000003000000, /* 2564 */
128'h6f632d67756265640100000002000000, /* 2565 */
128'h030000000000304072656c6c6f72746e, /* 2566 */
128'h65642c76637369721b00000010000000, /* 2567 */
128'h0800000003000000003331302d677562, /* 2568 */
128'h03000000ffff000002000000fd000000, /* 2569 */
128'h00000000000000006700000010000000, /* 2570 */
128'h08000000030000000010000000000000, /* 2571 */
128'h02000000006c6f72746e6f6311010000, /* 2572 */
128'h30303030303031407472617501000000, /* 2573 */
128'h1b000000080000000300000000000030, /* 2574 */
128'h1000000003000000003035373631736e, /* 2575 */
128'h00000000000000100000000067000000, /* 2576 */
128'h4b000000040000000300000000100000, /* 2577 */
128'h39010000040000000300000080f0fa02, /* 2578 */
128'h47010000040000000300000000c20100, /* 2579 */
128'h58010000040000000300000003000000, /* 2580 */
128'h63010000040000000300000001000000, /* 2581 */
128'h6d010000040000000300000002000000, /* 2582 */
128'h2d737078010000000200000004000000, /* 2583 */
128'h00000000303030303030303240697073, /* 2584 */
128'h786e6c781b0000002800000003000000, /* 2585 */
128'h00622e30302e322d6970732d7370782c, /* 2586 */
128'h302e322d6970732d7370782c786e6c78, /* 2587 */
128'h00000000040000000300000000612e30, /* 2588 */
128'h0f000000040000000300000001000000, /* 2589 */
128'h47010000040000000300000000000000, /* 2590 */
128'h58010000080000000300000003000000, /* 2591 */
128'h10000000030000000200000002000000, /* 2592 */
128'h00000000000000200000000067000000, /* 2593 */
128'h7a010000080000000300000000100000, /* 2594 */
128'h040000000300000000377865746e696b, /* 2595 */
128'h04000000030000000100000086010000, /* 2596 */
128'h04000000030000000100000096010000, /* 2597 */
128'h040000000300000008000000a7010000, /* 2598 */
128'h40636d6d0100000004000000be010000, /* 2599 */
128'h1b0000000d0000000300000000000030, /* 2600 */
128'h00000000746f6c732d6970732d636d6d, /* 2601 */
128'h00000000670000000400000003000000, /* 2602 */
128'h20bcbe00cd0100000400000003000000, /* 2603 */
128'he40c0000df0100000800000003000000, /* 2604 */
128'hee0100000000000003000000e40c0000, /* 2605 */
128'h72776f6c010000000200000002000000, /* 2606 */
128'h3030303030303033406874652d637369, /* 2607 */
128'h1b0000000c0000000300000000000000, /* 2608 */
128'h03000000006874652d63736972776f6c, /* 2609 */
128'h006b726f7774656e5b00000008000000, /* 2610 */
128'h03000000470100000400000003000000, /* 2611 */
128'h03000000580100000800000003000000, /* 2612 */
128'hf9010000060000000300000000000000, /* 2613 */
128'h100000000300000000007fe3023e1800, /* 2614 */
128'h00000000000000300000000067000000, /* 2615 */
128'h6f697067010000000200000000800000, /* 2616 */
128'h03000000000000303030303030303440, /* 2617 */
128'h03000000020000000b02000004000000, /* 2618 */
128'h7370782c786e6c781b00000015000000, /* 2619 */
128'h00000000612e30302e312d6f6970672d, /* 2620 */
128'h03000000170200000000000003000000, /* 2621 */
128'h00000040000000006700000010000000, /* 2622 */
128'h04000000030000000000010000000000, /* 2623 */
128'h04000000030000000000000027020000, /* 2624 */
128'h04000000030000000000000037020000, /* 2625 */
128'h04000000030000000000000049020000, /* 2626 */
128'h0400000003000000000000005b020000, /* 2627 */
128'h0400000003000000080000006f020000, /* 2628 */
128'h0400000003000000080000007f020000, /* 2629 */
128'h04000000030000000000000090020000, /* 2630 */
128'h040000000300000001000000a7020000, /* 2631 */
128'h0400000003000000ffffffffb4020000, /* 2632 */
128'h0400000003000000ffffffffc5020000, /* 2633 */
128'h040000000300000001000000b5000000, /* 2634 */
128'h020000000200000001000000bb000000, /* 2635 */
128'h73736572646461230900000002000000, /* 2636 */
128'h6c65632d657a69732300736c6c65632d, /* 2637 */
128'h6f6d00656c62697461706d6f6300736c, /* 2638 */
128'h00687461702d74756f647473006c6564, /* 2639 */
128'h6e6575716572662d65736162656d6974, /* 2640 */
128'h6e6575716572662d6b636f6c63007963, /* 2641 */
128'h7200657079745f656369766564007963, /* 2642 */
128'h2c766373697200737574617473006765, /* 2643 */
128'h626c7400657079742d756d6d00617369, /* 2644 */
128'h7075727265746e69230074696c70732d, /* 2645 */
128'h7075727265746e6900736c6c65632d74, /* 2646 */
128'h6e696c0072656c6c6f72746e6f632d74, /* 2647 */
128'h736f69706700656c646e6168702c7875, /* 2648 */
128'h742d746c75616665642c78756e696c00, /* 2649 */
128'h74732d6e696174657200726567676972, /* 2650 */
128'h6172006465646e65707375732d657461, /* 2651 */
128'h2d73747075727265746e69007365676e, /* 2652 */
128'h6d616e2d676572006465646e65747865, /* 2653 */
128'h6972702d78616d2c7663736972007365, /* 2654 */
128'h7665646e2c766373697200797469726f, /* 2655 */
128'h690064656570732d746e657272756300, /* 2656 */
128'h00746e657261702d747075727265746e, /* 2657 */
128'h732d6765720073747075727265746e69, /* 2658 */
128'h746469772d6f692d6765720074666968, /* 2659 */
128'h6c7800796c696d61662c786e6c780068, /* 2660 */
128'h6c780074736978652d6f6669662c786e, /* 2661 */
128'h7800737469622d73732d6d756e2c786e, /* 2662 */
128'h726566736e6172742d6d756e2c786e6c, /* 2663 */
128'h722d6b63732c786e6c7800737469622d, /* 2664 */
128'h6572662d78616d2d697073006f697461, /* 2665 */
128'h722d656761746c6f760079636e657571, /* 2666 */
128'h70772d656c6261736964007365676e61, /* 2667 */
128'h65726464612d63616d2d6c61636f6c00, /* 2668 */
128'h6700736c6c65632d6f69706723007373, /* 2669 */
128'h780072656c6c6f72746e6f632d6f6970, /* 2670 */
128'h7800737475706e692d6c6c612c786e6c, /* 2671 */
128'h322d737475706e692d6c6c612c786e6c, /* 2672 */
128'h75616665642d74756f642c786e6c7800, /* 2673 */
128'h6665642d74756f642c786e6c7800746c, /* 2674 */
128'h6f6970672c786e6c7800322d746c7561, /* 2675 */
128'h6f6970672c786e6c780068746469772d, /* 2676 */
128'h746e692c786e6c780068746469772d32, /* 2677 */
128'h7800746e65736572702d747075727265, /* 2678 */
128'h786e6c78006c6175642d73692c786e6c, /* 2679 */
128'h6e6c7800746c75616665642d6972742c, /* 2680 */
128'h00322d746c75616665642d6972742c78, /* 2681 */
128'h0000000000203a642520656369766544, /* 2682 */
128'h00203a6425206563697665642073250a, /* 2683 */
128'h00000000203a6425206563697665440a, /* 2684 */
128'h000a656369766564206e776f6e6b6e75, /* 2685 */
128'h00000a2973252c73252870756b6f6f6c, /* 2686 */
128'h7265206c616e7265746e692070636864, /* 2687 */
128'h00000000000000000a7025202c726f72, /* 2688 */
128'h5145525f5043484420676e69646e6553, /* 2689 */
128'h4b434120504348440000000a54534555, /* 2690 */
128'h696c432050434844000000000000000a, /* 2691 */
128'h203a7373657264644120504920746e65, /* 2692 */
128'h0000000a64252e64252e64252e642520, /* 2693 */
128'h73657264644120504920726576726553, /* 2694 */
128'h0a64252e64252e64252e642520203a73, /* 2695 */
128'h6120726574756f520000000000000000, /* 2696 */
128'h252e64252e642520203a737365726464, /* 2697 */
128'h6b73616d2074654e0000000a64252e64, /* 2698 */
128'h64252e642520203a7373657264646120, /* 2699 */
128'h697420657361654c000a64252e64252e, /* 2700 */
128'h00000000000000000a6425203d20656d, /* 2701 */
128'h00000a22732522203d206e69616d6f64, /* 2702 */
128'h00000a22732522203d20726576726573, /* 2703 */
128'h000000000a44455050494b53204b4341, /* 2704 */
128'h000000000000000a4b414e2050434844, /* 2705 */
128'h73657264646120646574736575716552, /* 2706 */
128'h0000000000000a646573756665722073, /* 2707 */
128'h000000000000000a732520726f727245, /* 2708 */
128'h6e6f6974706f2064656c646e61686e75, /* 2709 */
128'h656c646e61686e55000000000a642520, /* 2710 */
128'h64252065646f63706f20504348442064, /* 2711 */
128'h20676e69646e6553000000000000000a, /* 2712 */
128'h000a595245564f435349445f50434844, /* 2713 */
128'h00000000000a29732528726f72726570, /* 2714 */
128'h3a2043414d2073250000000030687465, /* 2715 */
128'h3a583230253a583230253a5832302520, /* 2716 */
128'h000a583230253a583230253a58323025, /* 2717 */
128'h484420646e65732074276e646c756f43, /* 2718 */
128'h206e6f20595245564f43534944205043, /* 2719 */
128'h00000a7325203a732520656369766564, /* 2720 */
128'h5043484420726f6620676e6974696157, /* 2721 */
128'h2020202020202020000a524546464f5f, /* 2722 */
128'h00000000000063250000000000000020, /* 2723 */
128'h0000005832302520000000000000002e, /* 2724 */
128'h00000000732573250000000000000a0a, /* 2725 */
128'h00000000007325203a646c697542202c, /* 2726 */
128'h73257a4820756c250000000000007325, /* 2727 */
128'h0000000000756c250000000000000000, /* 2728 */
128'h0073257a4863252000000000646c252e, /* 2729 */
128'h00000000007325736574794220756c25, /* 2730 */
128'h00003a786c3830250073254269632520, /* 2731 */
128'h000a73252020202000786c6c2a302520, /* 2732 */
128'h000000203a5d64255b6e6f6974636553, /* 2733 */
128'h25203d206465726975716572206e656c, /* 2734 */
128'h000a7825203d206c6175746361202c58, /* 2735 */
128'h302c782578302c7825287970636d656d, /* 2736 */
128'h25287465736d656d00000a3b29782578, /* 2737 */
128'h00000000000a3b29782578302c302c78, /* 2738 */
128'h0000000054455346464f5f4f4c43414d, /* 2739 */
128'h0000000054455346464f5f494843414d, /* 2740 */
128'h000000000054455346464f5f524c5054, /* 2741 */
128'h000000000054455346464f5f53434654, /* 2742 */
128'h0054455346464f5f4c5254434f49444d, /* 2743 */
128'h000000000054455346464f5f53434652, /* 2744 */
128'h00000000000054455346464f5f525352, /* 2745 */
128'h000000000054455346464f5f44414252, /* 2746 */
128'h000000000054455346464f5f524c5052, /* 2747 */
128'h46464f5f524c5052000000003f3f3f3f, /* 2748 */
128'h0000000000000047000064252b544553, /* 2749 */
128'h0a50495049203d206f746f7250205049, /* 2750 */
128'h00000000000000540000000000000000, /* 2751 */
128'h000a504745203d206f746f7250205049, /* 2752 */
128'h000a505550203d206f746f7250205049, /* 2753 */
128'h0000000a3a7265646165682074736574, /* 2754 */
128'h000a3a73746e65746e6f632074736574, /* 2755 */
128'h000a504449203d206f746f7250205049, /* 2756 */
128'h00000a5054203d206f746f7250205049, /* 2757 */
128'h0a50434344203d206f746f7250205049, /* 2758 */
128'h00000000000000360000000000000000, /* 2759 */
128'h0a50565352203d206f746f7250205049, /* 2760 */
128'h6f746f72502050490000000000000000, /* 2761 */
128'h6f746f7250205049000a455247203d20, /* 2762 */
128'h6f746f7250205049000a505345203d20, /* 2763 */
128'h6f746f725020504900000a4841203d20, /* 2764 */
128'h6f746f7250205049000a50544d203d20, /* 2765 */
128'h0000000000000a485054454542203d20, /* 2766 */
128'h5041434e45203d206f746f7250205049, /* 2767 */
128'h000000000000004d000000000000000a, /* 2768 */
128'h0a504d4f43203d206f746f7250205049, /* 2769 */
128'h6f746f72502050490000000000000000, /* 2770 */
128'h00000000000000000a50544353203d20, /* 2771 */
128'h494c504455203d206f746f7250205049, /* 2772 */
128'h6f746f725020504900000000000a4554, /* 2773 */
128'h00000000000000000a534c504d203d20, /* 2774 */
128'h000a574152203d206f746f7250205049, /* 2775 */
128'h7075736e75203d206f746f7270205049, /* 2776 */
128'h000000000a2978252820646574726f70, /* 2777 */
128'h257830203d20657079745f6f746f7270, /* 2778 */
128'h656c646e61686e750000000000000a78, /* 2779 */
128'h0000000a21747075727265746e692064, /* 2780 */
128'h000a726464612043414d207075746553, /* 2781 */
128'h00000a786c253a786c25203d2043414d, /* 2782 */
128'h3025203d20737365726464612043414d, /* 2783 */
128'h3230253a783230253a783230253a7832, /* 2784 */
128'h0000000a2e783230253a783230253a78, /* 2785 */
128'h75727265746e692074656e7265687445, /* 2786 */
128'h0a646c25203d20737574617473207470, /* 2787 */
128'h65687420746f6f420000000000000000, /* 2788 */
128'h2e6d6172676f727020646564616f6c20, /* 2789 */
128'h2c657962646f6f4700000000000a2e2e, /* 2790 */
128'h000000000a2e2e2e207265746f6f6220, /* 2791 */
128'h00007f7c5d5b3f3e3d3c3b3a2c2b2a22, /* 2792 */
128'h007f7c5d5b3f3e3d3c3b3a2e2c2b2a22, /* 2793 */
128'h66656463626139383736353433323130, /* 2794 */
128'h72776f6c2f6372730000000000000000, /* 2795 */
128'h00000000000000632e636d6d5f637369, /* 2796 */
128'h61625f6473203d3d20657361625f6473, /* 2797 */
128'h5f63736972776f6c00726464615f6573, /* 2798 */
128'h000a74756f656d6974207325203a6473, /* 2799 */
128'h616d202c6465766f6d65722064726143, /* 2800 */
128'h6425206f74206465676e616863206b73, /* 2801 */
128'h736e692064726143000000000000000a, /* 2802 */
128'h6e616863206b73616d202c6465747265, /* 2803 */
128'h0000000000000a6425206f7420646567, /* 2804 */
128'h25207461206465746165726320636d6d, /* 2805 */
128'h0000000a7825203d2074736f68202c78, /* 2806 */
128'h0000000000006f4e0000000000736559, /* 2807 */
128'h002020203a434d4d0000000052444420, /* 2808 */
128'h00000000000a7325203a656369766544, /* 2809 */
128'h3a4449207265727574636166756e614d, /* 2810 */
128'h0a7825203a4d454f000000000a782520, /* 2811 */
128'h6325203a656d614e0000000000000000, /* 2812 */
128'h0000000000000a206325632563256325, /* 2813 */
128'h00000a6425203a646565705320737542, /* 2814 */
128'h25203a79746963617061432068676948, /* 2815 */
128'h79746963617061430000000000000a73, /* 2816 */
128'h7464695720737542000000000000203a, /* 2817 */
128'h000000000a73257469622d6425203a68, /* 2818 */
128'h0000007825782520000000203a78250a, /* 2819 */
128'h00000000000064735f63736972776f6c, /* 2820 */
128'h0000000065646f6d206e776f6e6b6e55, /* 2821 */
128'h7830203a726f72724520737574617453, /* 2822 */
128'h2074756f656d69540000000a58383025, /* 2823 */
128'h616572206472616320676e6974696177, /* 2824 */
128'h6c69616620636d6d00000000000a7964, /* 2825 */
128'h6d6320706f747320646e6573206f7420, /* 2826 */
128'h6f6c62203a434d4d0000000000000a64, /* 2827 */
128'h20786c257830207265626d756e206b63, /* 2828 */
128'h6c2578302878616d2073646565637865, /* 2829 */
128'h203d3e20434d4d6500000000000a2978, /* 2830 */
128'h726f6620646572697571657220342e34, /* 2831 */
128'h642072657375206465636e61686e6520, /* 2832 */
128'h000000000000000a6165726120617461, /* 2833 */
128'h757320746f6e2073656f642064726143, /* 2834 */
128'h696e6f697469747261702074726f7070, /* 2835 */
128'h656f64206472614300000000000a676e, /* 2836 */
128'h20434820656e6966656420746f6e2073, /* 2837 */
128'h00000a657a69732070756f7267205057, /* 2838 */
128'h636e61686e6520617461642072657355, /* 2839 */
128'h5720434820746f6e2061657261206465, /* 2840 */
128'h696c6120657a69732070756f72672050, /* 2841 */
128'h72617020692550470000000a64656e67, /* 2842 */
128'h505720434820746f6e206e6f69746974, /* 2843 */
128'h67696c6120657a69732070756f726720, /* 2844 */
128'h656f642064726143000000000a64656e, /* 2845 */
128'h6e652074726f7070757320746f6e2073, /* 2846 */
128'h657475626972747461206465636e6168, /* 2847 */
128'h6e65206c61746f54000000000000000a, /* 2848 */
128'h6563786520657a6973206465636e6168, /* 2849 */
128'h20752528206d756d6978616d20736465, /* 2850 */
128'h656f64206472614300000a297525203e, /* 2851 */
128'h6f682074726f7070757320746f6e2073, /* 2852 */
128'h61702064656c6c6f72746e6f63207473, /* 2853 */
128'h6572206574697277206e6f6974697472, /* 2854 */
128'h6e6974746573207974696c696261696c, /* 2855 */
128'h726c61206472614300000000000a7367, /* 2856 */
128'h64656e6f697469747261702079646165, /* 2857 */
128'h206f6e203a434d4d000000000000000a, /* 2858 */
128'h0000000a746e65736572702064726163, /* 2859 */
128'h73657220746f6e206469642064726143, /* 2860 */
128'h20656761746c6f76206f7420646e6f70, /* 2861 */
128'h00000000000000000a217463656c6573, /* 2862 */
128'h7463656c6573206f7420656c62616e75, /* 2863 */
128'h00000000000000000a65646f6d206120, /* 2864 */
128'h646e756f66206473635f747865206f4e, /* 2865 */
128'h78363025206e614d0000000000000a21, /* 2866 */
128'h000000783430257834302520726e5320, /* 2867 */
128'h00000000632563256325632563256325, /* 2868 */
128'h6167656c20434d4d00000064252e6425, /* 2869 */
128'h636167654c2044530000000000007963, /* 2870 */
128'h6867694820434d4d0000000000000079, /* 2871 */
128'h0000297a484d36322820646565705320, /* 2872 */
128'h35282064656570532068676948204453, /* 2873 */
128'h6867694820434d4d000000297a484d30, /* 2874 */
128'h0000297a484d32352820646565705320, /* 2875 */
128'h7a484d32352820323552444420434d4d, /* 2876 */
128'h31524453205348550000000000000029, /* 2877 */
128'h00000000000000297a484d3532282032, /* 2878 */
128'h7a484d30352820353252445320534855, /* 2879 */
128'h35524453205348550000000000000029, /* 2880 */
128'h000000000000297a484d303031282030, /* 2881 */
128'h7a484d30352820303552444420534855, /* 2882 */
128'h31524453205348550000000000000029, /* 2883 */
128'h0000000000297a484d38303228203430, /* 2884 */
128'h0000297a484d30303228203030325348, /* 2885 */
128'h6f6e2064252065636976654420434d4d, /* 2886 */
128'h00000000000000000a646e756f662074, /* 2887 */
128'h000000000000445300000000434d4d65, /* 2888 */
128'h000000297325282000006425203a7325, /* 2889 */
128'h6e656c20656c69460000000000636d6d, /* 2890 */
128'h000000000000000a6425203d20687467, /* 2891 */
128'h6f6f7420687461702074736575716552, /* 2892 */
128'h00000000000a646c25202e676e6f6c20, /* 2893 */
128'h732522203a717277000000000000002f, /* 2894 */
128'h0a64253d657a69736b636f6c62202c22, /* 2895 */
128'h20657669656365520000000000000000, /* 2896 */
128'h0000000000000a2e646e6520656c6966, /* 2897 */
128'h656c6c6163207172775f656c646e6168, /* 2898 */
128'h206c6167656c6c4900000000000a2e64, /* 2899 */
128'h0a2e6e6f6974617265706f2050544654, /* 2900 */
128'h206f74206c6961460000000000000000, /* 2901 */
128'h2172657669726420445320746e756f6d, /* 2902 */
128'h6f6f622064616f4c000000000000000a, /* 2903 */
128'h726f6d656d206f746e69206e69622e74, /* 2904 */
128'h6e69622e746f6f620000000000000a79, /* 2905 */
128'h742064656c6961460000000000000000, /* 2906 */
128'h0000000a21746f6f62206e65706f206f, /* 2907 */
128'h69662065736f6c63206f74206c696166, /* 2908 */
128'h206f74206c696166000000000021656c, /* 2909 */
128'h00000000216b73696420746e756f6d75, /* 2910 */
128'h20736574796220642520646564616f4c, /* 2911 */
128'h7365726464612079726f6d656d206f74, /* 2912 */
128'h622e746f6f62206d6f72662078252073, /* 2913 */
128'h0a2e736574796220642520666f206e69, /* 2914 */
128'h666c652064616f6c0000000000000000, /* 2915 */
128'h000a79726f6d656d20524444206f7420, /* 2916 */
128'h2064656c696166206461657220666c65, /* 2917 */
128'h0000000064252065646f632068746977, /* 2918 */
128'h20746f6f622d750a000000005c2d2f7c, /* 2919 */
128'h67617473207473726966206465736162, /* 2920 */
128'h00000a726564616f6c20746f6f622065, /* 2921 */
128'h696166207325206e6f69747265737361, /* 2922 */
128'h696c202c732520656c6966202c64656c, /* 2923 */
128'h206e6f6974636e7566202c642520656e, /* 2924 */
128'h3a4552554c49414600000000000a7325, /* 2925 */
128'h74612078257830203d21207825783020, /* 2926 */
128'h00000a2e782578302074657366666f20, /* 2927 */
128'h7025203d203270202c7025203d203170, /* 2928 */
128'h2020202020202020000000000000000a, /* 2929 */
128'h08080808080808080000000000202020, /* 2930 */
128'h20676e69747465730000000000080808, /* 2931 */
128'h20676e69747365740000000000007525, /* 2932 */
128'h3a4552554c4941460000000000007525, /* 2933 */
128'h64612064616220656c626973736f7020, /* 2934 */
128'h666f20746120656e696c207373657264, /* 2935 */
128'h00000000000a2e782578302074657366, /* 2936 */
128'h7478656e206f7420676e697070696b53, /* 2937 */
128'h000000000000000a2e2e2e7473657420, /* 2938 */
128'h20202020200808080808080808080808, /* 2939 */
128'h08080808080808080808202020202020, /* 2940 */
128'h00000000000820080000000000000008, /* 2941 */
128'h78302073692065676e61722074736574, /* 2942 */
128'h00000000000a70257830206f74207025, /* 2943 */
128'h000000000075252f00752520706f6f4c, /* 2944 */
128'h6441206b637574530000000000000a3a, /* 2945 */
128'h0000203a732520200000007373657264, /* 2946 */
128'h00000a2e656e6f4400000000000a6b6f, /* 2947 */
128'h4d415244206c6174656d20657261420a, /* 2948 */
128'h65747365746d656d00000a7473657420, /* 2949 */
128'h20302e332e34206e6f69737265762072, /* 2950 */
128'h000000000000000a297469622d642528, /* 2951 */
128'h30322029432820746867697279706f43, /* 2952 */
128'h2073656c7261684320323130322d3130, /* 2953 */
128'h000000000000000a2e6e6f62617a6143, /* 2954 */
128'h74207265646e75206465736e6563694c, /* 2955 */
128'h50206c6172656e654720554e47206568, /* 2956 */
128'h65762065736e6563694c2063696c6275, /* 2957 */
128'h0a2e29796c6e6f282032206e6f697372, /* 2958 */
128'h5f676e696b726f770000000000000000, /* 2959 */
128'h20646c25202c424b6425203d20746573, /* 2960 */
128'h6c25202c736e6f697463757274736e69, /* 2961 */
128'h203d20495043202c73656c6379632064, /* 2962 */
128'h00000000000000000a646c252e646c25, /* 2963 */
128'h00000a0d21646c726f57206f6c6c6548, /* 2964 */
128'h3d20676e697474657320686374697753, /* 2965 */
128'h00000a0d70617274000000000a582520, /* 2966 */
128'hefcdab8967452301cccccccccccccccd, /* 2967 */
128'h10000000200000001032547698badcfe, /* 2968 */
128'h55555555555555555851f42d4c957f2d, /* 2969 */
128'h0000000000000000aaaaaaaaaaaaaaaa, /* 2970 */
128'h00000000000000000000000000000000, /* 2971 */
128'h00000000000000000000000000000000, /* 2972 */
128'h00000000000000000000000000000000, /* 2973 */
128'h00000000000000000000000000000000, /* 2974 */
128'h00000000000000000000000000000000, /* 2975 */
128'h00004b4d47545045000000030f060301, /* 2976 */
128'h000000003000000000000000004b4d47, /* 2977 */
128'h00000000ffffffff0000000000000000, /* 2978 */
128'h0000646d635f6473000000000c000000, /* 2979 */
128'h00000000ffffffff00006772615f6473, /* 2980 */
128'h000000002f7c5c2d0000000087feb2e8, /* 2981 */
128'hffffffff000000060000000087feb4a0, /* 2982 */
128'h0000000087fe70800000000000000000, /* 2983 */
128'h00000000000000000000000000000042, /* 2984 */
128'h00000000000000000000000000000000, /* 2985 */
128'h00000000000000000000000000000000, /* 2986 */
128'h00000000000000000000000000000000, /* 2987 */
128'h00000000000000000000000000000000, /* 2988 */
128'h00000000000000000000000000000000, /* 2989 */
128'h00000000000000000000000000000000, /* 2990 */
128'h00000000000000000000000000000000, /* 2991 */
128'h00000000000000000000000000000000, /* 2992 */
128'h00000000000000000000000000000000, /* 2993 */
128'h00000000000000000000000000000000, /* 2994 */
128'h00000000000000000000000000000000, /* 2995 */
128'h00000000000000000000000000000000, /* 2996 */
128'h00000000000000000000000000000000, /* 2997 */
128'h00000000000000000000000000000000, /* 2998 */
128'h00000000000000000000000000000000, /* 2999 */
128'h00000000000000000000000000000000, /* 3000 */
128'h00000000000000000000000000000000, /* 3001 */
128'h00000000000000000000000000000000, /* 3002 */
128'h00000000000000000000000000000000, /* 3003 */
128'h00000000000000000000000000000000, /* 3004 */
128'h00000000000000000000000000000000, /* 3005 */
128'h00000000000000000000000000000000, /* 3006 */
128'h00000000000000000000000000000000, /* 3007 */
128'h00000000000000000000000000000000, /* 3008 */
128'h00000000000000000000000000000000, /* 3009 */
128'h00000000000000000000000000000000, /* 3010 */
128'h00000000000000000000000000000000, /* 3011 */
128'h00000000000000000000000000000000, /* 3012 */
128'h00000000000000000000000000000000, /* 3013 */
128'h00000000000000000000000000000000, /* 3014 */
128'h00000000000000000000000000000000, /* 3015 */
128'h00000000000000000000000000000000, /* 3016 */
128'h00000000000000000000000000000000, /* 3017 */
128'h00000000000000000000000000000000, /* 3018 */
128'h00000000000000000000000000000000, /* 3019 */
128'h00000000000000000000000000000000, /* 3020 */
128'h00000000000000000000000000000000, /* 3021 */
128'h00000000000000000000000000000000, /* 3022 */
128'h00000000000000000000000000000000, /* 3023 */
128'h00000000000000000000000000000000, /* 3024 */
128'h00000000000000000000000000000000, /* 3025 */
128'h00000000000000000000000000000000, /* 3026 */
128'h00000000000000000000000000000000, /* 3027 */
128'h00000000000000000000000000000000, /* 3028 */
128'h00000000000000000000000000000000, /* 3029 */
128'h00000000000000000000000000000000, /* 3030 */
128'h00000000000000000000000000000000, /* 3031 */
128'h00000000000000000000000000000000, /* 3032 */
128'h00000000000000000000000000000000, /* 3033 */
128'h00000000000000000000000000000000, /* 3034 */
128'h00000000000000000000000000000000, /* 3035 */
128'h00000000000000000000000000000000, /* 3036 */
128'h00000000000000000000000000000000, /* 3037 */
128'h00000000000000000000000000000000, /* 3038 */
128'h00000000000000000000000000000000, /* 3039 */
128'h00000000000000000000000000000000, /* 3040 */
128'h00000000000000000000000000000000, /* 3041 */
128'h00000000000000000000000000000000, /* 3042 */
128'h00000000000000000000000000000000, /* 3043 */
128'h00000000000000000000000000000000, /* 3044 */
128'h00000000000000000000000000000000, /* 3045 */
128'h00000000000000000000000000000000, /* 3046 */
128'h00000000000000000000000000000000, /* 3047 */
128'h00000000000000000000000000000000, /* 3048 */
128'h00000000000000000000000000000000, /* 3049 */
128'h00000000000000000000000000000000, /* 3050 */
128'h00000000000000000000000000000000, /* 3051 */
128'h00000000000000000000000000000000, /* 3052 */
128'h00000000000000000000000000000000, /* 3053 */
128'h00000000000000000000000000000000, /* 3054 */
128'h00000000000000000000000000000000, /* 3055 */
128'h00000000000000000000000000000000, /* 3056 */
128'h00000000000000000000000000000000, /* 3057 */
128'h00000000000000000000000000000000, /* 3058 */
128'h00000000000000000000000000000000, /* 3059 */
128'h00000000000000000000000000000000, /* 3060 */
128'h00000000000000000000000000000000, /* 3061 */
128'h00000000000000000000000000000000, /* 3062 */
128'h00000000000000000000000000000000, /* 3063 */
128'h00000000000000000000000000000000, /* 3064 */
128'h00000000000000000000000000000000, /* 3065 */
128'h00000000000000000000000000000000, /* 3066 */
128'h00000000000000000000000000000000, /* 3067 */
128'h00000000000000000000000000000000, /* 3068 */
128'h00000000000000000000000000000000, /* 3069 */
128'h00000000000000000000000000000000, /* 3070 */
128'h00000000000000000000000000000000, /* 3071 */
128'h00000000000000000000000000000000, /* 3072 */
128'h00000000000000000000000000000000, /* 3073 */
128'h00000000000000000000000000000000, /* 3074 */
128'h00000000000000000000000000000000, /* 3075 */
128'h00000000000000000000000000000000, /* 3076 */
128'h00000000000000000000000000000000, /* 3077 */
128'h00000000000000000000000000000000, /* 3078 */
128'h00000000000000000000000000000000, /* 3079 */
128'h00000000000000000000000000000000, /* 3080 */
128'h00000000000000000000000000000000, /* 3081 */
128'h00000000000000000000000000000000, /* 3082 */
128'h00000000000000000000000000000000, /* 3083 */
128'h00000000000000000000000000000000, /* 3084 */
128'h00000000000000000000000000000000, /* 3085 */
128'h00000000000000000000000000000000, /* 3086 */
128'h00000000000000000000000000000000, /* 3087 */
128'h00000000000000000000000000000000, /* 3088 */
128'h00000000000000000000000000000000, /* 3089 */
128'h00000000000000000000000000000000, /* 3090 */
128'h00000000000000000000000000000000, /* 3091 */
128'h00000000000000000000000000000000, /* 3092 */
128'h00000000000000000000000000000000, /* 3093 */
128'h00000000000000000000000000000000, /* 3094 */
128'h00000000000000000000000000000000, /* 3095 */
128'h00000000000000000000000000000000, /* 3096 */
128'h00000000000000000000000000000000, /* 3097 */
128'h00000000000000000000000000000000, /* 3098 */
128'h00000000000000000000000000000000, /* 3099 */
128'h00000000000000000000000000000000, /* 3100 */
128'h00000000000000000000000000000000, /* 3101 */
128'h00000000000000000000000000000000, /* 3102 */
128'h00000000000000000000000000000000, /* 3103 */
128'h00000000000000000000000000000000, /* 3104 */
128'h00000000000000000000000000000000, /* 3105 */
128'h00000000000000000000000000000000, /* 3106 */
128'h00000000000000000000000000000000, /* 3107 */
128'h00000000000000000000000000000000, /* 3108 */
128'h00000000000000000000000000000000, /* 3109 */
128'h00000000000000000000000000000000, /* 3110 */
128'h00000000000000000000000000000000, /* 3111 */
128'h00000000000000000000000000000000, /* 3112 */
128'h00000000000000000000000000000000, /* 3113 */
128'h00000000000000000000000000000000, /* 3114 */
128'h00000000000000000000000000000000, /* 3115 */
128'h00000000000000000000000000000000, /* 3116 */
128'h00000000000000000000000000000000, /* 3117 */
128'h00000000000000000000000000000000, /* 3118 */
128'h00000000000000000000000000000000, /* 3119 */
128'h00000000000000000000000000000000, /* 3120 */
128'h00000000000000000000000000000000, /* 3121 */
128'h00000000000000000000000000000000, /* 3122 */
128'h00000000000000000000000000000000, /* 3123 */
128'h00000000000000000000000000000000, /* 3124 */
128'h00000000000000000000000000000000, /* 3125 */
128'h00000000000000000000000000000000, /* 3126 */
128'h00000000000000000000000000000000, /* 3127 */
128'h00000000000000000000000000000000, /* 3128 */
128'h00000000000000000000000000000000, /* 3129 */
128'h00000000000000000000000000000000, /* 3130 */
128'h00000000000000000000000000000000, /* 3131 */
128'h00000000000000000000000000000000, /* 3132 */
128'h00000000000000000000000000000000, /* 3133 */
128'h00000000000000000000000000000000, /* 3134 */
128'h00000000000000000000000000000000, /* 3135 */
128'h00000000000000000000000000000000, /* 3136 */
128'h00000000000000000000000000000000, /* 3137 */
128'h00000000000000000000000000000000, /* 3138 */
128'h00000000000000000000000000000000, /* 3139 */
128'h00000000000000000000000000000000, /* 3140 */
128'h00000000000000000000000000000000, /* 3141 */
128'h00000000000000000000000000000000, /* 3142 */
128'h00000000000000000000000000000000, /* 3143 */
128'h00000000000000000000000000000000, /* 3144 */
128'h00000000000000000000000000000000, /* 3145 */
128'h00000000000000000000000000000000, /* 3146 */
128'h00000000000000000000000000000000, /* 3147 */
128'h00000000000000000000000000000000, /* 3148 */
128'h00000000000000000000000000000000, /* 3149 */
128'h00000000000000000000000000000000, /* 3150 */
128'h00000000000000000000000000000000, /* 3151 */
128'h00000000000000000000000000000000, /* 3152 */
128'h00000000000000000000000000000000, /* 3153 */
128'h00000000000000000000000000000000, /* 3154 */
128'h00000000000000000000000000000000, /* 3155 */
128'h00000000000000000000000000000000, /* 3156 */
128'h00000000000000000000000000000000, /* 3157 */
128'h00000000000000000000000000000000, /* 3158 */
128'h00000000000000000000000000000000, /* 3159 */
128'h00000000000000000000000000000000, /* 3160 */
128'h00000000000000000000000000000000, /* 3161 */
128'h00000000000000000000000000000000, /* 3162 */
128'h00000000000000000000000000000000, /* 3163 */
128'h00000000000000000000000000000000, /* 3164 */
128'h00000000000000000000000000000000, /* 3165 */
128'h00000000000000000000000000000000, /* 3166 */
128'h00000000000000000000000000000000, /* 3167 */
128'h00000000000000000000000000000000, /* 3168 */
128'h00000000000000000000000000000000, /* 3169 */
128'h00000000000000000000000000000000, /* 3170 */
128'h00000000000000000000000000000000, /* 3171 */
128'h00000000000000000000000000000000, /* 3172 */
128'h00000000000000000000000000000000, /* 3173 */
128'h00000000000000000000000000000000, /* 3174 */
128'h00000000000000000000000000000000, /* 3175 */
128'h00000000000000000000000000000000, /* 3176 */
128'h00000000000000000000000000000000, /* 3177 */
128'h00000000000000000000000000000000, /* 3178 */
128'h00000000000000000000000000000000, /* 3179 */
128'h00000000000000000000000000000000, /* 3180 */
128'h00000000000000000000000000000000, /* 3181 */
128'h00000000000000000000000000000000, /* 3182 */
128'h00000000000000000000000000000000, /* 3183 */
128'h00000000000000000000000000000000, /* 3184 */
128'h00000000000000000000000000000000, /* 3185 */
128'h00000000000000000000000000000000, /* 3186 */
128'h00000000000000000000000000000000, /* 3187 */
128'h00000000000000000000000000000000, /* 3188 */
128'h00000000000000000000000000000000, /* 3189 */
128'h00000000000000000000000000000000, /* 3190 */
128'h00000000000000000000000000000000, /* 3191 */
128'h00000000000000000000000000000000, /* 3192 */
128'h00000000000000000000000000000000, /* 3193 */
128'h00000000000000000000000000000000, /* 3194 */
128'h00000000000000000000000000000000, /* 3195 */
128'h00000000000000000000000000000000, /* 3196 */
128'h00000000000000000000000000000000, /* 3197 */
128'h00000000000000000000000000000000, /* 3198 */
128'h00000000000000000000000000000000, /* 3199 */
128'h00000000000000000000000000000000, /* 3200 */
128'h00000000000000000000000000000000, /* 3201 */
128'h00000000000000000000000000000000, /* 3202 */
128'h00000000000000000000000000000000, /* 3203 */
128'h00000000000000000000000000000000, /* 3204 */
128'h00000000000000000000000000000000, /* 3205 */
128'h00000000000000000000000000000000, /* 3206 */
128'h00000000000000000000000000000000, /* 3207 */
128'h00000000000000000000000000000000, /* 3208 */
128'h00000000000000000000000000000000, /* 3209 */
128'h00000000000000000000000000000000, /* 3210 */
128'h00000000000000000000000000000000, /* 3211 */
128'h00000000000000000000000000000000, /* 3212 */
128'h00000000000000000000000000000000, /* 3213 */
128'h00000000000000000000000000000000, /* 3214 */
128'h00000000000000000000000000000000, /* 3215 */
128'h00000000000000000000000000000000, /* 3216 */
128'h00000000000000000000000000000000, /* 3217 */
128'h00000000000000000000000000000000, /* 3218 */
128'h00000000000000000000000000000000, /* 3219 */
128'h00000000000000000000000000000000, /* 3220 */
128'h00000000000000000000000000000000, /* 3221 */
128'h00000000000000000000000000000000, /* 3222 */
128'h00000000000000000000000000000000, /* 3223 */
128'h00000000000000000000000000000000, /* 3224 */
128'h00000000000000000000000000000000, /* 3225 */
128'h00000000000000000000000000000000, /* 3226 */
128'h00000000000000000000000000000000, /* 3227 */
128'h00000000000000000000000000000000, /* 3228 */
128'h00000000000000000000000000000000, /* 3229 */
128'h00000000000000000000000000000000, /* 3230 */
128'h00000000000000000000000000000000, /* 3231 */
128'h00000000000000000000000000000000, /* 3232 */
128'h00000000000000000000000000000000, /* 3233 */
128'h00000000000000000000000000000000, /* 3234 */
128'h00000000000000000000000000000000, /* 3235 */
128'h00000000000000000000000000000000, /* 3236 */
128'h00000000000000000000000000000000, /* 3237 */
128'h00000000000000000000000000000000, /* 3238 */
128'h00000000000000000000000000000000, /* 3239 */
128'h00000000000000000000000000000000, /* 3240 */
128'h00000000000000000000000000000000, /* 3241 */
128'h00000000000000000000000000000000, /* 3242 */
128'h00000000000000000000000000000000, /* 3243 */
128'h00000000000000000000000000000000, /* 3244 */
128'h00000000000000000000000000000000, /* 3245 */
128'h00000000000000000000000000000000, /* 3246 */
128'h00000000000000000000000000000000, /* 3247 */
128'h00000000000000000000000000000000, /* 3248 */
128'h00000000000000000000000000000000, /* 3249 */
128'h00000000000000000000000000000000, /* 3250 */
128'h00000000000000000000000000000000, /* 3251 */
128'h00000000000000000000000000000000, /* 3252 */
128'h00000000000000000000000000000000, /* 3253 */
128'h00000000000000000000000000000000, /* 3254 */
128'h00000000000000000000000000000000, /* 3255 */
128'h00000000000000000000000000000000, /* 3256 */
128'h00000000000000000000000000000000, /* 3257 */
128'h00000000000000000000000000000000, /* 3258 */
128'h00000000000000000000000000000000, /* 3259 */
128'h00000000000000000000000000000000, /* 3260 */
128'h00000000000000000000000000000000, /* 3261 */
128'h00000000000000000000000000000000, /* 3262 */
128'h00000000000000000000000000000000, /* 3263 */
128'h00000000000000000000000000000000, /* 3264 */
128'h00000000000000000000000000000000, /* 3265 */
128'h00000000000000000000000000000000, /* 3266 */
128'h00000000000000000000000000000000, /* 3267 */
128'h00000000000000000000000000000000, /* 3268 */
128'h00000000000000000000000000000000, /* 3269 */
128'h00000000000000000000000000000000, /* 3270 */
128'h00000000000000000000000000000000, /* 3271 */
128'h00000000000000000000000000000000, /* 3272 */
128'h00000000000000000000000000000000, /* 3273 */
128'h00000000000000000000000000000000, /* 3274 */
128'h00000000000000000000000000000000, /* 3275 */
128'h00000000000000000000000000000000, /* 3276 */
128'h00000000000000000000000000000000, /* 3277 */
128'h00000000000000000000000000000000, /* 3278 */
128'h00000000000000000000000000000000, /* 3279 */
128'h00000000000000000000000000000000, /* 3280 */
128'h00000000000000000000000000000000, /* 3281 */
128'h00000000000000000000000000000000, /* 3282 */
128'h00000000000000000000000000000000, /* 3283 */
128'h00000000000000000000000000000000, /* 3284 */
128'h00000000000000000000000000000000, /* 3285 */
128'h00000000000000000000000000000000, /* 3286 */
128'h00000000000000000000000000000000, /* 3287 */
128'h00000000000000000000000000000000, /* 3288 */
128'h00000000000000000000000000000000, /* 3289 */
128'h00000000000000000000000000000000, /* 3290 */
128'h00000000000000000000000000000000, /* 3291 */
128'h00000000000000000000000000000000, /* 3292 */
128'h00000000000000000000000000000000, /* 3293 */
128'h00000000000000000000000000000000, /* 3294 */
128'h00000000000000000000000000000000, /* 3295 */
128'h00000000000000000000000000000000, /* 3296 */
128'h00000000000000000000000000000000, /* 3297 */
128'h00000000000000000000000000000000, /* 3298 */
128'h00000000000000000000000000000000, /* 3299 */
128'h00000000000000000000000000000000, /* 3300 */
128'h00000000000000000000000000000000, /* 3301 */
128'h00000000000000000000000000000000, /* 3302 */
128'h00000000000000000000000000000000, /* 3303 */
128'h00000000000000000000000000000000, /* 3304 */
128'h00000000000000000000000000000000, /* 3305 */
128'h00000000000000000000000000000000, /* 3306 */
128'h00000000000000000000000000000000, /* 3307 */
128'h00000000000000000000000000000000, /* 3308 */
128'h00000000000000000000000000000000, /* 3309 */
128'h00000000000000000000000000000000, /* 3310 */
128'h00000000000000000000000000000000, /* 3311 */
128'h00000000000000000000000000000000, /* 3312 */
128'h00000000000000000000000000000000, /* 3313 */
128'h00000000000000000000000000000000, /* 3314 */
128'h00000000000000000000000000000000, /* 3315 */
128'h00000000000000000000000000000000, /* 3316 */
128'h00000000000000000000000000000000, /* 3317 */
128'h00000000000000000000000000000000, /* 3318 */
128'h00000000000000000000000000000000, /* 3319 */
128'h00000000000000000000000000000000, /* 3320 */
128'h00000000000000000000000000000000, /* 3321 */
128'h00000000000000000000000000000000, /* 3322 */
128'h00000000000000000000000000000000, /* 3323 */
128'h00000000000000000000000000000000, /* 3324 */
128'h00000000000000000000000000000000, /* 3325 */
128'h00000000000000000000000000000000, /* 3326 */
128'h00000000000000000000000000000000, /* 3327 */
128'h00000000000000000000000000000000, /* 3328 */
128'h00000000000000000000000000000000, /* 3329 */
128'h00000000000000000000000000000000, /* 3330 */
128'h00000000000000000000000000000000, /* 3331 */
128'h00000000000000000000000000000000, /* 3332 */
128'h00000000000000000000000000000000, /* 3333 */
128'h00000000000000000000000000000000, /* 3334 */
128'h00000000000000000000000000000000, /* 3335 */
128'h00000000000000000000000000000000, /* 3336 */
128'h00000000000000000000000000000000, /* 3337 */
128'h00000000000000000000000000000000, /* 3338 */
128'h00000000000000000000000000000000, /* 3339 */
128'h00000000000000000000000000000000, /* 3340 */
128'h00000000000000000000000000000000, /* 3341 */
128'h00000000000000000000000000000000, /* 3342 */
128'h00000000000000000000000000000000, /* 3343 */
128'h00000000000000000000000000000000, /* 3344 */
128'h00000000000000000000000000000000, /* 3345 */
128'h00000000000000000000000000000000, /* 3346 */
128'h00000000000000000000000000000000, /* 3347 */
128'h00000000000000000000000000000000, /* 3348 */
128'h00000000000000000000000000000000, /* 3349 */
128'h00000000000000000000000000000000, /* 3350 */
128'h00000000000000000000000000000000, /* 3351 */
128'h00000000000000000000000000000000, /* 3352 */
128'h00000000000000000000000000000000, /* 3353 */
128'h00000000000000000000000000000000, /* 3354 */
128'h00000000000000000000000000000000, /* 3355 */
128'h00000000000000000000000000000000, /* 3356 */
128'h00000000000000000000000000000000, /* 3357 */
128'h00000000000000000000000000000000, /* 3358 */
128'h00000000000000000000000000000000, /* 3359 */
128'h00000000000000000000000000000000, /* 3360 */
128'h00000000000000000000000000000000, /* 3361 */
128'h00000000000000000000000000000000, /* 3362 */
128'h00000000000000000000000000000000, /* 3363 */
128'h00000000000000000000000000000000, /* 3364 */
128'h00000000000000000000000000000000, /* 3365 */
128'h00000000000000000000000000000000, /* 3366 */
128'h00000000000000000000000000000000, /* 3367 */
128'h00000000000000000000000000000000, /* 3368 */
128'h00000000000000000000000000000000, /* 3369 */
128'h00000000000000000000000000000000, /* 3370 */
128'h00000000000000000000000000000000, /* 3371 */
128'h00000000000000000000000000000000, /* 3372 */
128'h00000000000000000000000000000000, /* 3373 */
128'h00000000000000000000000000000000, /* 3374 */
128'h00000000000000000000000000000000, /* 3375 */
128'h00000000000000000000000000000000, /* 3376 */
128'h00000000000000000000000000000000, /* 3377 */
128'h00000000000000000000000000000000, /* 3378 */
128'h00000000000000000000000000000000, /* 3379 */
128'h00000000000000000000000000000000, /* 3380 */
128'h00000000000000000000000000000000, /* 3381 */
128'h00000000000000000000000000000000, /* 3382 */
128'h00000000000000000000000000000000, /* 3383 */
128'h00000000000000000000000000000000, /* 3384 */
128'h00000000000000000000000000000000, /* 3385 */
128'h00000000000000000000000000000000, /* 3386 */
128'h00000000000000000000000000000000, /* 3387 */
128'h00000000000000000000000000000000, /* 3388 */
128'h00000000000000000000000000000000, /* 3389 */
128'h00000000000000000000000000000000, /* 3390 */
128'h00000000000000000000000000000000, /* 3391 */
128'h00000000000000000000000000000000, /* 3392 */
128'h00000000000000000000000000000000, /* 3393 */
128'h00000000000000000000000000000000, /* 3394 */
128'h00000000000000000000000000000000, /* 3395 */
128'h00000000000000000000000000000000, /* 3396 */
128'h00000000000000000000000000000000, /* 3397 */
128'h00000000000000000000000000000000, /* 3398 */
128'h00000000000000000000000000000000, /* 3399 */
128'h00000000000000000000000000000000, /* 3400 */
128'h00000000000000000000000000000000, /* 3401 */
128'h00000000000000000000000000000000, /* 3402 */
128'h00000000000000000000000000000000, /* 3403 */
128'h00000000000000000000000000000000, /* 3404 */
128'h00000000000000000000000000000000, /* 3405 */
128'h00000000000000000000000000000000, /* 3406 */
128'h00000000000000000000000000000000, /* 3407 */
128'h00000000000000000000000000000000, /* 3408 */
128'h00000000000000000000000000000000, /* 3409 */
128'h00000000000000000000000000000000, /* 3410 */
128'h00000000000000000000000000000000, /* 3411 */
128'h00000000000000000000000000000000, /* 3412 */
128'h00000000000000000000000000000000, /* 3413 */
128'h00000000000000000000000000000000, /* 3414 */
128'h00000000000000000000000000000000, /* 3415 */
128'h00000000000000000000000000000000, /* 3416 */
128'h00000000000000000000000000000000, /* 3417 */
128'h00000000000000000000000000000000, /* 3418 */
128'h00000000000000000000000000000000, /* 3419 */
128'h00000000000000000000000000000000, /* 3420 */
128'h00000000000000000000000000000000, /* 3421 */
128'h00000000000000000000000000000000, /* 3422 */
128'h00000000000000000000000000000000, /* 3423 */
128'h00000000000000000000000000000000, /* 3424 */
128'h00000000000000000000000000000000, /* 3425 */
128'h00000000000000000000000000000000, /* 3426 */
128'h00000000000000000000000000000000, /* 3427 */
128'h00000000000000000000000000000000, /* 3428 */
128'h00000000000000000000000000000000, /* 3429 */
128'h00000000000000000000000000000000, /* 3430 */
128'h00000000000000000000000000000000, /* 3431 */
128'h00000000000000000000000000000000, /* 3432 */
128'h00000000000000000000000000000000, /* 3433 */
128'h00000000000000000000000000000000, /* 3434 */
128'h00000000000000000000000000000000, /* 3435 */
128'h00000000000000000000000000000000, /* 3436 */
128'h00000000000000000000000000000000, /* 3437 */
128'h00000000000000000000000000000000, /* 3438 */
128'h00000000000000000000000000000000, /* 3439 */
128'h00000000000000000000000000000000, /* 3440 */
128'h00000000000000000000000000000000, /* 3441 */
128'h00000000000000000000000000000000, /* 3442 */
128'h00000000000000000000000000000000, /* 3443 */
128'h00000000000000000000000000000000, /* 3444 */
128'h00000000000000000000000000000000, /* 3445 */
128'h00000000000000000000000000000000, /* 3446 */
128'h00000000000000000000000000000000, /* 3447 */
128'h00000000000000000000000000000000, /* 3448 */
128'h00000000000000000000000000000000, /* 3449 */
128'h00000000000000000000000000000000, /* 3450 */
128'h00000000000000000000000000000000, /* 3451 */
128'h00000000000000000000000000000000, /* 3452 */
128'h00000000000000000000000000000000, /* 3453 */
128'h00000000000000000000000000000000, /* 3454 */
128'h00000000000000000000000000000000, /* 3455 */
128'h00000000000000000000000000000000, /* 3456 */
128'h00000000000000000000000000000000, /* 3457 */
128'h00000000000000000000000000000000, /* 3458 */
128'h00000000000000000000000000000000, /* 3459 */
128'h00000000000000000000000000000000, /* 3460 */
128'h00000000000000000000000000000000, /* 3461 */
128'h00000000000000000000000000000000, /* 3462 */
128'h00000000000000000000000000000000, /* 3463 */
128'h00000000000000000000000000000000, /* 3464 */
128'h00000000000000000000000000000000, /* 3465 */
128'h00000000000000000000000000000000, /* 3466 */
128'h00000000000000000000000000000000, /* 3467 */
128'h00000000000000000000000000000000, /* 3468 */
128'h00000000000000000000000000000000, /* 3469 */
128'h00000000000000000000000000000000, /* 3470 */
128'h00000000000000000000000000000000, /* 3471 */
128'h00000000000000000000000000000000, /* 3472 */
128'h00000000000000000000000000000000, /* 3473 */
128'h00000000000000000000000000000000, /* 3474 */
128'h00000000000000000000000000000000, /* 3475 */
128'h00000000000000000000000000000000, /* 3476 */
128'h00000000000000000000000000000000, /* 3477 */
128'h00000000000000000000000000000000, /* 3478 */
128'h00000000000000000000000000000000, /* 3479 */
128'h00000000000000000000000000000000, /* 3480 */
128'h00000000000000000000000000000000, /* 3481 */
128'h00000000000000000000000000000000, /* 3482 */
128'h00000000000000000000000000000000, /* 3483 */
128'h00000000000000000000000000000000, /* 3484 */
128'h00000000000000000000000000000000, /* 3485 */
128'h00000000000000000000000000000000, /* 3486 */
128'h00000000000000000000000000000000, /* 3487 */
128'h00000000000000000000000000000000, /* 3488 */
128'h00000000000000000000000000000000, /* 3489 */
128'h00000000000000000000000000000000, /* 3490 */
128'h00000000000000000000000000000000, /* 3491 */
128'h00000000000000000000000000000000, /* 3492 */
128'h00000000000000000000000000000000, /* 3493 */
128'h00000000000000000000000000000000, /* 3494 */
128'h00000000000000000000000000000000, /* 3495 */
128'h00000000000000000000000000000000, /* 3496 */
128'h00000000000000000000000000000000, /* 3497 */
128'h00000000000000000000000000000000, /* 3498 */
128'h00000000000000000000000000000000, /* 3499 */
128'h00000000000000000000000000000000, /* 3500 */
128'h00000000000000000000000000000000, /* 3501 */
128'h00000000000000000000000000000000, /* 3502 */
128'h00000000000000000000000000000000, /* 3503 */
128'h00000000000000000000000000000000, /* 3504 */
128'h00000000000000000000000000000000, /* 3505 */
128'h00000000000000000000000000000000, /* 3506 */
128'h00000000000000000000000000000000, /* 3507 */
128'h00000000000000000000000000000000, /* 3508 */
128'h00000000000000000000000000000000, /* 3509 */
128'h00000000000000000000000000000000, /* 3510 */
128'h00000000000000000000000000000000, /* 3511 */
128'h00000000000000000000000000000000, /* 3512 */
128'h00000000000000000000000000000000, /* 3513 */
128'h00000000000000000000000000000000, /* 3514 */
128'h00000000000000000000000000000000, /* 3515 */
128'h00000000000000000000000000000000, /* 3516 */
128'h00000000000000000000000000000000, /* 3517 */
128'h00000000000000000000000000000000, /* 3518 */
128'h00000000000000000000000000000000, /* 3519 */
128'h00000000000000000000000000000000, /* 3520 */
128'h00000000000000000000000000000000, /* 3521 */
128'h00000000000000000000000000000000, /* 3522 */
128'h00000000000000000000000000000000, /* 3523 */
128'h00000000000000000000000000000000, /* 3524 */
128'h00000000000000000000000000000000, /* 3525 */
128'h00000000000000000000000000000000, /* 3526 */
128'h00000000000000000000000000000000, /* 3527 */
128'h00000000000000000000000000000000, /* 3528 */
128'h00000000000000000000000000000000, /* 3529 */
128'h00000000000000000000000000000000, /* 3530 */
128'h00000000000000000000000000000000, /* 3531 */
128'h00000000000000000000000000000000, /* 3532 */
128'h00000000000000000000000000000000, /* 3533 */
128'h00000000000000000000000000000000, /* 3534 */
128'h00000000000000000000000000000000, /* 3535 */
128'h00000000000000000000000000000000, /* 3536 */
128'h00000000000000000000000000000000, /* 3537 */
128'h00000000000000000000000000000000, /* 3538 */
128'h00000000000000000000000000000000, /* 3539 */
128'h00000000000000000000000000000000, /* 3540 */
128'h00000000000000000000000000000000, /* 3541 */
128'h00000000000000000000000000000000, /* 3542 */
128'h00000000000000000000000000000000, /* 3543 */
128'h00000000000000000000000000000000, /* 3544 */
128'h00000000000000000000000000000000, /* 3545 */
128'h00000000000000000000000000000000, /* 3546 */
128'h00000000000000000000000000000000, /* 3547 */
128'h00000000000000000000000000000000, /* 3548 */
128'h00000000000000000000000000000000, /* 3549 */
128'h00000000000000000000000000000000, /* 3550 */
128'h00000000000000000000000000000000, /* 3551 */
128'h00000000000000000000000000000000, /* 3552 */
128'h00000000000000000000000000000000, /* 3553 */
128'h00000000000000000000000000000000, /* 3554 */
128'h00000000000000000000000000000000, /* 3555 */
128'h00000000000000000000000000000000, /* 3556 */
128'h00000000000000000000000000000000, /* 3557 */
128'h00000000000000000000000000000000, /* 3558 */
128'h00000000000000000000000000000000, /* 3559 */
128'h00000000000000000000000000000000, /* 3560 */
128'h00000000000000000000000000000000, /* 3561 */
128'h00000000000000000000000000000000, /* 3562 */
128'h00000000000000000000000000000000, /* 3563 */
128'h00000000000000000000000000000000, /* 3564 */
128'h00000000000000000000000000000000, /* 3565 */
128'h00000000000000000000000000000000, /* 3566 */
128'h00000000000000000000000000000000, /* 3567 */
128'h00000000000000000000000000000000, /* 3568 */
128'h00000000000000000000000000000000, /* 3569 */
128'h00000000000000000000000000000000, /* 3570 */
128'h00000000000000000000000000000000, /* 3571 */
128'h00000000000000000000000000000000, /* 3572 */
128'h00000000000000000000000000000000, /* 3573 */
128'h00000000000000000000000000000000, /* 3574 */
128'h00000000000000000000000000000000, /* 3575 */
128'h00000000000000000000000000000000, /* 3576 */
128'h00000000000000000000000000000000, /* 3577 */
128'h00000000000000000000000000000000, /* 3578 */
128'h00000000000000000000000000000000, /* 3579 */
128'h00000000000000000000000000000000, /* 3580 */
128'h00000000000000000000000000000000, /* 3581 */
128'h00000000000000000000000000000000, /* 3582 */
128'h00000000000000000000000000000000, /* 3583 */
128'h00000000000000000000000000000000, /* 3584 */
128'h00000000000000000000000000000000, /* 3585 */
128'h00000000000000000000000000000000, /* 3586 */
128'h00000000000000000000000000000000, /* 3587 */
128'h00000000000000000000000000000000, /* 3588 */
128'h00000000000000000000000000000000, /* 3589 */
128'h00000000000000000000000000000000, /* 3590 */
128'h00000000000000000000000000000000, /* 3591 */
128'h00000000000000000000000000000000, /* 3592 */
128'h00000000000000000000000000000000, /* 3593 */
128'h00000000000000000000000000000000, /* 3594 */
128'h00000000000000000000000000000000, /* 3595 */
128'h00000000000000000000000000000000, /* 3596 */
128'h00000000000000000000000000000000, /* 3597 */
128'h00000000000000000000000000000000, /* 3598 */
128'h00000000000000000000000000000000, /* 3599 */
128'h00000000000000000000000000000000, /* 3600 */
128'h00000000000000000000000000000000, /* 3601 */
128'h00000000000000000000000000000000, /* 3602 */
128'h00000000000000000000000000000000, /* 3603 */
128'h00000000000000000000000000000000, /* 3604 */
128'h00000000000000000000000000000000, /* 3605 */
128'h00000000000000000000000000000000, /* 3606 */
128'h00000000000000000000000000000000, /* 3607 */
128'h00000000000000000000000000000000, /* 3608 */
128'h00000000000000000000000000000000, /* 3609 */
128'h00000000000000000000000000000000, /* 3610 */
128'h00000000000000000000000000000000, /* 3611 */
128'h00000000000000000000000000000000, /* 3612 */
128'h00000000000000000000000000000000, /* 3613 */
128'h00000000000000000000000000000000, /* 3614 */
128'h00000000000000000000000000000000, /* 3615 */
128'h00000000000000000000000000000000, /* 3616 */
128'h00000000000000000000000000000000, /* 3617 */
128'h00000000000000000000000000000000, /* 3618 */
128'h00000000000000000000000000000000, /* 3619 */
128'h00000000000000000000000000000000, /* 3620 */
128'h00000000000000000000000000000000, /* 3621 */
128'h00000000000000000000000000000000, /* 3622 */
128'h00000000000000000000000000000000, /* 3623 */
128'h00000000000000000000000000000000, /* 3624 */
128'h00000000000000000000000000000000, /* 3625 */
128'h00000000000000000000000000000000, /* 3626 */
128'h00000000000000000000000000000000, /* 3627 */
128'h00000000000000000000000000000000, /* 3628 */
128'h00000000000000000000000000000000, /* 3629 */
128'h00000000000000000000000000000000, /* 3630 */
128'h00000000000000000000000000000000, /* 3631 */
128'h00000000000000000000000000000000, /* 3632 */
128'h00000000000000000000000000000000, /* 3633 */
128'h00000000000000000000000000000000, /* 3634 */
128'h00000000000000000000000000000000, /* 3635 */
128'h00000000000000000000000000000000, /* 3636 */
128'h00000000000000000000000000000000, /* 3637 */
128'h00000000000000000000000000000000, /* 3638 */
128'h00000000000000000000000000000000, /* 3639 */
128'h00000000000000000000000000000000, /* 3640 */
128'h00000000000000000000000000000000, /* 3641 */
128'h00000000000000000000000000000000, /* 3642 */
128'h00000000000000000000000000000000, /* 3643 */
128'h00000000000000000000000000000000, /* 3644 */
128'h00000000000000000000000000000000, /* 3645 */
128'h00000000000000000000000000000000, /* 3646 */
128'h00000000000000000000000000000000, /* 3647 */
128'h00000000000000000000000000000000, /* 3648 */
128'h00000000000000000000000000000000, /* 3649 */
128'h00000000000000000000000000000000, /* 3650 */
128'h00000000000000000000000000000000, /* 3651 */
128'h00000000000000000000000000000000, /* 3652 */
128'h00000000000000000000000000000000, /* 3653 */
128'h00000000000000000000000000000000, /* 3654 */
128'h00000000000000000000000000000000, /* 3655 */
128'h00000000000000000000000000000000, /* 3656 */
128'h00000000000000000000000000000000, /* 3657 */
128'h00000000000000000000000000000000, /* 3658 */
128'h00000000000000000000000000000000, /* 3659 */
128'h00000000000000000000000000000000, /* 3660 */
128'h00000000000000000000000000000000, /* 3661 */
128'h00000000000000000000000000000000, /* 3662 */
128'h00000000000000000000000000000000, /* 3663 */
128'h00000000000000000000000000000000, /* 3664 */
128'h00000000000000000000000000000000, /* 3665 */
128'h00000000000000000000000000000000, /* 3666 */
128'h00000000000000000000000000000000, /* 3667 */
128'h00000000000000000000000000000000, /* 3668 */
128'h00000000000000000000000000000000, /* 3669 */
128'h00000000000000000000000000000000, /* 3670 */
128'h00000000000000000000000000000000, /* 3671 */
128'h00000000000000000000000000000000, /* 3672 */
128'h00000000000000000000000000000000, /* 3673 */
128'h00000000000000000000000000000000, /* 3674 */
128'h00000000000000000000000000000000, /* 3675 */
128'h00000000000000000000000000000000, /* 3676 */
128'h00000000000000000000000000000000, /* 3677 */
128'h00000000000000000000000000000000, /* 3678 */
128'h00000000000000000000000000000000, /* 3679 */
128'h00000000000000000000000000000000, /* 3680 */
128'h00000000000000000000000000000000, /* 3681 */
128'h00000000000000000000000000000000, /* 3682 */
128'h00000000000000000000000000000000, /* 3683 */
128'h00000000000000000000000000000000, /* 3684 */
128'h00000000000000000000000000000000, /* 3685 */
128'h00000000000000000000000000000000, /* 3686 */
128'h00000000000000000000000000000000, /* 3687 */
128'h00000000000000000000000000000000, /* 3688 */
128'h00000000000000000000000000000000, /* 3689 */
128'h00000000000000000000000000000000, /* 3690 */
128'h00000000000000000000000000000000, /* 3691 */
128'h00000000000000000000000000000000, /* 3692 */
128'h00000000000000000000000000000000, /* 3693 */
128'h00000000000000000000000000000000, /* 3694 */
128'h00000000000000000000000000000000, /* 3695 */
128'h00000000000000000000000000000000, /* 3696 */
128'h00000000000000000000000000000000, /* 3697 */
128'h00000000000000000000000000000000, /* 3698 */
128'h00000000000000000000000000000000, /* 3699 */
128'h00000000000000000000000000000000, /* 3700 */
128'h00000000000000000000000000000000, /* 3701 */
128'h00000000000000000000000000000000, /* 3702 */
128'h00000000000000000000000000000000, /* 3703 */
128'h00000000000000000000000000000000, /* 3704 */
128'h00000000000000000000000000000000, /* 3705 */
128'h00000000000000000000000000000000, /* 3706 */
128'h00000000000000000000000000000000, /* 3707 */
128'h00000000000000000000000000000000, /* 3708 */
128'h00000000000000000000000000000000, /* 3709 */
128'h00000000000000000000000000000000, /* 3710 */
128'h00000000000000000000000000000000, /* 3711 */
128'h00000000000000000000000000000000, /* 3712 */
128'h00000000000000000000000000000000, /* 3713 */
128'h00000000000000000000000000000000, /* 3714 */
128'h00000000000000000000000000000000, /* 3715 */
128'h00000000000000000000000000000000, /* 3716 */
128'h00000000000000000000000000000000, /* 3717 */
128'h00000000000000000000000000000000, /* 3718 */
128'h00000000000000000000000000000000, /* 3719 */
128'h00000000000000000000000000000000, /* 3720 */
128'h00000000000000000000000000000000, /* 3721 */
128'h00000000000000000000000000000000, /* 3722 */
128'h00000000000000000000000000000000, /* 3723 */
128'h00000000000000000000000000000000, /* 3724 */
128'h00000000000000000000000000000000, /* 3725 */
128'h00000000000000000000000000000000, /* 3726 */
128'h00000000000000000000000000000000, /* 3727 */
128'h00000000000000000000000000000000, /* 3728 */
128'h00000000000000000000000000000000, /* 3729 */
128'h00000000000000000000000000000000, /* 3730 */
128'h00000000000000000000000000000000, /* 3731 */
128'h00000000000000000000000000000000, /* 3732 */
128'h00000000000000000000000000000000, /* 3733 */
128'h00000000000000000000000000000000, /* 3734 */
128'h00000000000000000000000000000000, /* 3735 */
128'h00000000000000000000000000000000, /* 3736 */
128'h00000000000000000000000000000000, /* 3737 */
128'h00000000000000000000000000000000, /* 3738 */
128'h00000000000000000000000000000000, /* 3739 */
128'h00000000000000000000000000000000, /* 3740 */
128'h00000000000000000000000000000000, /* 3741 */
128'h00000000000000000000000000000000, /* 3742 */
128'h00000000000000000000000000000000, /* 3743 */
128'h00000000000000000000000000000000, /* 3744 */
128'h00000000000000000000000000000000, /* 3745 */
128'h00000000000000000000000000000000, /* 3746 */
128'h00000000000000000000000000000000, /* 3747 */
128'h00000000000000000000000000000000, /* 3748 */
128'h00000000000000000000000000000000, /* 3749 */
128'h00000000000000000000000000000000, /* 3750 */
128'h00000000000000000000000000000000, /* 3751 */
128'h00000000000000000000000000000000, /* 3752 */
128'h00000000000000000000000000000000, /* 3753 */
128'h00000000000000000000000000000000, /* 3754 */
128'h00000000000000000000000000000000, /* 3755 */
128'h00000000000000000000000000000000, /* 3756 */
128'h00000000000000000000000000000000, /* 3757 */
128'h00000000000000000000000000000000, /* 3758 */
128'h00000000000000000000000000000000, /* 3759 */
128'h00000000000000000000000000000000, /* 3760 */
128'h00000000000000000000000000000000, /* 3761 */
128'h00000000000000000000000000000000, /* 3762 */
128'h00000000000000000000000000000000, /* 3763 */
128'h00000000000000000000000000000000, /* 3764 */
128'h00000000000000000000000000000000, /* 3765 */
128'h00000000000000000000000000000000, /* 3766 */
128'h00000000000000000000000000000000, /* 3767 */
128'h00000000000000000000000000000000, /* 3768 */
128'h00000000000000000000000000000000, /* 3769 */
128'h00000000000000000000000000000000, /* 3770 */
128'h00000000000000000000000000000000, /* 3771 */
128'h00000000000000000000000000000000, /* 3772 */
128'h00000000000000000000000000000000, /* 3773 */
128'h00000000000000000000000000000000, /* 3774 */
128'h00000000000000000000000000000000, /* 3775 */
128'h00000000000000000000000000000000, /* 3776 */
128'h00000000000000000000000000000000, /* 3777 */
128'h00000000000000000000000000000000, /* 3778 */
128'h00000000000000000000000000000000, /* 3779 */
128'h00000000000000000000000000000000, /* 3780 */
128'h00000000000000000000000000000000, /* 3781 */
128'h00000000000000000000000000000000, /* 3782 */
128'h00000000000000000000000000000000, /* 3783 */
128'h00000000000000000000000000000000, /* 3784 */
128'h00000000000000000000000000000000, /* 3785 */
128'h00000000000000000000000000000000, /* 3786 */
128'h00000000000000000000000000000000, /* 3787 */
128'h00000000000000000000000000000000, /* 3788 */
128'h00000000000000000000000000000000, /* 3789 */
128'h00000000000000000000000000000000, /* 3790 */
128'h00000000000000000000000000000000, /* 3791 */
128'h00000000000000000000000000000000, /* 3792 */
128'h00000000000000000000000000000000, /* 3793 */
128'h00000000000000000000000000000000, /* 3794 */
128'h00000000000000000000000000000000, /* 3795 */
128'h00000000000000000000000000000000, /* 3796 */
128'h00000000000000000000000000000000, /* 3797 */
128'h00000000000000000000000000000000, /* 3798 */
128'h00000000000000000000000000000000, /* 3799 */
128'h00000000000000000000000000000000, /* 3800 */
128'h00000000000000000000000000000000, /* 3801 */
128'h00000000000000000000000000000000, /* 3802 */
128'h00000000000000000000000000000000, /* 3803 */
128'h00000000000000000000000000000000, /* 3804 */
128'h00000000000000000000000000000000, /* 3805 */
128'h00000000000000000000000000000000, /* 3806 */
128'h00000000000000000000000000000000, /* 3807 */
128'h00000000000000000000000000000000, /* 3808 */
128'h00000000000000000000000000000000, /* 3809 */
128'h00000000000000000000000000000000, /* 3810 */
128'h00000000000000000000000000000000, /* 3811 */
128'h00000000000000000000000000000000, /* 3812 */
128'h00000000000000000000000000000000, /* 3813 */
128'h00000000000000000000000000000000, /* 3814 */
128'h00000000000000000000000000000000, /* 3815 */
128'h00000000000000000000000000000000, /* 3816 */
128'h00000000000000000000000000000000, /* 3817 */
128'h00000000000000000000000000000000, /* 3818 */
128'h00000000000000000000000000000000, /* 3819 */
128'h00000000000000000000000000000000, /* 3820 */
128'h00000000000000000000000000000000, /* 3821 */
128'h00000000000000000000000000000000, /* 3822 */
128'h00000000000000000000000000000000, /* 3823 */
128'h00000000000000000000000000000000, /* 3824 */
128'h00000000000000000000000000000000, /* 3825 */
128'h00000000000000000000000000000000, /* 3826 */
128'h00000000000000000000000000000000, /* 3827 */
128'h00000000000000000000000000000000, /* 3828 */
128'h00000000000000000000000000000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00000000000000000000000000000000, /* 3840 */
128'h00000000000000000000000000000000, /* 3841 */
128'h00000000000000000000000000000000, /* 3842 */
128'h00000000000000000000000000000000, /* 3843 */
128'h00000000000000000000000000000000, /* 3844 */
128'h00000000000000000000000000000000, /* 3845 */
128'h00000000000000000000000000000000, /* 3846 */
128'h00000000000000000000000000000000, /* 3847 */
128'h00000000000000000000000000000000, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule

