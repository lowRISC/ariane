/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module etherboot (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 5959;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_bffe7042,
        64'h00000000_bffe7080,
        64'h00000000_00000000,
        64'hffffffff_00000006,
        64'h00000000_bffeb3c0,
        64'h00000000_2f7c5c2d,
        64'h00000000_ffffffff,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_cc33aa55,
        64'h00000000_bffeb208,
        64'h00006772_615f6473,
        64'h0000646d_635f6473,
        64'h00000000_0c000000,
        64'h00000000_ffffffff,
        64'h00000000_00000000,
        64'h00000000_30000000,
        64'h00000000_004b4d47,
        64'h00004b4d_47545045,
        64'h00000003_0f060301,
        64'haaaaaaaa_aaaaaaaa,
        64'h55555555_55555555,
        64'h5851f42d_4c957f2d,
        64'h10000000_20000000,
        64'h10325476_98badcfe,
        64'hefcdab89_67452301,
        64'h00000002_464c457f,
        64'hcccccccc_cccccccd,
        64'h00000a0d_70617274,
        64'h00000000_000a7473,
        64'h65742065_68636143,
        64'h00000000_00000a74,
        64'h6f6f6220_50544654,
        64'h00000000_00000a74,
        64'h73657420_4d415244,
        64'h00000000_00000a74,
        64'h6f6f6220_49505351,
        64'h00000000_00000000,
        64'h0a746f6f_62204453,
        64'h00000000_0000000a,
        64'h5825203d_20646565,
        64'h73206d6f_646e6152,
        64'h000a5825_2c582520,
        64'h3d20676e_69747465,
        64'h73206863_74697753,
        64'h0000000a_5825203d,
        64'h205d6425_5b707773,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h0a646c25_2e646c25,
        64'h203d2049_5043202c,
        64'h73656c63_79632064,
        64'h6c25202c_736e6f69,
        64'h74637572_74736e69,
        64'h20646c25_202c424b,
        64'h6425203d_20746573,
        64'h5f676e69_6b726f77,
        64'h00000000_00000000,
        64'h0a2e2979_6c6e6f28,
        64'h2032206e_6f697372,
        64'h65762065_736e6563,
        64'h694c2063_696c6275,
        64'h50206c61_72656e65,
        64'h4720554e_47206568,
        64'h74207265_646e7520,
        64'h6465736e_6563694c,
        64'h00000000_0000000a,
        64'h2e6e6f62_617a6143,
        64'h2073656c_72616843,
        64'h20323130_322d3130,
        64'h30322029_43282074,
        64'h68676972_79706f43,
        64'h00000000_0000000a,
        64'h29746962_2d642528,
        64'h20302e33_2e34206e,
        64'h6f697372_65762072,
        64'h65747365_746d656d,
        64'h00000a74_73657420,
        64'h4d415244_206c6174,
        64'h656d2065_7261420a,
        64'h00000a2e_656e6f44,
        64'h00000000_000a6b6f,
        64'h0000203a_73252020,
        64'h00000073_73657264,
        64'h6441206b_63757453,
        64'h00000000_00000a3a,
        64'h00000000_0075252f,
        64'h00752520_706f6f4c,
        64'h00000000_000a7025,
        64'h7830206f_74207025,
        64'h78302073_69206567,
        64'h6e617220_74736574,
        64'h00000000_00082008,
        64'h00000000_00000008,
        64'h08080808_08080808,
        64'h08082020_20202020,
        64'h20202020_20080808,
        64'h08080808_08080808,
        64'h00000000_0000000a,
        64'h2e2e2e74_73657420,
        64'h7478656e_206f7420,
        64'h676e6970_70696b53,
        64'h00000000_000a2e78,
        64'h25783020_74657366,
        64'h666f2074_6120656e,
        64'h696c2073_73657264,
        64'h64612064_61622065,
        64'h6c626973_736f7020,
        64'h3a455255_4c494146,
        64'h00000000_00007525,
        64'h20676e69_74736574,
        64'h00000000_00007525,
        64'h20676e69_74746573,
        64'h00000000_00080808,
        64'h08080808_08080808,
        64'h00000000_00202020,
        64'h20202020_20202020,
        64'h00000000_0000000a,
        64'h7025203d_20327020,
        64'h2c702520_3d203170,
        64'h00000a2e_78257830,
        64'h20746573_66666f20,
        64'h74612078_25783020,
        64'h3d212078_25783020,
        64'h3a455255_4c494146,
        64'h00000000_000a7325,
        64'h206e6f69_74636e75,
        64'h66202c64_2520656e,
        64'h696c202c_73252065,
        64'h6c696620_2c64656c,
        64'h69616620_7325206e,
        64'h6f697472_65737361,
        64'h00000a72_6564616f,
        64'h6c20746f_6f622065,
        64'h67617473_20747372,
        64'h69662064_65736162,
        64'h20746f6f_622d750a,
        64'h00000000_216b7369,
        64'h6420746e_756f6d75,
        64'h206f7420_6c696166,
        64'h00000000_0021656c,
        64'h69662065_736f6c63,
        64'h206f7420_6c696166,
        64'h0000000a_21746f6f,
        64'h62206e65_706f206f,
        64'h74206465_6c696146,
        64'h00000000_00000000,
        64'h6e69622e_746f6f62,
        64'h00000000_00000a79,
        64'h726f6d65_6d206f74,
        64'h6e69206e_69622e74,
        64'h6f6f6220_64616f4c,
        64'h00000000_0000000a,
        64'h21726576_69726420,
        64'h44532074_6e756f6d,
        64'h206f7420_6c696146,
        64'h00000000_0000000a,
        64'h2e2e2e70_25207373,
        64'h65726464_61207461,
        64'h206d6172_676f7270,
        64'h20646564_616f6c20,
        64'h65687420_746f6f42,
        64'h00000000_5c2d2f7c,
        64'h000a7825_203d206c,
        64'h61757463_61202c58,
        64'h25203d20_64657269,
        64'h75716572_206e656c,
        64'h00000000_00000000,
        64'h0a2e6e6f_69746172,
        64'h65706f20_50544654,
        64'h206c6167_656c6c49,
        64'h00000000_000a2e64,
        64'h656c6c61_63207172,
        64'h775f656c_646e6168,
        64'h00000000_00000a2e,
        64'h646e6520_656c6966,
        64'h20657669_65636552,
        64'h00000000_00000000,
        64'h0a64253d_657a6973,
        64'h6b636f6c_62202c22,
        64'h73252220_3a717277,
        64'h00000000_0000002f,
        64'h00000000_000a646c,
        64'h25202e67_6e6f6c20,
        64'h6f6f7420_68746170,
        64'h20747365_75716552,
        64'h00000064_6c252065,
        64'h646f6320_68746977,
        64'h2064656c_69616620,
        64'h64616572_20666c65,
        64'h000a7972_6f6d656d,
        64'h20524444_206f7420,
        64'h666c6520_64616f6c,
        64'h00000000_00000000,
        64'h0a732520_3d202964,
        64'h252c7025_2835646d,
        64'h00000000_0000000a,
        64'h6425203d_20687467,
        64'h6e656c20_656c6946,
        64'h00000000_00636d6d,
        64'h00000029_73252820,
        64'h00006425_203a7325,
        64'h00000000_434d4d65,
        64'h00000000_00004453,
        64'h00000000_00000000,
        64'h0a646e75_6f662074,
        64'h6f6e2064_25206563,
        64'h69766544_20434d4d,
        64'h0000297a_484d3030,
        64'h32282030_30325348,
        64'h00000000_00297a48,
        64'h4d383032_28203430,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282030,
        64'h35524444_20534855,
        64'h00000000_0000297a,
        64'h484d3030_31282030,
        64'h35524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282035,
        64'h32524453_20534855,
        64'h00000000_00000029,
        64'h7a484d35_32282032,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d32_35282032,
        64'h35524444_20434d4d,
        64'h0000297a_484d3235,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000029_7a484d30,
        64'h35282064_65657053,
        64'h20686769_48204453,
        64'h0000297a_484d3632,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000000_00000079,
        64'h63616765_4c204453,
        64'h00000000_00007963,
        64'h6167656c_20434d4d,
        64'h00000064_252e6425,
        64'h00000000_63256325,
        64'h63256325_63256325,
        64'h00000078_34302578,
        64'h34302520_726e5320,
        64'h78363025_206e614d,
        64'h00000000_00000a21,
        64'h646e756f_66206473,
        64'h635f7478_65206f4e,
        64'h00000000_00000000,
        64'h0a65646f_6d206120,
        64'h7463656c_6573206f,
        64'h7420656c_62616e75,
        64'h00000000_00000000,
        64'h0a217463_656c6573,
        64'h20656761_746c6f76,
        64'h206f7420_646e6f70,
        64'h73657220_746f6e20,
        64'h64696420_64726143,
        64'h0000000a_746e6573,
        64'h65727020_64726163,
        64'h206f6e20_3a434d4d,
        64'h00000000_0000000a,
        64'h64656e6f_69746974,
        64'h72617020_79646165,
        64'h726c6120_64726143,
        64'h00000000_000a7367,
        64'h6e697474_65732079,
        64'h74696c69_6261696c,
        64'h65722065_74697277,
        64'h206e6f69_74697472,
        64'h61702064_656c6c6f,
        64'h72746e6f_63207473,
        64'h6f682074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000a29_7525203e,
        64'h20752528_206d756d,
        64'h6978616d_20736465,
        64'h65637865_20657a69,
        64'h73206465_636e6168,
        64'h6e65206c_61746f54,
        64'h00000000_0000000a,
        64'h65747562_69727474,
        64'h61206465_636e6168,
        64'h6e652074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0a64656e,
        64'h67696c61_20657a69,
        64'h73207075_6f726720,
        64'h50572043_4820746f,
        64'h6e206e6f_69746974,
        64'h72617020_69255047,
        64'h0000000a_64656e67,
        64'h696c6120_657a6973,
        64'h2070756f_72672050,
        64'h57204348_20746f6e,
        64'h20616572_61206465,
        64'h636e6168_6e652061,
        64'h74616420_72657355,
        64'h00000a65_7a697320,
        64'h70756f72_67205057,
        64'h20434820_656e6966,
        64'h65642074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_000a676e,
        64'h696e6f69_74697472,
        64'h61702074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0000000a,
        64'h61657261_20617461,
        64'h64207265_73752064,
        64'h65636e61_686e6520,
        64'h726f6620_64657269,
        64'h75716572_20342e34,
        64'h203d3e20_434d4d65,
        64'h00000000_000a2978,
        64'h6c257830_2878616d,
        64'h20736465_65637865,
        64'h20786c25_78302072,
        64'h65626d75_6e206b63,
        64'h6f6c6220_3a434d4d,
        64'h00000000_00000a64,
        64'h6d632070_6f747320,
        64'h646e6573_206f7420,
        64'h6c696166_20636d6d,
        64'h00000000_000a7964,
        64'h61657220_64726163,
        64'h20676e69_74696177,
        64'h2074756f_656d6954,
        64'h0000000a_58383025,
        64'h7830203a_726f7272,
        64'h45207375_74617453,
        64'h00000000_65646f6d,
        64'h206e776f_6e6b6e55,
        64'h00000000_00006473,
        64'h5f637369_72776f6c,
        64'h00000078_25782520,
        64'h00000020_3a78250a,
        64'h00000000_0a732574,
        64'h69622d64_25203a68,
        64'h74646957_20737542,
        64'h00000000_0000203a,
        64'h79746963_61706143,
        64'h00000000_00000a73,
        64'h25203a79_74696361,
        64'h70614320_68676948,
        64'h00000a64_25203a64,
        64'h65657053_20737542,
        64'h00000000_00000a20,
        64'h63256325_63256325,
        64'h6325203a_656d614e,
        64'h00000000_00000000,
        64'h0a782520_3a4d454f,
        64'h00000000_0a782520,
        64'h3a444920_72657275,
        64'h74636166_756e614d,
        64'h00000000_000a7325,
        64'h203a6563_69766544,
        64'h00202020_3a434d4d,
        64'h00000000_52444420,
        64'h00000000_00006f4e,
        64'h00000000_00736559,
        64'h0000000a_7825203d,
        64'h2074736f_68202c78,
        64'h25207461_20646574,
        64'h61657263_20636d6d,
        64'h00000000_00000a64,
        64'h25206f74_20646567,
        64'h6e616863_206b7361,
        64'h6d202c64_65747265,
        64'h736e6920_64726143,
        64'h00000000_0000000a,
        64'h6425206f_74206465,
        64'h676e6168_63206b73,
        64'h616d202c_6465766f,
        64'h6d657220_64726143,
        64'h000a7475_6f656d69,
        64'h74207325_203a6473,
        64'h5f637369_72776f6c,
        64'h00726464_615f6573,
        64'h61625f64_73203d3d,
        64'h20657361_625f6473,
        64'h00000000_00000063,
        64'h2e636d6d_5f637369,
        64'h72776f6c_2f637273,
        64'h00000000_00000000,
        64'h66656463_62613938,
        64'h37363534_33323130,
        64'h007f7c5d_5b3f3e3d,
        64'h3c3b3a2e_2c2b2a22,
        64'h00007f7c_5d5b3f3e,
        64'h3d3c3b3a_2c2b2a22,
        64'h0000000a_2e783230,
        64'h253a7832_30253a78,
        64'h3230253a_78323025,
        64'h3a783230_253a7832,
        64'h3025203d_20737365,
        64'h72646461_2043414d,
        64'h00000a78_6c253a78,
        64'h6c25203d_2043414d,
        64'h00000000_00000a78,
        64'h25203d20_5d64255b,
        64'h4d454f20_49505351,
        64'h000a7264_64612043,
        64'h414d2070_75746553,
        64'h0000000a_21747075,
        64'h72726574_6e692064,
        64'h656c646e_61686e75,
        64'h00000000_00000a78,
        64'h25783020_3d206570,
        64'h79745f6f_746f7270,
        64'h00000000_0a297825,
        64'h28206465_74726f70,
        64'h7075736e_75203d20,
        64'h6f746f72_70205049,
        64'h000a5741_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a534c50_4d203d20,
        64'h6f746f72_50205049,
        64'h00000000_000a4554,
        64'h494c5044_55203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505443_53203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a504d4f_43203d20,
        64'h6f746f72_50205049,
        64'h00000000_0000004d,
        64'h00000000_0000000a,
        64'h5041434e_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000a48,
        64'h50544545_42203d20,
        64'h6f746f72_50205049,
        64'h000a5054_4d203d20,
        64'h6f746f72_50205049,
        64'h00000a48_41203d20,
        64'h6f746f72_50205049,
        64'h000a5053_45203d20,
        64'h6f746f72_50205049,
        64'h000a4552_47203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505653_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000036,
        64'h00000000_00000000,
        64'h0a504343_44203d20,
        64'h6f746f72_50205049,
        64'h00000a50_54203d20,
        64'h6f746f72_50205049,
        64'h000a5044_49203d20,
        64'h6f746f72_50205049,
        64'h000a3a73_746e6574,
        64'h6e6f6320_74736574,
        64'h0000000a_3a726564,
        64'h61656820_74736574,
        64'h000a5055_50203d20,
        64'h6f746f72_50205049,
        64'h000a5047_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000054,
        64'h00000000_00000000,
        64'h0a504950_49203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000047,
        64'h00006425_2b544553,
        64'h46464f5f_524c5052,
        64'h00000000_3f3f3f3f,
        64'h00000000_00544553,
        64'h46464f5f_524c5052,
        64'h00000000_00544553,
        64'h46464f5f_44414252,
        64'h00000000_00005445,
        64'h5346464f_5f525352,
        64'h00000000_00544553,
        64'h46464f5f_53434652,
        64'h00544553_46464f5f,
        64'h4c525443_4f49444d,
        64'h00000000_00544553,
        64'h46464f5f_53434654,
        64'h00000000_00544553,
        64'h46464f5f_524c5054,
        64'h00000000_54455346,
        64'h464f5f49_4843414d,
        64'h00000000_54455346,
        64'h464f5f4f_4c43414d,
        64'h00000000_000a3b29,
        64'h78257830_2c302c78,
        64'h25287465_736d656d,
        64'h00000000_0a3b2978,
        64'h2578302c_78257830,
        64'h2c782528_6e666c65,
        64'h00000a70_2520726f,
        64'h72726520_7974696e,
        64'h61732072_64646170,
        64'h00000020_3a5d6425,
        64'h5b6e6f69_74636553,
        64'h000a7325_20202020,
        64'h00786c6c_2a302520,
        64'h00003a78_6c383025,
        64'h00732542_69632520,
        64'h00000000_00732573,
        64'h65747942_20756c25,
        64'h0073257a_48632520,
        64'h00000000_646c252e,
        64'h00000000_00756c25,
        64'h00000000_00000000,
        64'h73257a48_20756c25,
        64'h00000000_00007325,
        64'h00000000_00732520,
        64'h3a646c69_7542202c,
        64'h00000000_73257325,
        64'h00000000_00000a0a,
        64'h00000058_32302520,
        64'h00000000_0000002e,
        64'h00000000_00006325,
        64'h00000000_00000020,
        64'h20202020_20202020,
        64'h000a5245_46464f5f,
        64'h50434844_20726f66,
        64'h20676e69_74696157,
        64'h00000a73_25203a73,
        64'h25206563_69766564,
        64'h206e6f20_59524556,
        64'h4f435349_44205043,
        64'h48442064_6e657320,
        64'h74276e64_6c756f43,
        64'h000a5832_30253a58,
        64'h3230253a_58323025,
        64'h3a583230_253a5832,
        64'h30253a58_32302520,
        64'h3a204341_4d207325,
        64'h00000000_30687465,
        64'h00000000_000a2973,
        64'h2528726f_72726570,
        64'h000a5952_45564f43,
        64'h5349445f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_0000000a,
        64'h64252065_646f6370,
        64'h6f205043_48442064,
        64'h656c646e_61686e55,
        64'h00000000_0a642520,
        64'h6e6f6974_706f2064,
        64'h656c646e_61686e75,
        64'h00000000_0000000a,
        64'h73252072_6f727245,
        64'h00000000_00000a64,
        64'h65737566_65722073,
        64'h73657264_64612064,
        64'h65747365_75716552,
        64'h00000000_0000000a,
        64'h4b414e20_50434844,
        64'h00000000_0a444550,
        64'h50494b53_204b4341,
        64'h000a2273_2522203d,
        64'h20656d61_6e74736f,
        64'h4820746e_65696c43,
        64'h00000a22_73252220,
        64'h3d206e69_616d6f44,
        64'h00000000_0000000a,
        64'h7364253a_6d64253a,
        64'h68642520_3d20656d,
        64'h69742065_7361654c,
        64'h000a6425_2e64252e,
        64'h64252e64_2520203a,
        64'h73736572_64646120,
        64'h6b73616d_2074654e,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h61207265_74756f52,
        64'h00000000_00000000,
        64'h0a64252e_64252e64,
        64'h252e6425_20203a73,
        64'h73657264_64412050,
        64'h49207265_76726553,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h41205049_20746e65,
        64'h696c4320_50434844,
        64'h00000000_0000000a,
        64'h4b434120_50434844,
        64'h0000000a_54534555,
        64'h5145525f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_00000000,
        64'h0a702520_2c726f72,
        64'h7265206c_616e7265,
        64'h746e6920_70636864,
        64'h00000a29_73252c73,
        64'h25287075_6b6f6f6c,
        64'h000a6563_69766564,
        64'h206e776f_6e6b6e75,
        64'h00000000_203a6425,
        64'h20656369_7665440a,
        64'h00203a64_25206563,
        64'h69766564_2073250a,
        64'h00000000_00203a64,
        64'h25206563_69766544,
        64'h00000000_00000000,
        64'h73736572_6464612d,
        64'h63616d2d_6c61636f,
        64'h6c006874_6469772d,
        64'h6f692d67_65720074,
        64'h66696873_2d676572,
        64'h00737470_75727265,
        64'h746e6900_746e6572,
        64'h61702d74_70757272,
        64'h65746e69_00646565,
        64'h70732d74_6e657272,
        64'h75630076_65646e2c,
        64'h76637369_72007974,
        64'h69726f69_72702d78,
        64'h616d2c76_63736972,
        64'h0073656d_616e2d67,
        64'h65720064_65646e65,
        64'h7478652d_73747075,
        64'h72726574_6e690073,
        64'h65676e61_7200656c,
        64'h646e6168_702c7875,
        64'h6e696c00_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h00100000_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_00000064,
        64'h6e727768_2d637369,
        64'h72776f6c_1b000000,
        64'h0e000000_03000000,
        64'h00003030_30303030,
        64'h30344064_6e727768,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h00800000_00000000,
        64'h00000030_00000000,
        64'h67000000_10000000,
        64'h03000000_00007fe3,
        64'h023e1800_47010000,
        64'h06000000_03000000,
        64'h03000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_00636d6d,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_02000000,
        64'h25010000_04000000,
        64'h03000000_02000000,
        64'h14010000_04000000,
        64'h03000000_00000100,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40636d6d,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h04000000_3a010000,
        64'h04000000_03000000,
        64'h02000000_30010000,
        64'h04000000_03000000,
        64'h01000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h00c20100_06010000,
        64'h04000000_03000000,
        64'h80f0fa02_4b000000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000010_00000000,
        64'h67000000_10000000,
        64'h03000000_00303537,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000000,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'hffff0000_01000000,
        64'hca000000_08000000,
        64'h03000000_00333130,
        64'h2d677562_65642c76,
        64'h63736972_1b000000,
        64'h10000000_03000000,
        64'h00003040_72656c6c,
        64'h6f72746e_6f632d67,
        64'h75626564_01000000,
        64'h02000000_02000000,
        64'hbb000000_04000000,
        64'h03000000_02000000,
        64'hb5000000_04000000,
        64'h03000000_03000000,
        64'hfb000000_04000000,
        64'h03000000_07000000,
        64'he8000000_04000000,
        64'h03000000_00000004,
        64'h00000000_0000000c,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h09000000_01000000,
        64'h0b000000_01000000,
        64'hca000000_10000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00000c00,
        64'h00000000_00000002,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_01000000,
        64'h03000000_01000000,
        64'hca000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6e696c63,
        64'h01000000_c3000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h01000000_bb000000,
        64'h04000000_03000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00007663_73697200,
        64'h656e6169_7261202c,
        64'h7a687465_1b000000,
        64'h13000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha8060000_59010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'he0060000_38000000,
        64'h39080000_edfe0dd0,
        64'h00000000_fffff9da,
        64'hfffff9a0_fffff9c8,
        64'hfffff9a0_fffff9b6,
        64'hfffff9a2_fffff98e,
        64'h00000000_64726143,
        64'h2d445320_726f6620,
        64'h746f6f62_2d752064,
        64'h6573696d_696e696d,
        64'h20435349_52776f4c,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00020000_00010000,
        64'h0000c000_00008000,
        64'h00006000_00004000,
        64'h00002000_00001000,
        64'h00000800_00000400,
        64'h00000200_00000100,
        64'h00000080_00000040,
        64'h00000020_00000000,
        64'h0bebc200_0c65d400,
        64'h02faf080_05f5e100,
        64'h02faf080_017d7840,
        64'h03197500_03197500,
        64'h02faf080_018cba80,
        64'h017d7840_017d7840,
        64'h00989680_000f4240,
        64'h000186a0_00002710,
        64'h50463c37_322d2823,
        64'h1e19140f_0d0c0a00,
        64'h00000000_00000000,
        64'h00000000_10000000,
        64'h00000001_00000000,
        64'h20000000_00000002,
        64'h00000000_40000000,
        64'h00000005_00000001,
        64'h20000000_00000006,
        64'h00000001_40000000,
        64'h70000000_00000000,
        64'h70000000_00000002,
        64'h70000000_00000004,
        64'h60000000_00000005,
        64'h30000000_00000001,
        64'h30000000_00000003,
        64'h00000000_40050100,
        64'h40050000_40040500,
        64'h40040401_40040400,
        64'h40040300_40040200,
        64'h40040100_40040000,
        64'h00000000_bffeb370,
        64'h00000000_bffeb358,
        64'h00000000_bffeb340,
        64'h00000000_bffeb328,
        64'h00000000_bffeb310,
        64'h00000000_bffeb2f8,
        64'h00000000_bffeb2e0,
        64'h00000000_bffeb2c8,
        64'h00000000_bffeb2b0,
        64'h00000000_bffeb298,
        64'h00000000_bffeb288,
        64'h00000000_bffeb278,
        64'hffffcb68_ffffcb62,
        64'hffffcb5c_ffffc9b8,
        64'hffffbb46_ffffbb46,
        64'hffffbb46_ffffbb46,
        64'hffffbb42_ffffbb3e,
        64'hffffbb3e_ffffbb1a,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_bffe4cc6,
        64'h00000000_bffe4a68,
        64'h00000000_bffe4e58,
        64'h00646374_65675f63,
        64'h6d6d5f64_72616f62,
        64'h00000002_0000ffff,
        64'h004c4b40_004c4b40,
        64'h00300000_20000000,
        64'h00000000_bffe9c88,
        64'h00000000_bffeaf60,
        64'h00717269_5f646e65,
        64'h5f617461_645f6473,
        64'h5f637369_72776f6c,
        64'h00000000_00007172,
        64'h695f646d_635f6473,
        64'h5f637369_72776f6c,
        64'h00007172_695f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0067616c,
        64'h665f7470_75727265,
        64'h746e695f_74696177,
        64'h5f637369_72776f6c,
        64'h00000000_646d635f,
        64'h74726174_735f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0000006e,
        64'h655f7172_695f6473,
        64'h00000000_00007475,
        64'h6f656d69_745f6473,
        64'h00000000_0000657a,
        64'h69736b6c_625f6473,
        64'h00000000_00000074,
        64'h6e636b6c_625f6473,
        64'h00000000_00000000,
        64'h74657365_725f6473,
        64'h00000000_74726174,
        64'h735f646d_635f6473,
        64'h00000000_0000676e,
        64'h69747465_735f6473,
        64'h00000000_00007669,
        64'h645f6b6c_635f6473,
        64'h00000000_00000000,
        64'h6e67696c_615f6473,
        64'h00000000_00006465,
        64'h6c5f7465_735f6473,
        64'h5f637369_72776f6c,
        64'h09020b04_0d060f08,
        64'h010a030c_050e0700,
        64'h020f0c09_0603000d,
        64'h0a070401_0e0b0805,
        64'h0c07020d_08030e09,
        64'h040f0a05_000b0601,
        64'heb86d391_2ad7d2bb,
        64'hbd3af235_f7537e82,
        64'h4e0811a1_a3014314,
        64'hfe2ce6e0_6fa87e4f,
        64'h85845dd1_ffeff47d,
        64'h8f0ccc92_655b59c3,
        64'hfc93a039_ab9423a7,
        64'h432aff97_f4292244,
        64'hc4ac5665_1fa27cf8,
        64'he6db99e5_d9d4d039,
        64'h04881d05_d4ef3085,
        64'heaa127fa_289b7ec6,
        64'hbebfbc70_f6bb4b60,
        64'h4bdecfa9_a4beea44,
        64'hfde5380c_6d9d6122,
        64'h8771f681_fffa3942,
        64'h8d2a4c8a_676f02d9,
        64'hfcefa3f8_a9e3e905,
        64'h455a14ed_f4d50d87,
        64'hc33707d6_21e1cde6,
        64'he7d3fbc8_d8a1e681,
        64'h02441453_d62f105d,
        64'he9b6c7aa_265e5a51,
        64'hc040b340_f61e2562,
        64'h49b40821_a679438e,
        64'hfd987193_6b901122,
        64'h895cd7be_ffff5bb1,
        64'h8b44f7af_698098d8,
        64'hfd469501_a8304613,
        64'h4787c62a_f57c0faf,
        64'hc1bdceee_242070db,
        64'he8c7b756_d76aa478,
        64'h02020202_02020202,
        64'h10020202_02020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02010101_01010101,
        64'h10010101_01010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h08101010_10020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02424242_42424210,
        64'h10101010_10010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h01414141_41414110,
        64'h10101010_10100404,
        64'h04040404_04040404,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h08080808_08080808,
        64'h08080808_08080808,
        64'h08082828_28282808,
        64'h08080808_08080808,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_bf5dcfdf,
        64'hf0efedff_b0ef0ae5,
        64'h05130000_2517b7e1,
        64'hde2f80ef_ef1fb0ef,
        64'h0b050513_00002517,
        64'hbfe9c25f_f0eff03f,
        64'hb0ef0b25_05130000,
        64'h2517b7f5_edbff0ef,
        64'h8522f17f_b0ef0b65,
        64'h05130000_2517a001,
        64'hac3fe0ef_8522f2bf,
        64'hb0ef0ba5_05130000,
        64'h25178782_97ba439c,
        64'h97ba078a_68470713,
        64'h00000717_02f76463,
        64'h47190054_579b0ff4,
        64'h7413fd39_1be3f5bf,
        64'hb0ef2581_8552688c,
        64'h0004b823_f69fb0ef,
        64'h86222401_25816080,
        64'h608ce09c_09058556,
        64'h0007c783_016907b3,
        64'h49910faa_0a130000,
        64'h2a170eaa_8a930000,
        64'h2a974000_04b720eb,
        64'h0b130000_2b174901,
        64'hdb4f80ef_fe9416e3,
        64'hfadfb0ef_0405854a,
        64'h0004059b_639097ce,
        64'h00341793_449510e9,
        64'h09130000_29174000,
        64'h09b74401_94ffe0ef,
        64'h11050513_00002517,
        64'h929fe0ef_e05ae456,
        64'he852ec4e_f04af426,
        64'hf822fc06_7139971f,
        64'he06f1d25_05130000,
        64'h2517b69f_e06f0141,
        64'h60a2806f_c06f0141,
        64'hcc050513_00002517,
        64'h40a005b3_60a20005,
        64'h5c63d51f_70eff7c5,
        64'h05130000_051782af,
        64'hc0efe406_ccc50513,
        64'h00002517_1141bf4d,
        64'h008bb023_0921f3bf,
        64'hf0ef00c4_541b85ce,
        64'h24218082_61256be2,
        64'h7b027aa2_7a4279e2,
        64'h690664a6_644660e6,
        64'hed3fd0ef_9201854e,
        64'h002c1602_4084863b,
        64'hf6dff0ef_002c0344,
        64'h6863008a_853b012b,
        64'h09b30009_041b4000,
        64'h0bb7ff86_0a1b4901,
        64'h84b28aae_8b2afc4e,
        64'he8a2ec86_ec5ef05a,
        64'hf456f852_e0cae4a6,
        64'h711d8082_61056442,
        64'h60e2fee7_9ae30585,
        64'h37e100d5_802300f5,
        64'h56b35761_03800793,
        64'h85a2f49f_f0ef454d,
        64'h46010034_4589f55f,
        64'hf0efec06_c43e454d,
        64'h45894601_0034842e,
        64'hc62ae822_8fd90585,
        64'h65133007_07131101,
        64'h0085151b_67050185,
        64'h579b9d3d_00b007b7,
        64'ha45fe06f_014160a2,
        64'h64020004_4503943e,
        64'h24078793_00002797,
        64'h883dfedf_f0ef0045,
        64'h551b35fd_00b7d763,
        64'h842a4785_e406e022,
        64'h1141bfc1_f6180785,
        64'h00076703_97360027,
        64'h97138082_73884000,
        64'h07b7ffe5_37fdc319,
        64'h8b097a98_400006b7,
        64'h3e800793_00b76f63,
        64'h0007871b_40000637,
        64'h47812581_f7884000,
        64'h07b78d51_0106161b,
        64'h8d5d0085_979b8082,
        64'h25017b88_400007b7,
        64'h80822501_6b880007,
        64'hb8234000_07b78082,
        64'h25016388_400007b7,
        64'h8082e388_400007b7,
        64'h91011502_bff1f5df,
        64'hf0ef4541_f63ff0ef,
        64'h4521f69f_f0ef4511,
        64'hf6fff0ef_4509f75f,
        64'hf0ef4505_f7bff0ef,
        64'h4501e406_1141bf51,
        64'hc00028f3_c02026f3,
        64'hfac710e3_9f0fc06f,
        64'h2d050513_00002517,
        64'h02a74733_02a767b3,
        64'h02b345bb_02c74733,
        64'h40000593_02a68733,
        64'h411686b3_3e800513,
        64'hc00026f3_8e15c020,
        64'h267302b7_1d632705,
        64'hfe0813e3_97aa387d,
        64'h00078023_97aa0007,
        64'h802397aa_00078023,
        64'h97aa0007_80234000,
        64'h081387f2_45a901f6,
        64'h1e134681_48814701,
        64'h00c5131b_46058082,
        64'h80826145_69a26942,
        64'h64e27402_70a2ff24,
        64'h17e3e73f_f0ef2405,
        64'h01358533_46054685,
        64'h008495b3_497901f4,
        64'h99934441_a90fc0ef,
        64'h44850725_05130000,
        64'h2517a9ef_c0ef3365,
        64'h05130000_2517aaaf,
        64'hc0ef3125_05130000,
        64'h2517ab6f_c0ef2f65,
        64'h05130000_25170400,
        64'h0593c45f_e0efe44e,
        64'he84aec26_f022f406,
        64'h2f850513_00002517,
        64'h7179bf89_0485ae2f,
        64'hc0ef0c25_05130000,
        64'h2517b7d1_4a89af2f,
        64'hc0ef30a5_05130000,
        64'h25179782_852295a2,
        64'h00495613_00195593,
        64'h008a3783_b10fc0ef,
        64'h32050513_00002517,
        64'hc985000a_358302f7,
        64'h4c636722_010a2783,
        64'hb2cfc0ef_856ee129,
        64'h952ff0ef_85226582,
        64'hb3cfc0ef_856a85e6,
        64'hb44fc0ef_8562b4af,
        64'hc0ef855e_85ce0009,
        64'h8663b56f_c0ef855a,
        64'h85a68082_61096de2,
        64'h7d027ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_85567446,
        64'h70e6b7ef_c0ef39e5,
        64'h05130000_25170299,
        64'hf863eaaa_0a130000,
        64'h3a173aad_8d930000,
        64'h2d973aad_0d130000,
        64'h2d173a2c_8c930000,
        64'h2c973a2c_0c130000,
        64'h2c173a2b_8b930000,
        64'h2b973a2b_0b130000,
        64'h2b174485_4a81e03e,
        64'h00395793_bd0fc0ef,
        64'he436fc86_ec6ef06a,
        64'hf466f862_fc5ee0da,
        64'he4d6e8d2_f4a63ae5,
        64'h05130000_251785aa,
        64'h842a892e_962af0ca,
        64'hf8a2fff5_861389b2,
        64'hecce7119_80826505,
        64'hbfb1547d_bf050d85,
        64'he99fe0ef_0007c503,
        64'h97ea8b8d_00078b1b,
        64'h001b079b_eadfe0ef,
        64'h4521ef91_0ba1033d,
        64'hf7b3ff97_95e300d6,
        64'h102392c1_16c20789,
        64'h00fb8633_0006d683,
        64'h018786b3_4781e288,
        64'hf8a7b823_00003797,
        64'h8d4166e2_91011402,
        64'h15028c51_0106161b,
        64'h8d5d0105_151b6642,
        64'h67a2fe3f_d0efe42a,
        64'hfe9fd0ef_e82afeff,
        64'hd0ef842a_ff5fd0ef,
        64'hec36b775_4a058082,
        64'h61497da2_7d427ce2,
        64'h6c066ba6_6b466ae6,
        64'h7a0679a6_794674e6,
        64'h640a60aa_8522cb2f,
        64'hc0ef4725_05130000,
        64'h251702fa_18638aa6,
        64'h8bca4785_ed4d842a,
        64'ha94ff0ef_854a85a6,
        64'h866e04fd_966396d6,
        64'h003d9693_67824d81,
        64'h790d0d13_00002d17,
        64'h9c498993_4ca102ec,
        64'h0c130000_3c174b01,
        64'h4a098ba6_f85fe0ef,
        64'h8acae032_f46ee122,
        64'he506f86a_fc66e0e2,
        64'he4dee8da_ecd6f0d2,
        64'h69850200_051384ae,
        64'h892af4ce_f8cafca6,
        64'h7175bfb1_547dbf05,
        64'h0d85fbbf_e0ef0007,
        64'hc50397ea_8b8d0007,
        64'h8b1b001b_079bfcff,
        64'he0ef4521_ef910ba1,
        64'h033df7b3_ff9795e3,
        64'h00d60023_0ff6f693,
        64'h078500fb_86330006,
        64'hc6830187_86b34781,
        64'he2880aa7_b5230000,
        64'h37978d41_66e29101,
        64'h14021502_8c510106,
        64'h161b8d5d_0105151b,
        64'h664267a2_904fe0ef,
        64'he42a90af_e0efe82a,
        64'h910fe0ef_842a916f,
        64'he0efec36_b7754a05,
        64'h80826149_7da27d42,
        64'h7ce26c06_6ba66b46,
        64'h6ae67a06_79a67946,
        64'h74e6640a_60aa8522,
        64'hdd4fc0ef_59450513,
        64'h00002517_02fa1863,
        64'h8aa68bca_4785ed4d,
        64'h842abb6f_f0ef854a,
        64'h85a6866e_04fd9663,
        64'h96d6003d_96936782,
        64'h4d818b2d_0d130000,
        64'h3d179c49_89934ca1,
        64'h148c0c13_00003c17,
        64'h4b014a09_8ba68a6f,
        64'hf0ef8aca_e032f46e,
        64'he122e506_f86afc66,
        64'he0e2e4de_e8daecd6,
        64'hf0d26985_02000513,
        64'h84ae892a_f4cef8ca,
        64'hfca67175_b7e95b7d,
        64'hb7490605_00b83023,
        64'he30c85d6_e11185e2,
        64'h00167513_80826109,
        64'h6de27d02_7ca27c42,
        64'h7be26b06_6aa66a46,
        64'h69e67906_74a6855a,
        64'h744670e6_e88fc0ef,
        64'h62050513_00002517,
        64'hfafb90e3_04000793,
        64'h2b85fbb4_1be38c56,
        64'h2405e931_8b2ac72f,
        64'hf0ef854a_85ce6622,
        64'heb4fc0ef_856a85da,
        64'hebcfc0ef_e4328552,
        64'h06f61063_974e00e9,
        64'h08330036_17136782,
        64'h4601fffc_4a93edaf,
        64'hc0ef8566_85da0084,
        64'h8b3bee6f_c0ef8552,
        64'h4401003b_949b0177,
        64'h9c334785_4da1626d,
        64'h0d130000_2d1761ec,
        64'h8c930000_2c97616a,
        64'h0a130000_2a17f12f,
        64'hc0ef4b81_e03289ae,
        64'hf862e0da_e4d6f4a6,
        64'hf8a2fc86_ec6ef06a,
        64'hf466fc5e_e8d2ecce,
        64'h63050513_00002517,
        64'h892af0ca_7119bf75,
        64'h5dfdbfc5_859afe08,
        64'h0be385ba_b7610605,
        64'he10ce28c_85c60008,
        64'h036385be_008bea63,
        64'h00167813_80826109,
        64'h6de27d02_7ca27c42,
        64'h7be26b06_6aa66a46,
        64'h69e67906_74a6856e,
        64'h744670e6_f88fc0ef,
        64'h72050513_00002517,
        64'hf8f41be3_08000793,
        64'h2405ed29_8daad6af,
        64'hf0ef8526_85ca6622,
        64'hfacfc0ef_856685a2,
        64'hfb4fc0ef_e432854e,
        64'h05461c63_96ca00d4,
        64'h85330036_16934601,
        64'hfff7c893_fff74313,
        64'h8fd5008d_16b300fd,
        64'h17b30024_079b8f5d,
        64'h00ed1733_00fd17b3,
        64'h408b07bb_408a873b,
        64'hff4fc0ef_856285a2,
        64'hffcfc0ef_854e72ec,
        64'h8c930000_2c9703f0,
        64'h0b930810_0b134d05,
        64'h07f00a93_734c0c13,
        64'h00002c17_72c98993,
        64'h00002997_829fc0ef,
        64'h44018a32_892eec6e,
        64'hfc86f06a_f466f862,
        64'hfc5ee0da_e4d6e8d2,
        64'heccef0ca_f8a27465,
        64'h05130000_251784aa,
        64'hf4a67119_b7f15dfd,
        64'hbfe5e19c_e31cbf61,
        64'h0605e194_e314008c,
        64'h66638082_61096de2,
        64'h7d027ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_856e7446,
        64'h70e688ff_c0ef8265,
        64'h05130000_3517fb54,
        64'h17e32405_e1398daa,
        64'he6cff0ef_852685ca,
        64'h66228aff_c0ef856a,
        64'h85a28b7f_c0efe432,
        64'h85520566_1a63974a,
        64'h00e485b3_00361713,
        64'h4601fff6_c693fff7,
        64'hc7930089_96b300f9,
        64'h97b3408b_87bb8e3f,
        64'hc0ef8566_85a28ebf,
        64'hc0ef8552_08000a93,
        64'h820d0d13_00003d17,
        64'h03f00c13_498507f0,
        64'h0b93822c_8c930000,
        64'h3c9781aa_0a130000,
        64'h3a17917f_c0ef4401,
        64'h8b32892e_ec6efc86,
        64'hf06af466_f862fc5e,
        64'he0dae4d6_e8d2ecce,
        64'hf0caf8a2_83450513,
        64'h00003517_84aaf4a6,
        64'h7119b7f1_5dfdbfe5,
        64'he298e398_bf610605,
        64'he28ce38c_008c6663,
        64'h80826109_6de27d02,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e67906,
        64'h74a6856e_744670e6,
        64'h97dfc0ef_91450513,
        64'h00003517_fb541be3,
        64'h2405e139_8daaf5af,
        64'hf0ef8526_85ca6622,
        64'h99dfc0ef_856a85a2,
        64'h9a5fc0ef_e4328552,
        64'h05661a63_97ca00f4,
        64'h86b30036_17934601,
        64'h008995b3_00e99733,
        64'h408b873b_9c9fc0ef,
        64'h856685a2_9d1fc0ef,
        64'h85520800_0a93906d,
        64'h0d130000_3d1703f0,
        64'h0c134985_07f00b93,
        64'h908c8c93_00003c97,
        64'h900a0a13_00003a17,
        64'h9fdfc0ef_44018b32,
        64'h892eec6e_fc86f06a,
        64'hf466f862_fc5ee0da,
        64'he4d6e8d2_eccef0ca,
        64'hf8a291a5_05130000,
        64'h351784aa_f4a67119,
        64'hbff159fd_b74d0605,
        64'he29ce31c_80826125,
        64'h6c426be2_7b027aa2,
        64'h7a4279e2_690664a6,
        64'h854e6446_60e6a53f,
        64'hc0ef9ea5_05130000,
        64'h3517f94c_19e30c05,
        64'he91d89aa_831ff0ef,
        64'h852285a6_6622a73f,
        64'hc0ef855e_85cea7bf,
        64'hc0efe432_854a0556,
        64'h17639726_00e406b3,
        64'h00361713_46018fd9,
        64'h038c1713_8fd9030c,
        64'h17138fd9_028c1713,
        64'h8fd9020c_17138fd9,
        64'h018c1713_0187e7b3,
        64'h8fd9008c_1793010c,
        64'h1713abff_c0ef855a,
        64'h85ce000c_099bacbf,
        64'hc0ef854a_10000a13,
        64'ha00b8b93_00003b97,
        64'h9f8b0b13_00003b17,
        64'h9f090913_00003917,
        64'haedfc0ef_4c018ab2,
        64'h84aefc4e_ec86e862,
        64'hec5ef05a_f456f852,
        64'he0cae4a6_a0450513,
        64'h00003517_842ae8a2,
        64'h711db7e1_5d7db779,
        64'h0605e198_e398872a,
        64'hc291876a_00167693,
        64'hbf49000b_3d038082,
        64'h61656d42_6ce27c02,
        64'h7ba27b42_7ae26a06,
        64'h69a66946_64e6856a,
        64'h740670a6_b51fc0ef,
        64'hae850513_00003517,
        64'hfb441ae3_2405e529,
        64'h8d2a92ff_f0ef8526,
        64'h85ca6622_b71fc0ef,
        64'h856685a2_b79fc0ef,
        64'he432854e_05561c63,
        64'h97ca00f4_85b30036,
        64'h1793fffd_45134601,
        64'hb95fc0ef_856285a2,
        64'h000bbd03_cba50014,
        64'h7793ba7f_c0ef854e,
        64'h04000a13_adcc8c93,
        64'h00003c97_ad4c0c13,
        64'h00003c17_ddcb8b93,
        64'h00003b97_ddcb0b13,
        64'h00003b17_adc98993,
        64'h00003997_bd9fc0ef,
        64'h44018ab2_892ee86a,
        64'hf486ec66_f062f45e,
        64'hf85afc56_e0d2e4ce,
        64'he8caf0a2_af450513,
        64'h00003517_84aaeca6,
        64'h7159bfc1_54fdbf59,
        64'h0605e198_e3988726,
        64'hc2918766_00167693,
        64'h80826165_6ce27c02,
        64'h7ba27b42_7ae26a06,
        64'h69a664e6_69468526,
        64'h740670a6_c39fc0ef,
        64'hbd050513_00003517,
        64'hfb541be3_2405e129,
        64'h84aaa17f_f0ef854a,
        64'h85ce6622_c59fc0ef,
        64'h856285a2_c61fc0ef,
        64'he4328552_05661863,
        64'h97ce00f9_05b30036,
        64'h179314fd_46014090,
        64'h0cb3c7ff_c0ef8885,
        64'h855e85a2_fff44493,
        64'hc8dfc0ef_85520400,
        64'h0a93bc2c_0c130000,
        64'h3c17bbab_8b930000,
        64'h3b97bb2a_0a130000,
        64'h3a17caff_c0ef4401,
        64'h8b3289ae_ec66eca6,
        64'hf486f062_f45ef85a,
        64'hfc56e0d2_e4cef0a2,
        64'hbc850513_00003517,
        64'h892ae8ca_7159bfc9,
        64'h070500a8_3023e288,
        64'h00f70533_ab1ff06f,
        64'h6121863a_69e2854e,
        64'h790274a2_70e27442,
        64'h00c71c63_96ae00d9,
        64'h88330037_16934701,
        64'h8fc59081_178265a2,
        64'h66021482_8fc18cc9,
        64'h0109179b_0105151b,
        64'h891fe0ef_84aa897f,
        64'he0ef892a_89dfe0ef,
        64'h842a8a3f_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7f100e8_30238f69,
        64'h00083703_e3148ee9,
        64'h07856314_b29ff06f,
        64'h6121863e_69e2854e,
        64'h790274a2_70e27442,
        64'h00c79c63_974e00e5,
        64'h88330037_97134781,
        64'h8d5d9101_178265a2,
        64'h66021502_8fc18d45,
        64'h0109179b_0105151b,
        64'h909fe0ef_84aa90ff,
        64'he0ef892a_915fe0ef,
        64'h842a91bf_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7f100e8_30238f49,
        64'h00083703_e3148ec9,
        64'h07856314_ba1ff06f,
        64'h6121863e_69e2854e,
        64'h790274a2_70e27442,
        64'h00c79c63_974e00e5,
        64'h88330037_97134781,
        64'h8d5d9101_178265a2,
        64'h66021502_8fc18d45,
        64'h0109179b_0105151b,
        64'h981fe0ef_84aa987f,
        64'he0ef892a_98dfe0ef,
        64'h842a993f_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7d100e8_302302a7,
        64'h57330008_3703e314,
        64'h02a6d6b3_07856314,
        64'h4505e111_c21ff06f,
        64'h6121863e_69e2854e,
        64'h790274a2_70e27442,
        64'h00c79c63_974e00e5,
        64'h88330037_97134781,
        64'h8d5d9101_178265a2,
        64'h66021502_8fc18d45,
        64'h0109179b_0105151b,
        64'ha01fe0ef_84aaa07f,
        64'he0ef892a_a0dfe0ef,
        64'h842aa13f_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7e100e8_302302a7,
        64'h07330008_3703e314,
        64'h02a686b3_07856314,
        64'hc9dff06f_6121863e,
        64'h69e2854e_790274a2,
        64'h70e27442_00c79c63,
        64'h974e00e5_88330037,
        64'h97134781_8d5d9101,
        64'h178265a2_66021502,
        64'h8fc18d45_0109179b,
        64'h0105151b_a7dfe0ef,
        64'h84aaa83f_e0ef892a,
        64'ha89fe0ef_842aa8ff,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7f100e8,
        64'h30238f09_00083703,
        64'he3148e89_07856314,
        64'hd15ff06f_6121863e,
        64'h69e2854e_790274a2,
        64'h70e27442_00c79c63,
        64'h974e00e5_88330037,
        64'h97134781_8d5d9101,
        64'h178265a2_66021502,
        64'h8fc18d45_0109179b,
        64'h0105151b_af5fe0ef,
        64'h84aaafbf_e0ef892a,
        64'hb01fe0ef_842ab07f,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7f100e8,
        64'h30238f29_00083703,
        64'he3148ea9_07856314,
        64'hd8dff06f_6121863e,
        64'h69e2854e_790274a2,
        64'h70e27442_00c79c63,
        64'h974e00e5_88330037,
        64'h97134781_8d5d9101,
        64'h178265a2_66021502,
        64'h8fc18d45_0109179b,
        64'h0105151b_b6dfe0ef,
        64'h84aab73f_e0ef892a,
        64'hb79fe0ef_842ab7ff,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7ad0485,
        64'hab1ff0ef_0007c503,
        64'h97e20039_f7930985,
        64'hac1ff0ef_4521ef81,
        64'h00adb023_00acb023,
        64'h8d419101_14021502,
        64'h01a46433_00a96533,
        64'h010d1d1b_0105151b,
        64'h0344f7b3_bd5fe0ef,
        64'h892abdbf_e0ef8d2a,
        64'hbe1fe0ef_842abe7f,
        64'he0efe47f_f06f6165,
        64'h7ae28556_7b4264e6,
        64'h85da8626_6da26d42,
        64'h6ce27c02_7ba26a06,
        64'h69a66946_70a67406,
        64'h8a4fd0ef_06450513,
        64'h00003517_03749b63,
        64'h00fb0cb3_00fa8db3,
        64'h00349793_36cc0c13,
        64'h00003c17_9c4a0a13,
        64'h4981b53f_f0ef4481,
        64'h8bb28b2e_e46ee86a,
        64'hec66e8ca_f0a2f486,
        64'hf062f45e_f85ae4ce,
        64'heca60200_05138aaa,
        64'h6a05fc56_e0d27159,
        64'hb75107a1_05858082,
        64'h61616ba2_6b426ae2,
        64'h7a0279a2_794274e2,
        64'h640660a6_557d91af,
        64'hd0ef0925_05130000,
        64'h3517926f_d0ef0665,
        64'h05130000_3517058e,
        64'h02d60b63_fff7c693,
        64'hc31986be_8b056390,
        64'h00858733_bf6d07a1,
        64'h07056394_e390fff7,
        64'hc613c299_863e8a85,
        64'h008706b3_a0a94501,
        64'h964fd0ef_0fc50513,
        64'h00003517_fd4417e3,
        64'h04050325_99634581,
        64'h87a697ef_d0ef855a,
        64'h85de986f_d0ef854e,
        64'h03271863_470187a6,
        64'h994fd0ef_855685de,
        64'h00040b9b_9a0fd0ef,
        64'h854e4a41_0d4b0b13,
        64'h00003b17_0cca8a93,
        64'h00003a97_0c498993,
        64'h00003997_9c0fd0ef,
        64'h4401892e_e45ee486,
        64'he85aec56_f052f44e,
        64'hf84ae0a2_0d450513,
        64'h00003517_84aafc26,
        64'h715dbf5d_0785a001,
        64'h9ecfd0ef_0d450513,
        64'h00003517_85a28626,
        64'h9fcfd0ef_0bc50513,
        64'h00003517_6090600c,
        64'h02e80363_60980004,
        64'h38038082_61054501,
        64'h64a26442_60e200c7,
        64'h986300d5_043300d5,
        64'h84b30037_96934781,
        64'he426e822_ec061101,
        64'hbbbff06f_80824501,
        64'h80824501_80828082,
        64'h80828082_45098082,
        64'h45098082_4509bff9,
        64'h26052004_04136622,
        64'hdfffc0ef_e4328522,
        64'h85b28082_61454501,
        64'h64e27402_70a20096,
        64'h186300c6_84bb842e,
        64'hf406ec26_f0227179,
        64'h80824505_80824505,
        64'h80824505_80820141,
        64'h8d7d6402_60a29522,
        64'h408007b3_f57ff0ef,
        64'he406952e_842ae022,
        64'h1141a001_cbbff0ef,
        64'h4505abef_d0efe406,
        64'h14850513_00003517,
        64'h85aa862e_86b28736,
        64'h11418082_02f55533,
        64'h47a9b000_25738082,
        64'h45018082_45018082,
        64'h01414501_60a2eadf,
        64'hc0ef2000_0537afaf,
        64'hd0efe406_15c50513,
        64'h00003517_11418082,
        64'h80826105_644260e2,
        64'h8522936f_f0ef4581,
        64'h6622c509_842afd1f,
        64'hf0efe432_8532ec06,
        64'he8221101_02b50633,
        64'h8082953e_055e10d0,
        64'h0513e308_95360017,
        64'h86930075_6513157d,
        64'h631cc227_07130000,
        64'h47178082_45018082,
        64'h24050513_000f4537,
        64'ha001d69f_f0efe406,
        64'h25011141_90020000,
        64'h0023ee1f_f0ef8522,
        64'hb7811c25_05130000,
        64'h3517c511_2501c87f,
        64'ha0ef4501_e3c58593,
        64'h00003597_4605bfb9,
        64'h1c850513_00003517,
        64'hc5112501_b72fb0ef,
        64'ha5050513_00004517,
        64'hbb4fd06f_014106e5,
        64'h05130000_351760a2,
        64'h64024080_05b3cf81,
        64'h439ccae7_87930000,
        64'h47970005_4863842a,
        64'h90ef90ef_ca07ae23,
        64'h00004797_cc07a423,
        64'h00004797_e9850513,
        64'h00000517_bf8fd0ef,
        64'h09850513_00003517,
        64'hb7e121a5_05130000,
        64'h3517c511_2501d69f,
        64'ha0efaba5_05130000,
        64'h45172225_85930000,
        64'h35974605_c28fd0ef,
        64'h21050513_00003517,
        64'hc34fd06f_014160a2,
        64'h64022025_05130000,
        64'h3517c911_2501d47f,
        64'ha0efe022_e406d365,
        64'h05130000_4517f065,
        64'h85930000_35974605,
        64'h11418302_0141bce5,
        64'h85930000_259760a2,
        64'h64028322_f1402573,
        64'h0ff0000f_0000100f,
        64'hc84fd0ef_e40621e5,
        64'h05130000_3517842a,
        64'h85aae022_1141bf95,
        64'hd687ac23_00004797,
        64'h9c25bf5d_2f4010ef,
        64'h854ede7f_f0ef0009,
        64'h4503993e_00397913,
        64'h24878793_00003797,
        64'h0009099b_00c4591b,
        64'he05ff0ef_4521b775,
        64'hdaf72a23_00004717,
        64'h4785cdef_d0ef24e5,
        64'h05130000_351785a6,
        64'h04967563_4632dca7,
        64'ha9230000_4797c50d,
        64'h2501fe3f_a0efba65,
        64'h05130000_451785ca,
        64'h86260074_def72623,
        64'h00004717_57fd8082,
        64'h612169e2_790274a2,
        64'h744270e2_e0a7a423,
        64'h00004797_c10d2501,
        64'hf08fb0ef_bdc50513,
        64'h00004517_02b78563,
        64'h84b2842e_892aec4e,
        64'hfc06f04a_f426f822,
        64'h7139439c_e3478793,
        64'h00004797_80826105,
        64'h60e2e9ff_f0ef0091,
        64'h4503ea7f_f0ef0081,
        64'h4503f13f_f0efec06,
        64'h002c1101_80826145,
        64'h694264e2_740270a2,
        64'hfe9410e3_ec9ff0ef,
        64'h00914503_ed1ff0ef,
        64'h34610081_4503f3ff,
        64'hf0ef0ff5_7513002c,
        64'h00895533_54e10380,
        64'h0413892a_f406e84a,
        64'hec26f022_71798082,
        64'h61456942_64e27402,
        64'h70a2fe94_10e3f0bf,
        64'hf0ef0091_4503f13f,
        64'hf0ef3461_00814503,
        64'hf81ff0ef_0ff57513,
        64'h002c0089_553b54e1,
        64'h4461892a_f406e84a,
        64'hec26f022_71798082,
        64'h61056442_60e2f43f,
        64'hf0ef0091_4503f4bf,
        64'hf0ef0081_4503fb7f,
        64'hf0ef0ff4_7513002c,
        64'hf5dff0ef_00914503,
        64'hf65ff0ef_00814503,
        64'hfd1ff0ef_ec068121,
        64'h842a002c_e8221101,
        64'h808200f5_802300e5,
        64'h80a30007_c7830007,
        64'h470397aa_973e8111,
        64'h00f57713_d6c78793,
        64'h00002797_b7f50405,
        64'hfa5ff0ef_80820141,
        64'h640260a2_e5090004,
        64'h4503842a_e406e022,
        64'h11418082_00e78823,
        64'h02000713_00e78423,
        64'hfc700713_00e78623,
        64'h470d0007_822300e7,
        64'h8023476d_00e78623,
        64'hf8000713_00078223,
        64'h100007b7_808200a7,
        64'h0023dfe5_0207f793,
        64'h01474783_10000737,
        64'h80820205_75130147,
        64'hc5031000_07b78082,
        64'h00054503_808200b5,
        64'h00238082_61056902,
        64'h64a26442_60e2f47d,
        64'hfa1ff0ef_41240433,
        64'h854a8926_0084f363,
        64'h89226804_8493842a,
        64'he04aec06_e8220098,
        64'h94b7e426_11018082,
        64'h61056902_64a26442,
        64'h60e2fe85_6ee3f45f,
        64'hf0ef0405_944a0285,
        64'h54332404_0413000f,
        64'h443702a4_85333e20,
        64'h00ef892a_f63ff0ef,
        64'h84aae04a_e426e822,
        64'hec061101_808202a7,
        64'hd5330141_91011502,
        64'h640260a2_02f407b3,
        64'h24078793_000f47b7,
        64'h414000ef_842af95f,
        64'hf0efe022_e4061141,
        64'h80826105_64a28d05,
        64'h02a7d533_644260e2,
        64'h91011502_02f407b3,
        64'h3e800793_440000ef,
        64'h842afc1f_f0ef84aa,
        64'he426e822_ec061101,
        64'h80824501_80820141,
        64'h8d5d9101_17821502,
        64'h60a21007_e78310a7,
        64'ha22310e1_a0232705,
        64'h1001a703_00e57763,
        64'h878e1041_e7035040,
        64'h00efe406_11418082,
        64'hcf1ff06f_c7458593,
        64'h00004597_4611cb81,
        64'he8c7d783_00004797,
        64'h80822401_01132201,
        64'h39032281_34832301,
        64'h34032381_3083f63f,
        64'hf0ef8522_002ce90f,
        64'hf0efe802_c44a0828,
        64'h20400613_85a6e52f,
        64'hf0ef2211_3c230028,
        64'h21800613_45818932,
        64'h84ae842a_23213023,
        64'h22913423_22813823,
        64'hdc010113_ebfff06f,
        64'h614505c1_70a24190,
        64'h7402d8bf_f06f6145,
        64'h70a265a2_74028522,
        64'h875fd0ef_e42e5ae5,
        64'h05130000_3517842a,
        64'h885fd06f_61455d65,
        64'h05130000_351770a2,
        64'h740202f7_0a63478d,
        64'h00d70e63_01e15703,
        64'h00e10f23_0115c703,
        64'h00e10fa3_46890105,
        64'hc703f022_f4067179,
        64'h80826105_690264a2,
        64'h644260e2_d47ff06f,
        64'h61056902_64a260e2,
        64'h64428d7f_d0ef5f65,
        64'h05130000_35170087,
        64'hcf63278d_439cf767,
        64'h87930000_4797f8f7,
        64'h11230000_47172785,
        64'h0007d783_f9078793,
        64'h00004797_240000ef,
        64'h02000513_d19ff0ef,
        64'h4515fa65_d5830000,
        64'h45972560_00ef4535,
        64'he29ff0ef_854adae5,
        64'h85930000_4597daa7,
        64'h9c230000_47974611,
        64'hcf3ff0ef_fd055503,
        64'h00004517_dca79623,
        64'h00004797_d07ff0ef,
        64'h4511da9f_f0ef0044,
        64'h8513ffc4_059b06a7,
        64'h9a632501_0024d783,
        64'hd23ff0ef_00055503,
        64'h00004517_08a79563,
        64'h25010004_d783d39f,
        64'hf0ef84ae_450d892a,
        64'h08c7df63_8432478d,
        64'he04ae426_ec06e822,
        64'h1101b791_02f71823,
        64'h00004717_4785eaff,
        64'hf0ef854e_e3458593,
        64'h00004597_4611e4a7,
        64'h90230000_4797d79f,
        64'hf0ef4501_e4a79623,
        64'h00004797_d87ff0ef,
        64'h06f73823_00004717,
        64'h06f73823_00004717,
        64'h451107e2_08100793,
        64'h9edfd0ef_6ec50513,
        64'h00003517_858a4390,
        64'h08878793_00004797,
        64'hdecff0ef_850a85a2,
        64'hdf4ff0ef_850a7065,
        64'h85930000_359700f7,
        64'h096302f0_07930129,
        64'h4703de0f_f0ef850a,
        64'h4d858593_00003597,
        64'h855ff0ef_850a4581,
        64'h10000613_b7550cf7,
        64'h27230000_47172000,
        64'h07938082_615569b2,
        64'h695264f2_741270b2,
        64'ha5dfd0ef_73450513,
        64'h00003517_00a405b3,
        64'hf1cff0ef_51c50513,
        64'h00003517_842af2af,
        64'hf0ef8522_04a7f263,
        64'h0ff00793_9526f3af,
        64'hf0ef53a5_05130000,
        64'h351784aa_f48ff0ef,
        64'h852212a7_a5230000,
        64'h479704e7_ee631ff0,
        64'h0793fff5_071be93f,
        64'hf0ef9526_0505f6af,
        64'hf0ef8526_00a404b3,
        64'h0505f76f_f0ef892e,
        64'hea4aee26_f6068522,
        64'h89aae64e_01258413,
        64'hf2227169_80824501,
        64'h80820141_640260a2,
        64'h8522547d_00850363,
        64'h874fa0ef_8432e406,
        64'he0221141_66a0006f,
        64'h610564a2_60e26442,
        64'hb0dfd06f_61057c65,
        64'h05130000_351740a0,
        64'h05b364a2_60e26442,
        64'h00055e63_85bf90ef,
        64'hef850513_00000517,
        64'hb35fd0ef_7d450513,
        64'h00003517_b41fd0ef,
        64'h7c850513_00003517,
        64'h862286aa_608ce2df,
        64'hc0ef85a2_6088b5bf,
        64'hd0ef85a2_9c11ec06,
        64'h7d050513_00003517,
        64'h6380e822_60902064,
        64'h84930000_4497e426,
        64'h21878793_00004797,
        64'h11018082_610564a2,
        64'h6442e00c_95a660e2,
        64'h600ca05f_f0efec06,
        64'h600885aa_84ae862e,
        64'he4262424_04130000,
        64'h4417e822_11018082,
        64'h24f73823_00004717,
        64'h24f73823_00004717,
        64'h07e20810_07935020,
        64'h006f0305_05130141,
        64'h60a26402_02a4753b,
        64'h4529fe7f_f0ef357d,
        64'h02b455bb_45a900b7,
        64'hf86347a5_00a04563,
        64'h842ee406_e0221141,
        64'hb7c50505_fd07879b,
        64'h9fb902f6_07bb00b6,
        64'he763fd07_059b2701,
        64'h8082853e_e3190005,
        64'h47034629_46a54781,
        64'ha93ff06f_95be9201,
        64'h16029181_1582639c,
        64'h2c878793_00004797,
        64'h80820141_91411542,
        64'h11418d5d_05220085,
        64'h579bfa5f_f06f4581,
        64'hd7dff06f_01410505,
        64'h45814629_60a26402,
        64'hf77d8b11_00074703,
        64'h973e0005_4703fea4,
        64'h7ae3157d_80820141,
        64'h557d6402_60a2e719,
        64'h8b110007_4703973e,
        64'hfff58513_e3478793,
        64'h00002797_fff5c703,
        64'h00a405b3_951ff0ef,
        64'he589842a_e406e022,
        64'h1141bfd5_0789bff1,
        64'h052a052a_b7e9e01c,
        64'h078d00e6_98630420,
        64'h07130027_c683fce6,
        64'h9fe3052a_06900713,
        64'h0017c683_fed716e3,
        64'h06b00693_02d70763,
        64'h04d00693_80820141,
        64'h640260a2_02d70e63,
        64'h04700693_00e6ea63,
        64'h02d70463_0007c703,
        64'h04b00693_601cf87f,
        64'hf0ef842e_e406e022,
        64'h1141b7e1_e008b7cd,
        64'hfc97879b_0ff7f793,
        64'hfe07079b_c6098a09,
        64'hb7d196be_050502d5,
        64'h86b3feb7_f4e3fd07,
        64'h879b0008_8b630046,
        64'h78938082_61058536,
        64'h644260e2_ec050008,
        64'h98630446_78930006,
        64'h460300f8_06330007,
        64'h079b0005_4703f0e8,
        64'h08130000_28174681,
        64'h00c16583_e0dff0ef,
        64'hc632ec06_006c842e,
        64'he8221101_bfd50789,
        64'hbff1052a_052ab7e9,
        64'he01c078d_00e69863,
        64'h04200713_0027c683,
        64'hfce69fe3_052a0690,
        64'h07130017_c683fed7,
        64'h16e306b0_069302d7,
        64'h076304d0_06938082,
        64'h01416402_60a202d7,
        64'h0e630470_069300e6,
        64'hea6302d7_04630007,
        64'hc70304b0_0693601c,
        64'hf0dff0ef_842ee406,
        64'he0221141_80820141,
        64'h40a00533_60a2f23f,
        64'hf0efe406_05051141,
        64'hf2dff06f_00e68463,
        64'h02d00713_00054683,
        64'hb7e94501_e088fcf7,
        64'h18e347a9_fd279be3,
        64'h07858f81_cb010007,
        64'hc703fe87_82e367e2,
        64'hf5dff0ef_8522082c,
        64'h892a862e_80826121,
        64'h790274a2_744270e2,
        64'h5529e901_65a2b03f,
        64'hf0ef84b2_842ae42e,
        64'h00063023_f04afc06,
        64'hf426f822_7139b7e1,
        64'he008b7cd_fc97879b,
        64'h0ff7f793_fe07079b,
        64'hc6098a09_b7d196be,
        64'h050502d5_86b3feb7,
        64'hf4e3fd07_879b0008,
        64'h8b630046_78938082,
        64'h61058536_644260e2,
        64'hec050008_98630446,
        64'h78930006_460300f8,
        64'h06330007_079b0005,
        64'h47030628_08130000,
        64'h28174681_00c16583,
        64'hf61ff0ef_c632ec06,
        64'h006c842e_e8221101,
        64'h8082fae7_8fe34741,
        64'hbfed47a9_8082c19c,
        64'h47a1a809_050900e7,
        64'h9c630780_07130ff7,
        64'hf7930207_879bc709,
        64'h8b050007_4703973e,
        64'h0b070713_00002717,
        64'h00154783_02f71f63,
        64'h03000793_00054703,
        64'hc19c47c1_cf950447,
        64'hf7930007_c78397ba,
        64'h00254703_04d71763,
        64'h07800693_0ff77713,
        64'h0207071b_c6898a85,
        64'h0006c683_00e786b3,
        64'h0f878793_00002797,
        64'h00154703_06f71e63,
        64'h03000793_00054703,
        64'he7c9419c_b7f1377d,
        64'h87aabfa5_fef51be3,
        64'h0785f8b7_12e30007,
        64'hc70300d8_0a630087,
        64'h85130007_b803bfcd,
        64'h367d0785_f8b71fe3,
        64'h0007c703_d24d8a1d,
        64'heb1187aa_27018edd,
        64'h00365713_02079693,
        64'h8fd90107_179300b7,
        64'he7330085_97938e19,
        64'h953a9301_1702fed8,
        64'h19e30007_869b0785,
        64'hfcb69de3_0007c683,
        64'h87aa00a7_083b9f1d,
        64'h4721c39d_00757793,
        64'hb7f5367d_0785feb7,
        64'h1ce30007_c7038082,
        64'h853e4781_e60187aa,
        64'h260100c7_ef630ff5,
        64'hf59347c1_b7ed853e,
        64'hfeb70be3_00150793,
        64'h00054703_80824501,
        64'h00c51463_0ff5f593,
        64'h962abfe1_0405d17d,
        64'hf83ff0ef_852285ca,
        64'h86268082_614569a2,
        64'h694264e2_740270a2,
        64'h85224401_0097db63,
        64'h408987bb_008509bb,
        64'hd0dff0ef_8522c899,
        64'h0005049b_d19ff0ef,
        64'h892ee44e_f406e84a,
        64'hec26852e_842af022,
        64'h7179bfc5_0505feb7,
        64'h8de30005_47838082,
        64'h00c51363_962a8082,
        64'h853ed3f5_9f950705,
        64'h0006c683_0007c783,
        64'h00e586b3_00e507b3,
        64'ha8214781_00e61463,
        64'h4701b7e5_00b70023,
        64'h97220005_c58300e6,
        64'h85b300f8_0733fef6,
        64'h05e317fd_4781fff6,
        64'h461386ae_88328082,
        64'h01416402_60a28522,
        64'hf53ff0ef_00a5e963,
        64'h842ae406_e0221141,
        64'h80826145_64e26942,
        64'h85267402_70a20004,
        64'h0023f75f_f0ef944a,
        64'h864a8522_fff60913,
        64'h00c56463_6582892a,
        64'hce1184aa_6622dd3f,
        64'hf0efe02e_e84af406,
        64'he432ec26_852e842a,
        64'hf0227179_b7e50106,
        64'h80230785_00f706b3,
        64'h0006c803_00f586b3,
        64'h808200f6_13634781,
        64'h00f50733_963a95be,
        64'h078e02e7_87335761,
        64'h00365793_fed765e3,
        64'h40f606b3_0106b023,
        64'h07a100f5_06b30006,
        64'hb80300f5_86b3a811,
        64'h471d4781_eb9d872a,
        64'h8b9d00b5_67b304b5,
        64'h0463b7f5_feb78fa3,
        64'h0785bfe9_fee7bc23,
        64'h07a18082_00c79763,
        64'h963e963a_97aa078e,
        64'h02e78733_57610036,
        64'h57930106_ee6340f8,
        64'h8833469d_00c508b3,
        64'h87aaffed_8f5537fd,
        64'h07220ff5_f69347a1,
        64'heb0587aa_00757713,
        64'h80824501_b7e50789,
        64'h00d780a3_00e78023,
        64'h8082e311_0017c703,
        64'hce810007_c68387aa,
        64'hcf990005_4783c11d,
        64'h80826105_64a28526,
        64'h644260e2_e0080505,
        64'h00050023_c501f73f,
        64'hf0ef8526_842ac891,
        64'he822ec06_6104e426,
        64'h1101bfd9_6aa7ba23,
        64'h00004797_05050005,
        64'h0023c781_00054783,
        64'hc519f9ff_f0ef8522,
        64'h85a68082_610564a2,
        64'h644260e2_85224401,
        64'h6e07b023_00004797,
        64'hef810004_4783942a,
        64'hfa1ff0ef_85a68522,
        64'hcc116380_6fc78793,
        64'h00004797_e519842a,
        64'h84aeec06_e426e822,
        64'h1101bfd5_87aeb7e5,
        64'h0505fafd_0007c683,
        64'h0785fee6_8fe38082,
        64'h4501eb19_00054703,
        64'hb7c50785_8082853e,
        64'hfa7d0007_46030705,
        64'h00d60863_a021872e,
        64'hca890007_468300f5,
        64'h07334781_bfd5872e,
        64'hb7d50785_fa7d0007,
        64'h46030705_fed60ee3,
        64'h8082853e_ea990007,
        64'h468300f5_07334781,
        64'hb7fd0785_808240a7,
        64'h8533e701_0007c703,
        64'h00b78563_87aa95aa,
        64'h80826105_644260e2,
        64'h4501fe85_7be3157d,
        64'h00b78663_00054783,
        64'h0ff5f593_952265a2,
        64'hfe5ff0ef_ec06842a,
        64'he42ee822_1101bfcd,
        64'h07858082_40a78533,
        64'he7010007_c70387aa,
        64'hbfcd0505_dffd8082,
        64'h00b79363_00054783,
        64'h0ff5f593_80824501,
        64'hbfcd0505_c3998082,
        64'h00b79363_00054783,
        64'h0ff5f593_8082853e,
        64'hfee10705_e3994187,
        64'hd79b0187_979b40f6,
        64'h87bb0007_c78300e5,
        64'h87b30007_c68300e5,
        64'h07b3a015_478100e6,
        64'h14634701_8082853e,
        64'hf37d0505_e3994187,
        64'hd79b0187_979b40f7,
        64'h07bbfff5_c7830005,
        64'h47030585_80820007,
        64'h8023fec7_99e3d375,
        64'hfee78fa3_0785fff5,
        64'hc7030585_963efb7d,
        64'h00178693_0007c703,
        64'h87b68082_e21987aa,
        64'hb7d587b6_8082fb75,
        64'hfee78fa3_0785fff5,
        64'hc7030585_eb090017,
        64'h86930007_c70387aa,
        64'h8082f76d_00e68023,
        64'h078500f5_06b30007,
        64'h470300f5_873300c7,
        64'h8c634781_8082fb75,
        64'hfee78fa3_0785fff5,
        64'hc7030585_87aa8082,
        64'h01416402_60a28d41,
        64'h15029001_fd1ff0ef,
        64'h14020005_041bfdbf,
        64'hf0efe022_e4061141,
        64'h80820141_25016402,
        64'h60a28d41_0105151b,
        64'hfe9ff0ef_842afeff,
        64'hf0efe022_e4061141,
        64'hfc3ff06f_8fc50513,
        64'h00005517_80822501,
        64'h8d5d00f7_17bb40f0,
        64'h07bb00f7_553b93ed,
        64'h836d8f3d_0127d713,
        64'he1189736_00176713,
        64'h02d786b3_65186294,
        64'h611c6d26_86930000,
        64'h46971c60_106f8082,
        64'h61056902_64a26442,
        64'h60e28522_e99ff0ef,
        64'h10f40023_0247c783,
        64'h85220ea4_2e23681c,
        64'h18f43423_2b878793,
        64'h00001797_18f43023,
        64'h2c878793_00001797,
        64'h16f43c23_8fa78793,
        64'hfffff797_e65ff0ef,
        64'h04052823_03253023,
        64'he90410f5_02a34785,
        64'h0ef52c23_4799c57c,
        64'h57fdcd21_842a20a0,
        64'h10ef4505_1c000593,
        64'h84aa892e_c7ad639c,
        64'hc7bd651c_cbad511c,
        64'hcbbd4d5c_cfad4401,
        64'h4d1cc141_4401e04a,
        64'he426ec06_e8221101,
        64'hb7716000_334010ef,
        64'h7b850513_00003517,
        64'h01a98863_d80fe0ef,
        64'h856685e2_00978e63,
        64'h601cd8ef_e0ef855e,
        64'h85ca0009_0663d9af,
        64'he0ef638c_855a0fc4,
        64'h2603681c_89560007,
        64'hc3638952_4c1cc791,
        64'h4901541c_db8fe06f,
        64'h612539a5_05130000,
        64'h45176d02_6ca26c42,
        64'h6be27b02_7aa27a42,
        64'h79e26906_64a660e6,
        64'h64460294_15634d29,
        64'h830c8c93_00004c97,
        64'h00050c1b_24cb8b93,
        64'h00004b97_24cb0b13,
        64'h00004b17_24ca8a93,
        64'h00004a97_24ca0a13,
        64'h00004a17_89aae0ca,
        64'hec86e06a_e466e862,
        64'hec5ef05a_f456f852,
        64'hfc4e6080_e8a2a864,
        64'h84930000_5497e4a6,
        64'h711d8082_e308e518,
        64'he11ce788_6798a9e7,
        64'h87930000_5797e508,
        64'h80828e07_a9230000,
        64'h5797e79c_e39cab67,
        64'h87930000_5797b7d5,
        64'h6000a8cf_f0ef8522,
        64'hc78119a4_47838082,
        64'h610564a2_644260e2,
        64'h00941763_84beec06,
        64'he4266380_e822ae67,
        64'h87930000_57971101,
        64'h80824388_93c78793,
        64'h00005797_80820f85,
        64'h05138082_c3980015,
        64'h071b4388_95478793,
        64'h00005797_bfd55535,
        64'h80826105_64a26442,
        64'h60e2e080_0f840413,
        64'he501ce0f_f0ef842a,
        64'hcd09f7df_f0ef84ae,
        64'he822ec06_e4261101,
        64'hbfcdf840_0513bfe5,
        64'h45018082_610560e2,
        64'h5535e97f_e06f6105,
        64'h60e200f7_0c630ff0,
        64'h07930815_470302b7,
        64'h006365a2_10354703,
        64'hc105fbdf_f0efe42e,
        64'hec061101_41488082,
        64'h853ebfd1_87b600a6,
        64'h04630fc7_a6038082,
        64'h0141853e_478160a2,
        64'hf3cfe0ef_e4063665,
        64'h05130000_451785aa,
        64'h114102e7_90636394,
        64'h631cbb27_07130000,
        64'h57178082_45018082,
        64'h01414501_640260a2,
        64'h0dc000ef_13e000ef,
        64'h02c00513_fc5ff0ef,
        64'h85220005_5563ac0f,
        64'he0ef8522_12a000ef,
        64'hbef72223_00005717,
        64'h842ae406_e0224785,
        64'h1141ef9d_439cbfa7,
        64'h87930000_57978082,
        64'h18b50d23_8082557d,
        64'h8082557d_80824501,
        64'hc56c8702_972a4318,
        64'h972a8379_d3c50513,
        64'h00003517_1702ef05,
        64'h6863450d_0007081b,
        64'h377d8b3d_01a6571b,
        64'hf0e51c63_40000737,
        64'h06bba423_06dba223,
        64'h06fba023_04cbae23,
        64'h018ba503_45e646d6,
        64'h47c64636_e8051763,
        64'h842a90ff_e0efc4be,
        64'h855e0107_979b008c,
        64'h460107cb_d783c2be,
        64'h479d04f1_102347a5,
        64'h06fb9e23_04e15783,
        64'h0007d663_018ba783,
        64'hec051163_842a943f,
        64'he0efc2be_47d5855e,
        64'hc4be0107_979b008c,
        64'h460107cb_d78304f1,
        64'h1023478d_6ce000ef,
        64'h06cb8513_00ec4641,
        64'hef2ff06f_fa100413,
        64'hbf6d1187_25839752,
        64'h83790207_9713fcfc,
        64'h65e34581_bfa1d171,
        64'hd13fe0ef_855e4585,
        64'h0b700613_0ff6f693,
        64'hbb35f53d_9d9fe0ef,
        64'h855ec9af_f0ef855e,
        64'h460118fb_ae2308bb,
        64'ha2230017_b79317ed,
        64'h088ba583_ef8d1afb,
        64'ha823409c_e79d0046,
        64'hf7930089_2683f14d,
        64'hfeffe0ef_855e408c,
        64'h913fe0ef_855e02eb,
        64'haa230017_b71341b7,
        64'h87b301a7_86634711,
        64'h00d78963_47214000,
        64'h06b70009_2783bfa5,
        64'hfb9910e3_0931941f,
        64'he0ef855e_035baa23,
        64'h08fba223_180bae23,
        64'h1a0ba823_088ba783,
        64'hdabfe0ef_855e4585,
        64'h0b700613_4681c90d,
        64'hdbbfe0ef_855e0fb6,
        64'hf6934585_0b700613,
        64'h00894683_c3a12781,
        64'h8ff900f9_f7b30009,
        64'h270340dc_04f71963,
        64'h0017b793_17ed0049,
        64'h4703409c_10000db7,
        64'h20000d37_fac90913,
        64'h00003917_bd2197bf,
        64'he0ef4325_05130000,
        64'h4517ff64_98e304a1,
        64'heb992781_00f9f7b3,
        64'h00fa97bb_409c012c,
        64'h8c930000_3c974c2d,
        64'hfe0b0b13_00003b17,
        64'h4a85fca4_84930000,
        64'h3497daaf_f0ef2981,
        64'h855e00f9_f9b34601,
        64'h088ba583_044ba783,
        64'h040ba983_e6f769e3,
        64'h400407b7_04fba023,
        64'h00c7e793_040ba783,
        64'hd7dd8b85_04dba023,
        64'h0106e693_040ba683,
        64'h04dba023_0216869b,
        64'hc58900c7_f593cd91,
        64'h0027f593_1abba423,
        64'h03f7f593_0c464783,
        64'h04fba023_0016879b,
        64'h700006b7_b1294f65,
        64'h05130000_4517e611,
        64'hb5f1e225_ecf769e3,
        64'h400407b7_00f77863,
        64'h1a0bb603_400407b7,
        64'h04fba023_27851000,
        64'h07b7b0cd_02fba423,
        64'h478500d0_10ef8526,
        64'ha39fe0ef_8a3d8abd,
        64'h0146561b_0106569b,
        64'h06248513_58458593,
        64'h00004597_074ba603,
        64'ha59fe0ef_04d48513,
        64'h58858593_00004597,
        64'h0186d69b_0ff77713,
        64'h0ff7f793_0ff6f813,
        64'h0106d71b_0086d79b,
        64'h06cbc603_077bc883,
        64'h070ba683_a8dfe0ef,
        64'hfef53623_02450513,
        64'h5a858593_00004597,
        64'h84aa06fb_c603074b,
        64'hd68307ab_d70302c7,
        64'hd7b3ed10_92010a8b,
        64'hb783d11c_9fb90712,
        64'h00e03733_8f750207,
        64'h161376c1_9fb5068e,
        64'h00d036b3_8ef9f006,
        64'h8693ff01_06b79fb5,
        64'h068a00d0_36b38ef9,
        64'h0f068693_f0f0f6b7,
        64'h9fb500f0_37b30686,
        64'h00d036b3_27818ef9,
        64'h8ff9ccc6_8693aaa7,
        64'h8793cccc_d6b7aaaa,
        64'hb7b708cb_a7030005,
        64'h06230005_15234a00,
        64'h00ef855e_08fba823,
        64'h08fba623_20000793,
        64'hc79919cb_a7831afb,
        64'haa231b0b_a7830adb,
        64'ha2230afb_a02302d6,
        64'h06bb02f7_57bb8a8d,
        64'h0106d69b_02e6073b,
        64'h3e800613_c30503f7,
        64'h77130126_d71bc78d,
        64'h27818fd1_8ff90186,
        64'hd61b17fd_67c100cd,
        64'ha68308fb_ae230087,
        64'h171b1487_a78397b6,
        64'h078a1326_86930000,
        64'h369704d6_1c638003,
        64'h06b7018b_a60300f6,
        64'hf8638bbd_00c7579b,
        64'h46a5008d_a703fda5,
        64'h9ee3fefd_2e238fd9,
        64'h8ff58f51_0087d79b,
        64'h8e690087_961b8f51,
        64'h0187971b_0187d61b,
        64'h0d11000d_2783f006,
        64'h869300ff_0537040d,
        64'h059366c1_bf911187,
        64'h25839752_83790207,
        64'h9713f6f7_62e34581,
        64'h472db575_def98be3,
        64'h10bc0991_81dff0ef,
        64'h855e8405_85934601,
        64'h180bae23_096ba223,
        64'h1afba823_017d85b7,
        64'h4785f3f5_37fd6702,
        64'h67a2c521_d51fe0ef,
        64'he03ac93a_e556e16a,
        64'he43e855e_110c0110,
        64'h04000713_4791d502,
        64'h8dead33a_0af11023,
        64'hfe0c7d13_47b56702,
        64'hed05d7ff_e0efd53e,
        64'he03ad33a_855e110c,
        64'h0107979b_46014755,
        64'h07cbd783_0af11023,
        64'h03700793_895ff0ef,
        64'h855e4601_18fbae23,
        64'h08bba223_0017b793,
        64'h17ed088b_a583efd9,
        64'h1afba823_409c09b7,
        64'h90638bbd_010cc783,
        64'he541dcff_e0efc93e,
        64'he556e166_855e110c,
        64'h04000793_0110d53e,
        64'h00fde7b3_17c12d81,
        64'h810007b7_d33e47d5,
        64'h0af11023_47994d85,
        64'h0ae79d63_470d00e7,
        64'h86634705_409cd41f,
        64'he0ef855e_02fbaa23,
        64'h001d3793_40fd0d33,
        64'h100007b7_00ed0863,
        64'h47912000_073700ed,
        64'h0d6347a1_40000737,
        64'h0e051963_8daa8bff,
        64'hf0ef855e_0015b593,
        64'h40bd05b3_100005b7,
        64'h00fd0863_45912000,
        64'h07b700fd_0d6345a1,
        64'h400007b7_12078e63,
        64'h278101a7_f7b300f9,
        64'h77b30009_ad0340dc,
        64'h840b0b1b_06010993,
        64'h017d8b37_bf0104fb,
        64'ha0230087_e793040b,
        64'ha783f207_50e302e7,
        64'h97138fd5_8ff90087,
        64'hd79b0087_969bf007,
        64'h07136741_44dcfbe1,
        64'h8b8583a5_4cdce605,
        64'h1de3eb7f_e0efdc3e,
        64'hf84af426_c556855e,
        64'h010c0400_07931030,
        64'hc33e47d5_08f11023,
        64'h47990209_886339fd,
        64'h09053ac5_49959881,
        64'h19020100_0ab70ff1,
        64'h04934905_bfa98003,
        64'h0737b785_80020737,
        64'h00074563_03079713,
        64'hb7bda007_071b8001,
        64'h1737b949_df400413,
        64'he15fe0ef_8cc50513,
        64'h00005517_fef493e3,
        64'h44078793_00003797,
        64'h04a1ebc5_278100f9,
        64'h77b300e7_97bb4785,
        64'h40980a85_83f97913,
        64'h02079a93_478500f9,
        64'h7933fe0c_7c9345e4,
        64'h84930000_3497044b,
        64'ha783f0be_0ff10c13,
        64'h040ba903_639c06e7,
        64'h87930000_579708f7,
        64'h13638001_07b7018b,
        64'ha70304fb_a0238fd9,
        64'h20000737_040ba783,
        64'h00075963_02d79713,
        64'h00ebac23_80010737,
        64'h08d70e63_4689c701,
        64'h09270d63_8b3d0187,
        64'hd71b04eb_ac238f55,
        64'h8f718ecd_0087571b,
        64'h8de90087_159b8ecd,
        64'h0187169b_0187559b,
        64'h40d804fb_aa232781,
        64'h8fd58ef1_f0070613,
        64'h8fd16741_0087569b,
        64'h8e698fd5_0087161b,
        64'h0187179b_0187569b,
        64'h00ff0537_4098bd79,
        64'h8a9d9381_00f6d69b,
        64'h17828fd9_01e6d71b,
        64'h8ff90027_979b1771,
        64'h6705b545_08bba823,
        64'h00b515bb_89bd0165,
        64'hd59bbd91_40040737,
        64'hbda94003_0737bd89,
        64'h40020737_bb75842a,
        64'hfe0996e3_39fdc529,
        64'h844ff0ef_d05aec56,
        64'he826855e_108c0810,
        64'h4b210a85_4991d482,
        64'h06f11023_98810209,
        64'h1a930330_07930bf1,
        64'h04934905_d2caed05,
        64'h874ff0ef_d4bed2ca,
        64'h855e0107_979b108c,
        64'h460107cb_d78306f1,
        64'h10230370_079304fb,
        64'ha0232789_100007b7,
        64'h54075963_018ba703,
        64'he20515e3_842aff3f,
        64'he0ef855e_00b54583,
        64'h113000ef_855ee405,
        64'h10e3842a_c94ff0ef,
        64'h855e08fb_80a357fd,
        64'h08fbaa23_4785e405,
        64'h1ce3842a_8d8ff0ef,
        64'hc4bec2ca_855e008c,
        64'h0107979b_46014955,
        64'h07cbd783_04f11023,
        64'h479d8f6f_f0efc282,
        64'hc4be04e1_1023855e,
        64'h008c4601_0107979b,
        64'h471100e7_8e63577d,
        64'h04cba783_c21508fb,
        64'ha82300e7_f4632000,
        64'h0793090b_a70308fb,
        64'ha6230107_d4632000,
        64'h07930afb_b8230e0b,
        64'hb0230c0b_bc230c0b,
        64'hb8230c0b_b4230c0b,
        64'hb0230a0b_bc230307,
        64'h87b300d7_97b32689,
        64'h078546a1_8fd90106,
        64'hd79b8f7d_003f0737,
        64'h0107979b_14070f63,
        64'h02cba703_090ba823,
        64'h1408dd63_090ba623,
        64'h00e5183b_8b3d0107,
        64'hd71b08eb_a22308eb,
        64'ha42304cb_a823180b,
        64'hae231a0b_a8238a05,
        64'h00c7d61b_02c7073b,
        64'h018ba883_45050f87,
        64'h47031086_26039652,
        64'h9752060a_8b3d646a,
        64'h0a130000_3a178a1d,
        64'h0036571b_00ebac23,
        64'h4007071b_40010737,
        64'ha0292007_071b4001,
        64'h0737bf05_06fb9e23,
        64'h478502fb_a6238b85,
        64'h41e7d79b_048ba783,
        64'h00fbac23_400007b7,
        64'hbfe91f10_10ef0640,
        64'h051308a9_6fe31630,
        64'h10ef8526_0007cc63,
        64'h048ba783_f155842a,
        64'hb1eff0ef_855e4585,
        64'h3e800913_90810205,
        64'h14931870_10ef4501,
        64'hafeff0ef_855e0407,
        64'hc163180b_8c23048b,
        64'ha7838082_615d6db6,
        64'h6d566cf6_7c167bb6,
        64'h7b567af6_6a1a69ba,
        64'h695a64fa_741a70ba,
        64'h8522d55d_842ad99f,
        64'hf0ef855e_a031020b,
        64'ha423f4fd_34fd1005,
        64'h0de3842a_a88ff0ef,
        64'h855e008c_46014495,
        64'hcf818b85_1b8ba783,
        64'h12050ae3_842aaa2f,
        64'hf0efc482_c2be855e,
        64'h008c479d_460104f1,
        64'h10234789_e7b5180b,
        64'h8ca3198b_c783c7b1,
        64'h199bc783_219010ef,
        64'h45018baa_e3b54401,
        64'he6eeeaea_eee6f2e2,
        64'hf6defada_fed6e352,
        64'he74eeb4a_ef26f706,
        64'hf3227161_551cb585,
        64'h84aab595_fa100493,
        64'h9fcff0ef_c8450513,
        64'h00005517_d965c04f,
        64'hf0ef8522_4585bfd1,
        64'h18f40c23_47850007,
        64'hd663443c_ed09c1cf,
        64'hf0ef8522_4581becf,
        64'hf0ef8522_02f51f63,
        64'hf9200793_b55d18f4,
        64'h0ca34785_06041e23,
        64'hd45c8b85_41e7d79b,
        64'hc43ccc18_80010737,
        64'h00e68563_80020737,
        64'h4c14bf45_34b010ef,
        64'h3e800513_06090863,
        64'h397d0007_ca6347b2,
        64'hed1db76f_f0ef8522,
        64'h858a4601_c43e0197,
        64'he7b30187_1563c43e,
        64'h0177f7b3_c25a4bdc,
        64'h01511023_4c18681c,
        64'he13db9ef_f0efc402,
        64'hc2520131_10238522,
        64'h858a4601_40000cb7,
        64'h80020c37_00ff8bb7,
        64'h4b050290_0a934a55,
        64'h03700993_3e900913,
        64'hcc1c8002_07b700f7,
        64'h15630aa0_079300c1,
        64'h4703e911_be0ff0ef,
        64'hc23ec43a_8522858a,
        64'h460147d5_0aa00713,
        64'he3991aa0_07138ff9,
        64'h4bdc00ff_8737681c,
        64'h00f11023_47a10005,
        64'h05a346d0_00ef8522,
        64'hf14984aa_cdaff0ef,
        64'h8522f13f_f0ef8522,
        64'h45814601_b5eff0ef,
        64'h8522d85c_478508f4,
        64'h22231a04_28231804,
        64'h2e230884_2783f945,
        64'h84aa9782_6b9c679c,
        64'h8522681c_43b010ef,
        64'h7d000513_b8eff0ef,
        64'h85220204_2c2302f4,
        64'h08234785_1af42c23,
        64'h478df93f_f0eff3e5,
        64'h4481541c_80826109,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e674a6,
        64'h79068526_744670e6,
        64'hf8500493_b98ff0ef,
        64'he0850513_00005517,
        64'h02042423_eb8d6b9c,
        64'h679c681c_c509f07f,
        64'hf0ef842a_c17c8fd9,
        64'hf466f862_fc5ee0da,
        64'he4d6e8d2_eccef0ca,
        64'hf4a6fc86_f8a2070d,
        64'h4b9c7119_10000737,
        64'h691c8082_8082c18f,
        64'hf06f02c5_0823dd0c,
        64'h0007859b_87ba00d5,
        64'hf3630007_069b0007,
        64'h859b4f18_87ae00d5,
        64'hf3630007_869b4f5c,
        64'h6918e215_b7cdc402,
        64'hfef414e3_47858082,
        64'h61217902_74a27442,
        64'h70e2d26f_f0ef8526,
        64'h858a4601_c43e4789,
        64'h00f41f63_4791c24a,
        64'h00f11023_4799ed19,
        64'hd44ff0ef_c43ec24a,
        64'h8526858a_46010107,
        64'h979b4955_842e07c4,
        64'hd78300f1_10230370,
        64'h079304f5_92635529,
        64'h478500f5_866384aa,
        64'h4791f04a_f822fc06,
        64'hf4267139_80820141,
        64'h640260a2_45058302,
        64'h014160a2_64028522,
        64'h00030763_0187b303,
        64'h679c681c_00055e63,
        64'hffdfe0ef_842ae406,
        64'he0221141_b325842a,
        64'hb335dd79_842a941f,
        64'hf0ef8526_45850a70,
        64'h061386ca_b381842a,
        64'h953ff0ef_85264585,
        64'h09b00613_46850127,
        64'h9b630a79_c783d4fb,
        64'h0ee34785_ed19971f,
        64'hf0ef8526_458509c0,
        64'h061386de_fdba18e3,
        64'h0c110ffa_7a132a0d,
        64'hffac90e3_0ffafa93,
        64'h2ca12a85_e139999f,
        64'hf0ef8526_0ff6f693,
        64'h0196d6bb_45858656,
        64'h000c2683_4c818ad2,
        64'h09b00d93_4d6108f0,
        64'h0a13ff9a_10e32a05,
        64'he92d9c5f_f0ef8526,
        64'h45850ff6_76130ff6,
        64'hf693f8ca_061b00da,
        64'hd6bb003a_169b4c8d,
        64'hfdbd1fe3_2d05e945,
        64'h8a2a9edf_f0ef8526,
        64'h45850ff6_76130ff6,
        64'hf693f88d_061b00dc,
        64'hd6bb003d_169b4d91,
        64'h4d0108f4_aa2300a7,
        64'h979b0e09_c7830af9,
        64'h87a34785_e579a21f,
        64'hf0ef8526_45850af0,
        64'h06134685_e3958b85,
        64'h0af9c783_e20b05e3,
        64'hb535547d_db8ff0ef,
        64'h00850513_00005517,
        64'hcb898b85_09b9c783,
        64'hbfd100f9_7933fff7,
        64'hc793b5a9_39c020ef,
        64'hfd850513_00005517,
        64'hef898b85_0a69c783,
        64'h02d90263_fcb614e3,
        64'h87b20ff9_79130127,
        64'he933c70d_4189591b,
        64'h4187d79b_8b050189,
        64'h191b0187_979b0027,
        64'h571b00c5_17bbc39d,
        64'h8b850017_579b4b98,
        64'h97d2078e_0017861b,
        64'h45914505_47810016,
        64'he913c399_0fe6f913,
        64'h8b89c719_89360017,
        64'hf7130a79_c683008a,
        64'h4783b5c9_e50ff0ef,
        64'h02050513_00005517,
        64'h85ca0126_7a63963e,
        64'h09d9c783_9e3d0087,
        64'h979b0106_161b09e9,
        64'hc78309f9_c603ee05,
        64'h1ae3842a_f8aff0ef,
        64'h852685ce_ee068de3,
        64'h02850513_00005517,
        64'h8a89000b_8963fa65,
        64'h96e387ae_06110521,
        64'h0128893b_0ffbfb93,
        64'h00fbebb3_00be17bb,
        64'hcb898b85_0107c783,
        64'h97d2078e_02080063,
        64'h01162023_02e858bb,
        64'hb7f14b81_4a814c81,
        64'hb7c9ed6f_f0ef0465,
        64'h05130000_55170008,
        64'h8d6302e8_78bb0017,
        64'h859b0005_28034311,
        64'h4e054781_89568662,
        64'h00ca0513_8c0a009c,
        64'h9c9be399_4b8502ea,
        64'hdabb54dc_b7615429,
        64'hf14ff0ef_04c50513,
        64'h00005517_cb8902ec,
        64'hf7bb0005_ac83e791,
        64'h02eaf7bb_060a8063,
        64'hfe09f993_02f10993,
        64'h0045aa83_db4504e5,
        64'h05130000_55170984,
        64'ha7038082_2a010113,
        64'h23813d83_24013d03,
        64'h24813c83_25013c03,
        64'h25813b83_26013b03,
        64'h26813a83_27013a03,
        64'h27813983_28013903,
        64'h28813483_29013403,
        64'h29813083_8522f840,
        64'h0413f8ef_f0ef0765,
        64'h05130000_5517e7b9,
        64'h0016f793_07e4c683,
        64'h00e7eb63_05450513,
        64'h00005517_8a2e8b32,
        64'h84aabfe7_87933ffc,
        64'h07b79f3d_bff7879b,
        64'hbffc07b7_4d180ac7,
        64'hed634789_23b13c23,
        64'h25a13023_25913423,
        64'h25813823_25713c23,
        64'h27613023_27513423,
        64'h27413823_27313c23,
        64'h29213023_28913423,
        64'h28813823_28113c23,
        64'hd6010113_80826145,
        64'h69a26942_64e27402,
        64'h70a28522_013505a3,
        64'h17a010ef_8526842a,
        64'h86dff0ef_852685ca,
        64'h00091c63_00f51e63,
        64'h842a57b5_c519cc1f,
        64'hf0ef84aa_45850b30,
        64'h06138edd_892e9be1,
        64'h0079f693_0ff5f993,
        64'h08154783_f022f406,
        64'he44ee84a_ec267179,
        64'hbfd984aa_b7554685,
        64'hfef760e3_54a94705,
        64'hffc5879b_80822401,
        64'h01132281_34832201,
        64'h39038526_23013403,
        64'h23813083_df400493,
        64'he3990b94_4783e915,
        64'h9a7ff0ef_854a85a2,
        64'h980101f1_0413ed91,
        64'h258199f5_ffe4059b,
        64'he11d84aa_d3fff0ef,
        64'h892a4585_0b900613,
        64'h842eed85_54a94681,
        64'h04b7ec63_06f58463,
        64'h47892321_30232291,
        64'h34232281_38232211,
        64'h3c23dc01_0113b765,
        64'h5929b775_5951bf45,
        64'h1a04b023_5f0020ef,
        64'hdd4d1a04_b503892a,
        64'hb75d08f4_aa2302f7,
        64'h07bb2785_27058bfd,
        64'h8b7d0057_d79b00a7,
        64'hd71b50fc_f3dd8b85,
        64'h0af44783_80822501,
        64'h01132281_39832301,
        64'h39032381_3483854a,
        64'h24013403_24813083,
        64'h08f48023_0a744783,
        64'h08f4ac23_00a7979b,
        64'h02e787bb_0dd44703,
        64'h0e044783_f8dc07a6,
        64'h0d442783_00098663,
        64'hc79954dc_08f4aa23,
        64'h00a7979b_0e044783,
        64'h0af407a3_4785e141,
        64'he0bff0ef_85264585,
        64'h0af00613_4685c6b5,
        64'he3918bfd_09c44783,
        64'hc7898b85_0a044783,
        64'hf4fc07a6_c319f4fc,
        64'h54d89fb9_08844703,
        64'h9fb90087_171b0894,
        64'h47039fb9_0107171b,
        64'h0187979b_08a44703,
        64'h08b44783_f8fc07ce,
        64'h02e787b3_0dd44783,
        64'h02f70733_0e044703,
        64'h97ba08c4_47039fb9,
        64'h0087171b_0107979b,
        64'h468508d4_470308e4,
        64'h47830409_8f63fce5,
        64'h14e30621_070de21c,
        64'h07ce02b7_87b30dd4,
        64'h478302f5_85b30e04,
        64'h45830009_8c634685,
        64'hc39197ae_ffe74583,
        64'h9fad0105_959b0087,
        64'h979b0007_4583fff7,
        64'h4783e0fc_07c64681,
        64'h09d40513_0a844783,
        64'hfcdc07c6_0c848613,
        64'h09140713_0e244783,
        64'h06f48fa3_09c44783,
        64'hc7898b89_0a044783,
        64'h00098a63_08f480a3,
        64'h0b344783_c7890e24,
        64'h4783e781_0019f993,
        64'h8b8506f4_8f2309b4,
        64'h49830a04_4783f8dc,
        64'h00d77363_0147d693,
        64'h07a68007_07136705,
        64'h0d442783_00e7fd63,
        64'hcc981ff7_87934004,
        64'h07b753b8_97ba078a,
        64'h04070713_00004717,
        64'h1cf76d63_47210c04,
        64'h478313d0_10ef85a2,
        64'h20000613_1e050563,
        64'h1a04b503_1aa4b023,
        64'h792020ef_20000513,
        64'he7991a04_b7831e05,
        64'h1a63892a_c03ff0ef,
        64'h84aa85a2_980101f1,
        64'h04131ce7_f3634901,
        64'h3ffc0737_23313423,
        64'h22913c23_24813023,
        64'h24113423_9fb92321,
        64'h3823bffc_07b7db01,
        64'h01134d18_bfcdfc79,
        64'h347d8082_612174a2,
        64'h744270e2_d8bff0ef,
        64'h85263e80_0593e919,
        64'hc4dff0ef_8526858a,
        64'h4601440d_c432c23e,
        64'h84aafc06_f426f822,
        64'h47f58e55_00f11023,
        64'h030006b7_8e554799,
        64'h71390106_161b0086,
        64'h969b8082_61216aa2,
        64'h6a4269e2_74a27902,
        64'h85267442_70e2fc09,
        64'h99e39aa2_02878433,
        64'h9a224089_89b308c9,
        64'h6783fc85_1ae3f01f,
        64'hf0ef854a_85d68652,
        64'h86a2844e_0089f363,
        64'h0207e403_01093783,
        64'h89a6f96d_ecdff0ef,
        64'h854a08c9_2583a089,
        64'h4481bd7f_f0ef4565,
        64'h05130000_551700b6,
        64'h7a630144_85b36810,
        64'h00054d63_905fa0ef,
        64'h852200b4_4583c11d,
        64'h892a4a40_10ef8ab6,
        64'h84b28a2e_4148842a,
        64'hce05e456_e852ec4e,
        64'hf04af426_f822fc06,
        64'h7139b7c5_4401b7d5,
        64'h0004841b_b74d02f6,
        64'h063bbf61_47c58082,
        64'h61256906_64a66446,
        64'h60e68522_c41ff0ef,
        64'h4a050513_00005517,
        64'hc11dd4ff_f0efd23e,
        64'hd402854a_100c47f5,
        64'h460102f1_102347b1,
        64'h0497f063_4785e529,
        64'h842ad6ff_f0efc83e,
        64'hca26d23a_854a100c,
        64'h47850030_cc3ee42e,
        64'h4755d432_cf3108c9,
        64'h27832601_02f11023,
        64'h02c92703_47c906d7,
        64'hf66384b6_892a4785,
        64'he8a2ec86_e0cae4a6,
        64'h711d8082_4501bfd5,
        64'h45018082_612174a2,
        64'h744270e2_f8ed34fd,
        64'hc901dc7f_f0ef8522,
        64'h858a4601_4495cb91,
        64'h8b891b84_2783c11d,
        64'hdddff0ef_c23e842a,
        64'hf426fc06_f822858a,
        64'h460147d5_c42e00f1,
        64'h102347c1_7139e7a9,
        64'h19c52783_bf6df920,
        64'h0513d07f_f0ef5465,
        64'h05130000_5517fc80,
        64'h47e34501_8456b74d,
        64'h84566080_20ef3e80,
        64'h05130080_5863fff4,
        64'h0a9bfe04_c5e334fd,
        64'h80826125_7b027aa2,
        64'h7a4279e2_690664a6,
        64'h644660e6_fba00513,
        64'hd4dff0ef_57450513,
        64'h00005517_c7950125,
        64'hf7b30547_95630135,
        64'hf7b3c789_1005f793,
        64'h45b2ed15_e71ff0ef,
        64'h855a858a_4601e00a,
        64'h0a13e009_89930809,
        64'h09134495_c43e842e,
        64'h8b2af456_ec86f05a,
        64'he4a6e8a2_6a056989,
        64'hfdf94937_0107979b,
        64'hf852fc4e_e0ca07c5,
        64'h5783c23e_47d500f1,
        64'h102347b5_711d8082,
        64'h61457402_70a2c43c,
        64'h47b2e119_ec9ff0ef,
        64'h8522858a_4601c43e,
        64'h8fd94000_07378fd9,
        64'h8f756000_06b78ff5,
        64'h8ff9f806_86934bdc,
        64'h008006b7_4538691c,
        64'hc195842a_c402c23e,
        64'hf406f022_478500f1,
        64'h10234785_71798082,
        64'h61457402_70a28522,
        64'h6fe020ef_7d000513,
        64'he509842a_f21ff0ef,
        64'hc202c402_00011023,
        64'h858a4601_852271c0,
        64'h20eff406_3e800513,
        64'h842af022_71798082,
        64'h4501bf65_4501fd45,
        64'h59b010ef_0d448513,
        64'h0d440593_4611fcf7,
        64'h15e30e04_47830e04,
        64'hc703fcf7_1be30c04,
        64'h47830c04_c703fef7,
        64'h11e30dd4_47830dd4,
        64'hc7038082_24010113,
        64'h22813483_23013403,
        64'h23813083_fb600513,
        64'h00f70d63_0a044783,
        64'h0a04c703_e909fadf,
        64'hf0ef1a05_34832211,
        64'h3c232291_342385a2,
        64'h980101f1_04132281,
        64'h3823dc01_011308e6,
        64'he0634004_07374d14,
        64'h80826161_60a6fd3f,
        64'hf0efcc3e_d402e486,
        64'h100c2000_07930030,
        64'he83ee42e_07851782,
        64'h4785d23e_47d502f1,
        64'h102347a1_715d8302,
        64'h0007b303_679c691c,
        64'h808271a5_05130000,
        64'h55178082_6108953e,
        64'h817549a7_87930000,
        64'h47971502_00a7eb63,
        64'h47ad8082_557d8082,
        64'h01416402_60a24501,
        64'h83020141_60a26402,
        64'h85220003_07630207,
        64'hb303679c_681c0005,
        64'h5e63ff5f_f0ef842a,
        64'he406e022_11418082,
        64'h557d8082_557db7f1,
        64'h659c95aa_058e05e1,
        64'h35f1bfe1_617cbff1,
        64'h7d5c8082_61054501,
        64'h6442e900_64a260e2,
        64'h02945433_0e7010ef,
        64'h90811482_7540f55c,
        64'h08c52483_795c8782,
        64'h97b6e426_e822ec06,
        64'h1101431c_97360025,
        64'h97135026_86930000,
        64'h469704b7_ec63479d,
        64'h80824501_83020003,
        64'h03630087_b303679c,
        64'h691c8082_61356452,
        64'h60f28522_157020ef,
        64'h0808842a_e3fff0ef,
        64'he436eec6_eac2e6be,
        64'he2baea22_ee060808,
        64'h10000593_1234862a,
        64'hfe36fa32_f62e710d,
        64'h80826161_60e2e69f,
        64'hf0efe436_e4c6e0c2,
        64'hfc3ef83a_ec061000,
        64'h05931014_862ef436,
        64'hf032715d_80826161,
        64'h60e2e8df_f0efe436,
        64'he4c6e0c2_fc3ef83a,
        64'hec061034_f436715d,
        64'hb7f18522_02010393,
        64'h0005059b_501010ef,
        64'h85220124_74336000,
        64'h00840b13_b5fd845a,
        64'hd89ff0ef_00840b13,
        64'h02010393_00044503,
        64'ha809dd1f_f0ef0028,
        64'h02010393_0005059b,
        64'he31ff0ef_400845a9,
        64'h46010016_b6930038,
        64'h00840b13_f8b50693,
        64'ha81145c1_00163613,
        64'h46850038_00840b13,
        64'hfa850613_f6e510e3,
        64'h07800713_02e50063,
        64'h07500713_a00d4601,
        64'h46850038_00840b13,
        64'hf6e51ee3_07000713,
        64'h00a76c63_06e50e63,
        64'h07300713_b74d048d,
        64'h0024c503_80826109,
        64'h0007051b_6b066aa6,
        64'h6a4669e6_790674a6,
        64'h744670e6_f55d08f5,
        64'h09630630_079304d5,
        64'h0f630580_069302a6,
        64'heb6306d5_0f630640,
        64'h06930489_0014c503,
        64'h478100f6_f36346a5,
        64'h0ff7f793_fd07879b,
        64'hcb9d0004_c7830355,
        64'h10634781_04890545,
        64'h0f630014_c503bfe1,
        64'he71ff0ef_02010393,
        64'h04850135_086304d7,
        64'hff639381_17827682,
        64'h0017079b_c52d8f1d,
        64'h0004c503_77a27742,
        64'h02095913_03000a93,
        64'h06c00a13_02500993,
        64'hf82af02e_f42afc3e,
        64'h843684b2_e0dafc86,
        64'he4d6e8d2_eccef4a6,
        64'hf8a2597d_011cf0ca,
        64'h7119b7e1_01178023,
        64'h00660023_06850006,
        64'h48830007_c30300d7,
        64'h063397ba_93811782,
        64'h40f807bb_b7d1feb5,
        64'h0fa30505_bf4500c8,
        64'h063b8082_00b7ea63,
        64'h0006879b_fff5081b,
        64'h46810015_559b9d19,
        64'h00050023_050500f5,
        64'h002302d0_07930003,
        64'h076302f6_e96300a6,
        64'h06bb0300_059340e0,
        64'h063b8536_fcb8ffe3,
        64'h02b8d53b_fec68fa3,
        64'h06850ff6_76130306,
        64'h061b04ae_6a630ff5,
        64'h761302b8_f53b0005,
        64'h089b3859_86ba4e25,
        64'h0ff6f813_04100693,
        64'hc2190610_06934305,
        64'h40a0053b_e6810005,
        64'h56634301_bfd900d7,
        64'h00230785_0006c683,
        64'h00f506b3_00d3b823,
        64'h00170693_8082852e,
        64'h00070023_00b6e663,
        64'h0103b703_0007869b,
        64'h47819d9d_fff7059b,
        64'h00c6f563_8e9dfff7,
        64'h06930003_b7038f99,
        64'h92010205_96130103,
        64'hb7830083_b7038082,
        64'h45018082_00078023,
        64'h45050103_b78300a7,
        64'h002300f3_b8230017,
        64'h079300d7_fe639381,
        64'h17822785_40f707b3,
        64'h0003b683_0083b783,
        64'h0103b703_80826145,
        64'h45016a02_69a26942,
        64'h64e27402_70a22f20,
        64'h00ef0d25_05130000,
        64'h6517fd24_1de33020,
        64'h00ef8191_00f5f613,
        64'h0405854e_0007c583,
        64'h008487b3_318000ef,
        64'h8552e781_0004059b,
        64'h01f47793_20000913,
        64'hb2898993_00006997,
        64'hb28a0a13_00006a17,
        64'h4401ed9f_f0ef8526,
        64'h45813460_00efb265,
        64'h05130000_6517dfe6,
        64'h06130000_6617e789,
        64'haa060613_00006617,
        64'h584c19c4_2783e01f,
        64'hb0ef14a5_85930000,
        64'h65977448_13c030ef,
        64'hb4850513_00006517,
        64'h384000ef_b3c50513,
        64'h00006517_ac458593,
        64'h00006597_c789ad65,
        64'h85930000_6597545c,
        64'h3a4000ef_b4c50513,
        64'h00006517_5c0c3b20,
        64'h00ef0186_561b0ff6,
        64'hf6930ff7_77130ff6,
        64'h77930106_569b0086,
        64'h571bb5a5_05130000,
        64'h651706c4_45835830,
        64'h3dc000ef_91c115c2,
        64'h0085d59b_b6450513,
        64'h00006517_546c3f20,
        64'h00efb5a5_05130000,
        64'h651706f4_45834020,
        64'h00ef638c_b5c50513,
        64'h00006517_681c2240,
        64'h10ef842a_4bf010ef,
        64'h45014790_10ef0001,
        64'hb5031ea0_30efb765,
        64'h05130000_651784aa,
        64'h0e2030ef_e052e44e,
        64'he84aec26_f022f406,
        64'h20000513_71797a00,
        64'h006f6105_468560e2,
        64'h66226442_85a25010,
        64'h10efe42e_ec064501,
        64'h842ae822_11018082,
        64'h01416402_60a2557d,
        64'he3914505_703c1a80,
        64'h30efb125_05130000,
        64'h6517b025_85930000,
        64'h659734c0_06139ae6,
        64'h86930000_569702f4,
        64'h02632000_07b7e406,
        64'h6380e022_1141711c,
        64'h80822501_638897aa,
        64'h200007b7_050ef73f,
        64'hf06f2000_05374581,
        64'h46098082_b7f9c45c,
        64'h4785d8f1_45018885,
        64'hbfe94501_c45c4789,
        64'hc7890024_f793f404,
        64'h01242423_e01c2000,
        64'h07b78082_614569a2,
        64'h694264e2_740270a2,
        64'h557d1f60_30ef8522,
        64'h00099d63_508000ef,
        64'hc2050513_00006517,
        64'h862285aa_89aa7b30,
        64'h10efa125_05130000,
        64'h551785a2_c41d5551,
        64'h842a1dc0_30ef892e,
        64'h84b2e44e_f406e84a,
        64'hec26f022_04800513,
        64'h717908b0_41635535,
        64'hb7dd87ca_14e109a1,
        64'h3c2020ef_e43e002c,
        64'h4621854e_639c0087,
        64'h8913dcd5_01096483,
        64'h00093983_97a667a1,
        64'hbf41b1bf_f0ef8522,
        64'hb77100f9_26230009,
        64'hb783dbd9_8b85bd85,
        64'h677020ef_4505d809,
        64'h8ce3c43f_f0ef8522,
        64'h484cc85c_9bf54985,
        64'h485cb4bf_f0ef8522,
        64'hef8d8b85_00892783,
        64'h00090963_04043023,
        64'h2ea030ef_855a85d6,
        64'h0ca00613_aa468693,
        64'h00005697_01848c63,
        64'h04043903_6004cc9d,
        64'h49858889_c85c9bf9,
        64'h485cc85c_0027e793,
        64'h485ccbb5_603cfeb6,
        64'h90e30791_872a2685,
        64'hc3988f51_8361ff87,
        64'h37030106_8763c390,
        64'h0086161b_ff870513,
        64'h63104591_480d4681,
        64'h00c90793_01898713,
        64'h08e69f63_0037f693,
        64'h470d0204_3c230049,
        64'h2783cba9_7c1c3680,
        64'h30ef855a_85d609c0,
        64'h0613b0a6_86930000,
        64'h56970189_8c630384,
        64'h39030004_3983cfb5,
        64'h0014f793_660000ef,
        64'hd5050513_00006517,
        64'h85cad1bf_f0ef85ca,
        64'h29010049_6913ff39,
        64'h79138522_01442903,
        64'hc39d0084_f79368a0,
        64'h00efd525_05130000,
        64'h651785ca_d45ff0ef,
        64'h85ca2901_00896913,
        64'hff397913_85220144,
        64'h2903c39d_0044f793,
        64'hb29ff0ef_85224581,
        64'hb71ff0ef_85224581,
        64'hcc5cf920_0793c781,
        64'h7c1c00f7_6f630c89,
        64'h37830209_37031404,
        64'h80632481_8cfd4981,
        64'h485c0709_34834180,
        64'h30ef855a_85d60f20,
        64'h061386e6_01890963,
        64'h00043903_b7117020,
        64'h00efdb25_05130000,
        64'h6517ba25_85930000,
        64'h5597000b_9d633bfd,
        64'h20000c37_8bd2bd61,
        64'h00c4e493_bd854580,
        64'h30efdc25_05130000,
        64'h6517db25_85930000,
        64'h65971490_0613bbe6,
        64'h86930000_5697b765,
        64'h47014781_2585e31c,
        64'h97469381_83751782,
        64'h170200be_873b8fd9,
        64'h8fe90107_67330087,
        64'hd79b01c8_78330087,
        64'h981b0107_67330187,
        64'h971b0187_d81bf2e5,
        64'h00670363_16fd0605,
        64'h27810107_e7b301e8,
        64'h183b0705_00371f1b,
        64'h00064803_ec0689e3,
        64'h6e89f005_051300ff,
        64'h0e374311_47014781,
        64'h45816390_0107e683,
        64'h65410004_3883603c,
        64'hee079be3_8b85449c,
        64'hdf5ff0ef_8522488c,
        64'hdb9ff0ef_e0248522,
        64'h44cc8082_61654501,
        64'h6ce27c02_7ba27b42,
        64'h7ae26a06_69a66946,
        64'h64e67406_70a6efe9,
        64'h485ce92b_0b130000,
        64'h6b17e82a_8a930000,
        64'h6a97ebbf_f0ef2581,
        64'h0015e593_cccc8c93,
        64'h00005c97_85220d89,
        64'hb583cdbf_f0ef8522,
        64'h4585e9bf_f0ef8522,
        64'h24058593_000f45b7,
        64'hd31ff0ef_85224581,
        64'h46054685_4705cfff,
        64'hf0ef8522_4581cc7f,
        64'hf0ef8522_85a6c8bf,
        64'hf0ef681a_0a138522,
        64'h00095583_c55ff0ef,
        64'h00989a37_85220089,
        64'h2583be3f_f0ef8522,
        64'h4581d73f_f0ef8522,
        64'h45814605_46814705,
        64'h0144e493_16078663,
        64'h8b85008a_2783000a,
        64'h09638cdd_03243c23,
        64'h4c1c4485_e391448d,
        64'h8b89c709_0017f713,
        64'h44810049_278316f9,
        64'h9a630404_3a032000,
        64'h07b70004_3983bf7f,
        64'hf0ef4585_60080e04,
        64'h9c636f60_20ef00c9,
        64'h05134581_4611d01c,
        64'he03084b2_892e0005,
        64'hd7830204_08a3ec66,
        64'hf062f45e_f85afc56,
        64'he0d2e4ce_f486e8ca,
        64'heca67100_f0a27159,
        64'h80826105_690264a2,
        64'h644260e2_c8440499,
        64'h3c2364c0_30effb65,
        64'h05130000_6517fa65,
        64'h85930000_65970760,
        64'h0613da26_86930000,
        64'h569702f9_026384ae,
        64'h842a2000_07b7ec06,
        64'he426e822_00053903,
        64'he04a1101_80826105,
        64'h64a26442_60e2e424,
        64'h692030ef_ffc50513,
        64'h00006517_fec58593,
        64'h00006597_06f00613,
        64'hdd868693_00005697,
        64'h02f40263_84ae2000,
        64'h07b7ec06_e4266100,
        64'he8221101_80826105,
        64'h64a26442_60e2e0a0,
        64'h90511452_6d6030ef,
        64'h04050513_00006517,
        64'h03058593_00006597,
        64'h06800613_e0c68693,
        64'h00005697_02f48263,
        64'h842e2000_07b7ec06,
        64'he8226104_e4261101,
        64'h80826105_64a26442,
        64'h60e2fc80_90411442,
        64'h71a030ef_08450513,
        64'h00006517_07458593,
        64'h00006597_06100613,
        64'he4068693_00005697,
        64'h02f48263_842e2000,
        64'h07b7ec06_e8226104,
        64'he4261101_d4dff06f,
        64'h01414581_60a26402,
        64'h6008f23f_f0ef4605,
        64'h46854705_45818522,
        64'hef1ff0ef_45818522,
        64'hf39ff0ef_842a4581,
        64'h04053023_02053c23,
        64'h46054681_4705e022,
        64'he4061141_80820141,
        64'h45016402_60a2d97f,
        64'hf0ef4581_6008f67f,
        64'hf0ef4581_46054685,
        64'h47058522_f35ff0ef,
        64'h45818522_f7dff0ef,
        64'he4064581_85224605,
        64'h46814705_7100e022,
        64'h11418082_612169e2,
        64'h790274a2_744270e2,
        64'h0289b823_8c4588a1,
        64'h01246433_0034949b,
        64'h8c590049_79130029,
        64'h191b8b05_88090014,
        64'h141b6722_7fe030ef,
        64'he43a16a5_05130000,
        64'h651715a5_85930000,
        64'h659705a0_0613f166,
        64'h86930000_569702f9,
        64'h84638436_893284ae,
        64'h200007b7_fc06f04a,
        64'hf426f822_00053983,
        64'hec4e7139_80826105,
        64'h64a26442_60e2f404,
        64'h04b030ef_1b450513,
        64'h00006517_1a458593,
        64'h00006597_05300613,
        64'hf5068693_00005697,
        64'h02f40263_84ae2000,
        64'h07b7ec06_e4266100,
        64'he8221101_80826105,
        64'h64a26442_60e2f004,
        64'h08b030ef_1f450513,
        64'h00006517_1e458593,
        64'h00006597_04c00613,
        64'hf8068693_00005697,
        64'h02f40263_84ae2000,
        64'h07b7ec06_e4266100,
        64'he8221101_80826105,
        64'h64a26442_60e2ec80,
        64'h90011402_0cf030ef,
        64'h23850513_00006517,
        64'h22858593_00006597,
        64'h04500613_e1468693,
        64'h00007697_02f48263,
        64'h842e2000_07b7ec06,
        64'he8226104_e4261101,
        64'h80826105_64a26442,
        64'h60e2e880_90011402,
        64'h113030ef_27c50513,
        64'h00006517_26c58593,
        64'h00006597_03e00613,
        64'he6068693_00007697,
        64'h02f48263_842e2000,
        64'h07b7ec06_e8226104,
        64'he4261101_80826105,
        64'h64a26442_60e2e404,
        64'h153030ef_2bc50513,
        64'h00006517_2ac58593,
        64'h00006597_03600613,
        64'h03868693_00005697,
        64'h02f40263_84ae2000,
        64'h07b7ec06_e4266100,
        64'he8221101_80826105,
        64'h64a26442_60e2e004,
        64'h193030ef_2fc50513,
        64'h00006517_2ec58593,
        64'h00006597_02f00613,
        64'h06868693_00005697,
        64'h02f40263_84ae2000,
        64'h07b7ec06_e4266100,
        64'he8221101_80826105,
        64'h64a26442_60e2fc24,
        64'h1d3030ef_33c50513,
        64'h00006517_32c58593,
        64'h00006597_08800613,
        64'h09068693_00005697,
        64'h02f50263_84ae842a,
        64'h200007b7_ec06e426,
        64'he8221101_8082556d,
        64'hbfe50007_ac238082,
        64'h4501cf98_02000713,
        64'h00d71763_469100d7,
        64'h0d63711c_46a15958,
        64'h80826149_640a60aa,
        64'hf83ff0ef_0808f01f,
        64'hf0ef0808_e85ff0ef,
        64'h080885a2_6622f71f,
        64'hf0efe42e_e5060808,
        64'h842ae122_71758082,
        64'h61051625_05130000,
        64'h751760e2_fca71de3,
        64'hfef68fa3_fec68f23,
        64'h0007c783_97ae0006,
        64'h46038bbd_962e0047,
        64'hd6130705_06890007,
        64'hc78300e1_07b34541,
        64'h3c858593_00006597,
        64'h1a068693_00007697,
        64'h47013e50_20efec06,
        64'h850a4641_05050593,
        64'h11018082_e13cb807,
        64'h87930000_0797ed3c,
        64'h639cf927_87930000,
        64'h7797e93c_04053423,
        64'h639cf9a7_87930000,
        64'h77978082_614569a2,
        64'h694264e2_740270a2,
        64'hfd24fde3_45019782,
        64'h8522603c_fc1c078e,
        64'h643c0124_f5633f30,
        64'h20ef9522_45819201,
        64'h16020006_091b40a9,
        64'h863b449d_04000993,
        64'h00e78023_97a2f800,
        64'h07130017_8513e84a,
        64'hf406e44e_ec26842a,
        64'h03f7f793_f0227179,
        64'h653c8082_61616ba2,
        64'h6b426ae2_7a0279a2,
        64'h794274e2_640660a6,
        64'hb7c99782_44018526,
        64'h60bc0174_176399d6,
        64'h41590933_4a7020ef,
        64'h0144043b_86560084,
        64'h853385ce_020ada93,
        64'h020a1a93_00090a1b,
        64'h00f97463_93811782,
        64'h00078a1b_408b07bb,
        64'h04000b93_04000b13,
        64'he53c8932_89ae84aa,
        64'h97b203f7_f413ec56,
        64'hf052e486_e45ee85a,
        64'hf44ef84a_fc26e0a2,
        64'h715d653c_80826105,
        64'h692264c2_cd70cd34,
        64'hc97c0505_282300c8,
        64'h863b00d3_06bb00fe,
        64'h07bb010e_883b6462,
        64'hf3ff1de3_00e587bb,
        64'h0005869b_0003861b,
        64'h0f918f5d_0157171b,
        64'h00b7579b_9f3d0077,
        64'h47339fa1_8f4dfff7,
        64'h47130007_081b00b3,
        64'h85bb4080_9fa18dd5,
        64'h0115d59b_94aa00f5,
        64'h969b048a_9db5ffc2,
        64'ha4038db9_02c10075,
        64'he5b3fff7_c593023f,
        64'hc4839ead_00c703bb,
        64'h00c3e633_400c9ead,
        64'h0166561b_00a6139b,
        64'h0082a583_9e2d8e3d,
        64'h8e59fff6_c6139db1,
        64'h00f8073b_01076833,
        64'h01a8581b_0003a583,
        64'h9e2d0068_171b0107,
        64'h083b0042_a5839f2d,
        64'h942a040a_418c95aa,
        64'h058a93aa_038a020f,
        64'hc5839f2d_022fc403,
        64'h021fc383_0002a703,
        64'h00d745b3_8f5dfff6,
        64'h47132e22_82930000,
        64'h5297f45f_17e300e4,
        64'h07bb0004_069b0005,
        64'h861b0291_8f5d0177,
        64'h171b0097_579b9f3d,
        64'h8f219fa5_8f2d0007,
        64'h081b00d5_843b8ec1,
        64'h00092483_0106d69b,
        64'h9fa50106_941b992a,
        64'h9ea1090a_8ead00e7,
        64'hc6b3ffc3_a4839c35,
        64'h00c705bb_03c18e4d,
        64'h0156561b_0132c903,
        64'h00b6159b_40809e2d,
        64'h9ea194aa_8db9048a,
        64'h00f8073b_0083a403,
        64'h9e210107_683301c8,
        64'h581b0048_171b0122,
        64'hc4830107_083b4080,
        64'h9e2194aa_048a0043,
        64'ha4039f21_0112c483,
        64'h9f254000_00c5c4b3,
        64'h942a040a_00d7c5b3,
        64'h0003a703_0102c403,
        64'h36038393_00005397,
        64'h82fe3eaf_8f930000,
        64'h5f97f25f_1ee300e4,
        64'h07bb0004_069b0003,
        64'h861b0005_881b8f5d,
        64'h0147171b_00c7579b,
        64'h9f3d0077_47338f6d,
        64'h0083c733_9fb900d3,
        64'h843b8ec1_40980126,
        64'hd69b9fb9_00e6941b,
        64'h94aa048a_ffcfa703,
        64'h9eb90fc1_8eadffff,
        64'h44838efd_0075c6b3,
        64'h0f119f35_00c583bb,
        64'h00c3e633_40189eb9,
        64'h0176561b_0096139b,
        64'h008fa703_9e398e3d,
        64'h8e7500b7_c6339f31,
        64'h00f805bb_0105e833,
        64'h0003a703_01b8581b,
        64'h9e390058_159b0105,
        64'h883b004f_a7039db9,
        64'h942a040a_4318972a,
        64'h070a93aa_038a000f,
        64'h47039db9_002f4403,
        64'h001f4383_000fa583,
        64'h00b6c733_8df100d7,
        64'hc5b34ca2_82930000,
        64'h5297402f_8f930000,
        64'h5f974caf_0f130000,
        64'h5f17f45f_17e300e3,
        64'h87bb0003_869b0005,
        64'h881b0f41_8f5d0167,
        64'h171b00a7_579b9f3d,
        64'h8f2d9fa1_00777733,
        64'h8f2d0007_061b00d7,
        64'h03bbffcf_a4039fa1,
        64'h00d3e6b3_0116969b,
        64'h00f6d39b_007686bb,
        64'h8ebd00cf_24038ef9,
        64'h00b7c6b3_00d383bb,
        64'h00c5873b_008383bb,
        64'h8e590146_561b00c6,
        64'h171b9e39_008f2383,
        64'h8e358e6d_00f6c633,
        64'h9f3100f8_05bb0077,
        64'h073b0105_e8330198,
        64'h581b0078_159b0105,
        64'h883b004f_2703ff4f,
        64'ha3839db9_007585bb,
        64'h0fc1008f_a403000f,
        64'h2583000f_a38300b6,
        64'h47338dfd_00c6c5b3,
        64'h488f8f93_00005f97,
        64'h887687f2_869a8646,
        64'h04050293_8f2ae44a,
        64'he826ec22_110105c5,
        64'h28830585_23030545,
        64'h2e030505_2e83bf81,
        64'h842abdd1_00e785a3,
        64'h47216786_a8dfd0ef,
        64'h082c462d_6506ab7f,
        64'hd0ef4581_02000613,
        64'h6506f835_0005041b,
        64'ha19fe0ef_1028d3c1,
        64'h01814783_02f51b63,
        64'h4791b771_0005041b,
        64'h8b2fe0ef_00f50223,
        64'h47857522_00f50023,
        64'h5795b7c5_078500c6,
        64'h802396be_0834b77d,
        64'hf0f713e3_0e500793,
        64'h01814703_00d77963,
        64'h0007869b_02000613,
        64'h47299381_02061793,
        64'hf8f6e9e3_0007069b,
        64'h00d58023_070595ba,
        64'h082cfe67_02e3b7dd,
        64'hffc81be3_00080563,
        64'h0005c803_05858082,
        64'h61256446_60e68522,
        64'h4419feb0_45e34185,
        64'hd59b0185_959ba831,
        64'h00068e1b_92c58593,
        64'h00007597_92c116c2,
        64'h36810108_ec630308,
        64'h58131842_f9f6881b,
        64'h92c10305_96930017,
        64'h061b0006_c58300e5,
        64'h06b3432d_48e54701,
        64'hfec686e3_0006c683,
        64'h96aa9281_02071693,
        64'hfff7871b_b77d87ba,
        64'hb7452785_a0e900e7,
        64'h8ca30007_8ba30007,
        64'h8b230460_071300e7,
        64'h8c230210_07136786,
        64'hbb1fd0ef_082c462d,
        64'hc7e56506_01814783,
        64'h10051563_2501ac3f,
        64'he0ef1028_4585e045,
        64'h0005041b_bccfe0ef,
        64'hda021028_4581ebb1,
        64'h02000613_eb290007,
        64'h4703972a_93010207,
        64'h97134781_00010c23,
        64'h6522e471_0005041b,
        64'heddfd0ef_ec86e8a2,
        64'h1028002c_4605e42a,
        64'h711db7d5_842abf55,
        64'h00048023_00f51563,
        64'h47918082_61256906,
        64'h64a66446_60e68522,
        64'h00a92023_c15fd0ef,
        64'h953e0347_87930270,
        64'h079300e6_84630005,
        64'h46830430_0793470d,
        64'h6562e015_0005041b,
        64'he63fd0ef_510c6562,
        64'h02090a63_fec783e3,
        64'h177d0007_c78397a6,
        64'h93811782_0007869b,
        64'hfff6879b_ce890007,
        64'h00230200_061346ad,
        64'h00b48713_c8dfd0ef,
        64'h8526462d_75c2e93d,
        64'h2501b97f_e0ef0828,
        64'h4585e559_2501c9ef,
        64'he0efd202_08284581,
        64'hc4b9e051_0005041b,
        64'hf95fd0ef_ec86e8a2,
        64'h08284601_002c8932,
        64'h84aee42a_e0cae4a6,
        64'h711d8082_61256446,
        64'h60e62501_acefe0ef,
        64'h00f50223_478500e7,
        64'h8ca30087_571b00e7,
        64'h8c230044_570300e7,
        64'h8ba30087_571b00e7,
        64'h8b237522_00645703,
        64'hcb856786_eb950207,
        64'hf79300b7_c7834519,
        64'h67a6e129_250199df,
        64'he0efe4be_1028083c,
        64'h65a2e929_250180af,
        64'he0efec86_1028002c,
        64'h4605842e_e42ae8a2,
        64'h711dbfcd_47a18082,
        64'h614d853e_64ea740a,
        64'h70aa0005_079bb48f,
        64'he0ef6506_e7910005,
        64'h079be18f_e0ef0088,
        64'h00f70223_06d707a3,
        64'h478506f7_04a30086,
        64'hd69b0106_d69b0087,
        64'hd79b0107_d79b0107,
        64'h979b06f7_04230107,
        64'hd79b06f7_07230107,
        64'h969b57d6_02f69c63,
        64'h05574683_02e00793,
        64'h6706efa9_0005079b,
        64'hfbbfd0ef_8522c1bd,
        64'h47890005_059bca4f,
        64'he0ef8522_0005059b,
        64'hf25fd0ef_85a60004,
        64'h450306f7_076357d6,
        64'h4736cbb5_8bc100b4,
        64'hc78300f4_02234785,
        64'h00f485a3_0207e793,
        64'h64060281_4783df7f,
        64'hd0ef00d4_851302a1,
        64'h0593464d_648aebdd,
        64'h0005079b_dcbfe0ef,
        64'h10a80ce7_92634711,
        64'hcbf10005_079ba9df,
        64'he0ef10a8_65820c05,
        64'h4c6347ad_efdfd0ef,
        64'h850ae33f_d0ef10a8,
        64'h008c0280_0613e3ff,
        64'hd0ef1028_05ad4655,
        64'h0e058d63_479165e6,
        64'h10071163_02077713,
        64'h479900b7_c7037786,
        64'h10079963_0005079b,
        64'hae7fe0ef_f0be083c,
        64'hf4be0088_65a26786,
        64'h12079563_0005079b,
        64'h95cfe0ef_ed26f122,
        64'hf5060088_002c4605,
        64'he02ee42a_71718082,
        64'h616564e6_740670a6,
        64'h2501c94f_e0ef00f5,
        64'h02234785_008705a3,
        64'h8c3d0274_74138c65,
        64'h8cbd7522_00b74783,
        64'hc30d6706_e39d0207,
        64'hf79300b7_c7834519,
        64'h67a6e915_2501b55f,
        64'he0efe4be_1028083c,
        64'h65a2e131_25019c2f,
        64'he0eff486_10284605,
        64'h002c8432_84aee42a,
        64'heca6f0a2_7159b7c5,
        64'h44218082_614d6d46,
        64'h6ce67c06_7ba67b46,
        64'h7ae66a0a_69aa694a,
        64'h64ea740a_70aa8522,
        64'hf2bfe0ef_85a67522,
        64'h441db749_8c6a0ffb,
        64'hfb93f53f_d0ef3bfd,
        64'h855a4581_20000613,
        64'hec090005_041b8d4f,
        64'he0ef0195_02230385,
        64'h2823001c_0d1b7522,
        64'ha82d0005_041bd50f,
        64'he0ef00f5_02234785,
        64'h01278aa3_01578a23,
        64'h01378da3_01478d23,
        64'h00e78ca3_00078ba3,
        64'h00078b23_04600713,
        64'h00e78c23_02100713,
        64'h00e785a3_75224741,
        64'h6786e835_0005041b,
        64'hf5ffe0ef_1028040b,
        64'h99634c85_00274b83,
        64'h06f404a3_06d407a3,
        64'h0087d79b_0086d69b,
        64'h0107d79b_0106d69b,
        64'h0107979b_06f40423,
        64'h0107d79b_0107969b,
        64'h06f40723_478100f6,
        64'h93635714_00d61663,
        64'h57d20007_4603468d,
        64'h05740aa3_7722ff7f,
        64'hd0ef0544_051385da,
        64'h052404a3_05540423,
        64'h053407a3_05440723,
        64'h040405a3_04040523,
        64'h03740a23_02000613,
        64'h04f406a3_0089591b,
        64'h0089d99b_04600793,
        64'h0ff4fa13_04f40623,
        64'h02e00b93_0109591b,
        64'h02100793_0109d99b,
        64'h02f40fa3_0109191b,
        64'h0104999b_0ff97a93,
        64'h47c187af_e0ef855a,
        64'h02000593_462d886f,
        64'he0ef855a_00050c1b,
        64'h45812000_06130344,
        64'h0b13f60f_e0ef8522,
        64'h0104d91b_85a67422,
        64'h16041263_0005041b,
        64'ha8cfe0ef_16f48863,
        64'h440557fd_16f48c63,
        64'h44097522_47851804,
        64'h80630005_049bb33f,
        64'he0ef4581_75221807,
        64'h9d630207_f79300b7,
        64'hc7834419_67a61af4,
        64'h15634791_1c040763,
        64'h0005041b_d53fe0ef,
        64'he4be1028_083c65a2,
        64'h1c041263_0005041b,
        64'hbc4fe0ef_e8eaece6,
        64'hf0e2f4de_f8dafcd6,
        64'he152e54e_e94aed26,
        64'hf506f122_1028002c,
        64'h4605e42a_7171b7ed,
        64'hf5512501_91eff0ef,
        64'h85a27502_bf612501,
        64'hf12fe0ef_7502e411,
        64'hf1552501_9e3fe0ef,
        64'h1008faf5_18e34791,
        64'hd94d2501_838ff0ef,
        64'h00a84581_f1612501,
        64'h941fe0ef_caa200a8,
        64'h4589952f_e0ef00a8,
        64'h100c0280_0613fc87,
        64'h8de30149_2783c89d,
        64'h88c1cc0d_0005041b,
        64'haccfe0ef_00094503,
        64'h79028082_61497946,
        64'h74e6640a_60aa451d,
        64'hcb810014_f79300b5,
        64'hc483c599_75e2eb89,
        64'h0207f793_00b7c783,
        64'h45196786_e1052501,
        64'he27fe0ef_e0be1008,
        64'h081c65a2_e9052501,
        64'hc94fe0ef_f8cafca6,
        64'he122e506_1008002c,
        64'h4605e42a_7175b7b1,
        64'h00f40523_fbf7f793,
        64'h00a44783_f55d2501,
        64'h71e040ef_03040593,
        64'h0017c503_46854c50,
        64'h601cdba5_0407f793,
        64'h00a44783_fcf96ae3,
        64'h4d1c6008_fcf900e3,
        64'h45094785_b769449d,
        64'hb7e12501_a1eff0ef,
        64'h85ca6008_f9792501,
        64'hb25fe0ef_167d1000,
        64'h06374c0c_b7dd4505,
        64'h02f91463_57fd0005,
        64'h091b941f_e0ef4c0c,
        64'hbf7d84aa_00a405a3,
        64'hc5390004_2a232501,
        64'ha5aff0ef_484cef01,
        64'h600800f4_0523c818,
        64'h0207e793_fed772e3,
        64'h48144458_cf390027,
        64'hf71300a4_47838082,
        64'h610564a2_69028526,
        64'h644260e2_0007849b,
        64'hcb9100b4_4783e491,
        64'h0005049b_bb8fe0ef,
        64'h842ae04a_ec06e426,
        64'he8221101_bfad8a2a,
        64'hbfbd4a09_b7494a05,
        64'hb7c539f1_09112485,
        64'he1116582_01557533,
        64'h2501aa2f_e0efe02e,
        64'h854ab745_fc0c94e3,
        64'h3cfd39f9_09092485,
        64'he3918fd9_0087979b,
        64'h00094703_00194783,
        64'h038b9163_20000993,
        64'h03440913_85cee921,
        64'h2501d04f_e0ef0015,
        64'h899b8522_00099e63,
        64'h1afd4c09_44814981,
        64'h49011000_0ab7504c,
        64'hb74d009b_202300f4,
        64'h02a30017_e793c804,
        64'h00544783_fef963e3,
        64'h29054c1c_2485e111,
        64'h09550863_09350863,
        64'h2501a49f_e0ef8522,
        64'h85ca4a85_59fd4481,
        64'h490902fb_9f634785,
        64'h00044b83_80826165,
        64'h6ce27c02_7ba27b42,
        64'h7ae26a06_69a66946,
        64'h64e68552_740670a6,
        64'h00fb2023_02f76263,
        64'hffec871b_481c0184,
        64'h2c836000_000a1c63,
        64'h00050a1b_e70fe0ef,
        64'hec66f062_f45efc56,
        64'he4cee8ca_eca6f486,
        64'he0d28522_002c4601,
        64'h8b2ee42a_f85a8432,
        64'hf0a27159_bfcd4419,
        64'h80826165_64e67406,
        64'h70a68522_c00fe0ef,
        64'h102885a6_c489cf81,
        64'h6786e801_0005041b,
        64'h85eff0ef_e4be1028,
        64'h083c65a2_e00d0005,
        64'h041becef_e0eff486,
        64'hf0a21028_002c4601,
        64'h84aee42a_eca67159,
        64'hbf6584aa_d16dbf7d,
        64'h00042a23_00f51663,
        64'h47912501_f77fe0ef,
        64'h85224581_c58fe0ef,
        64'h852285ca_00042a23,
        64'h02f51363_47912501,
        64'hb34ff0ef_85224581,
        64'h02243023_80826145,
        64'h64e26942_85267402,
        64'h70a20005_049bc4ff,
        64'he0ef8522_45810009,
        64'h1f63e889_0005049b,
        64'hd8cfe0ef_892e842a,
        64'hf406e84a_ec26f022,
        64'h71798082_01416402,
        64'h60a20004_3023e119,
        64'h2501daef_e0ef842a,
        64'he406e022_1141b7c1,
        64'hfcf501e3_4791bfdd,
        64'h45258082_61217442,
        64'h70e2f971_fcf50be3,
        64'h47912501_cadfe0ef,
        64'h00f41423_0067d783,
        64'h85224581_67e2c448,
        64'he24fe0ef_0007c503,
        64'h67e2a02d_00043023,
        64'h4515e789_8bc100b5,
        64'hc783cd99_6c0ce529,
        64'h2501968f_f0eff01c,
        64'h101ce01c_852265a2,
        64'h67e2e115_2501fdaf,
        64'he0ef0828_002c4601,
        64'h842ac52d_e42ef822,
        64'hfc067139_b7bdc45c,
        64'h013787bb_413484bb,
        64'hcc0c445c_faf5fae3,
        64'h4f9c601c_fabafee3,
        64'hfd4588e3_0005059b,
        64'hc3ffe0ef_bf6984ce,
        64'he5990005_059bfcbf,
        64'he0efcb81_8b896008,
        64'h00a44783_b765cc0c,
        64'hc84cb5ed_490500f4,
        64'h05a34785_00f59763,
        64'h57fdbded_490900f4,
        64'h05a34789_00f59763,
        64'h47850005_059b802f,
        64'hf0efe595_484cbfb1,
        64'h9ca90094_d49bcd11,
        64'h2501c79f_e0ef6008,
        64'hd7b51ff4_f793c45c,
        64'h9fa5445c_0499ea63,
        64'h4a855a7d_d1c19c9d,
        64'hc45c2781_4c0c8ff9,
        64'h413007bb_02c6ed63,
        64'h0337563b_0336d6bb,
        64'hfff4869b_377dc729,
        64'h0097999b_00254783,
        64'h6008bf59_cc44ed35,
        64'h25012ef0_40ef85ce,
        64'h0017c503_86264685,
        64'h601c00f4_0523fbf7,
        64'hf79300a4_4783ed51,
        64'h25013410_40ef0017,
        64'hc50385ce_4685601c,
        64'hc3850407_f7930304,
        64'h099300a4_4783fc96,
        64'h0ee34c50_d3e51ff7,
        64'hf793445c_4481bf7d,
        64'h00f40523_0207e793,
        64'h00a44783_c81cfcf7,
        64'h78e34818_445ce4bd,
        64'h00042623_445884ba,
        64'he3918b89_00a44783,
        64'h00977763_48188082,
        64'h61216aa2_6a4269e2,
        64'h790274a2_854a7442,
        64'h70e20007_891bcf89,
        64'h00b44783_00091763,
        64'h0005091b_fa8fe0ef,
        64'h84ae842a_e456e852,
        64'hec4efc06_f04af426,
        64'hf8227139_b721fe94,
        64'h65e3fee7_8fa32405,
        64'h07850007_47039736,
        64'h92810204_16936722,
        64'h0789bdf5_4545b7e9,
        64'h00e60023_fc974703,
        64'h972a1088_93011702,
        64'h0007059b_fff5871b,
        64'hb7e12785_bf199c3d,
        64'h01260023_fff7c793,
        64'he989963a_93010206,
        64'h97136622_36fd86a2,
        64'h85be04e4_60630037,
        64'h871be705_fc974703,
        64'h97361094_93010207,
        64'h97134781_f48fe0ef,
        64'h1828100c_b7614509,
        64'hf6e512e3_67a24711,
        64'hdd612501_a86ff0ef,
        64'h18284581_01350e63,
        64'h2501897f_e0ef0007,
        64'hc50365c6_77e2e105,
        64'h2501e46f_f0ef1828,
        64'h4581f951_2501f4ff,
        64'he0ef1828_4581c2aa,
        64'h8bdfe0ef_0007c503,
        64'h65c677e2_f55d2501,
        64'he6cff0ef_18284581,
        64'hfd4d2501_f75fe0ef,
        64'h18284585_80826149,
        64'h79a67946_74e6640a,
        64'h60aa0007_8023078d,
        64'h00e78123_02f00713,
        64'h0e941563_00e780a3,
        64'h03a00713_00e78023,
        64'h0307071b_37474703,
        64'h00008717_e50567a2,
        64'h45010409_91634996,
        64'hc2be4bdc_02f00913,
        64'h842677e2_ecbe081c,
        64'he5212501_ab9fe0ef,
        64'h1828002c_460184ae,
        64'h00050023_f4cef8ca,
        64'he122e506_e42afca6,
        64'h7175bfd9_4415fcf4,
        64'h1ee34791_b7c5c8c8,
        64'h965fe0ef_0004c503,
        64'h74a2cb99_8bc100b5,
        64'hc7838082_616564e6,
        64'h740670a6_8522cbd8,
        64'h575277a2_e9916586,
        64'he41d0005_041bcb4f,
        64'hf0efe4be_1028083c,
        64'h65a2ec19_0005041b,
        64'hb25fe0ef_eca6f486,
        64'hf0a21028_002c4601,
        64'he42a7159_bfe5452d,
        64'h80826105_60e24501,
        64'h42a78423_00008797,
        64'h00054a63_945fe0ef,
        64'hec060028_e42a1101,
        64'h80820141_640260a2,
        64'h00043023_e1192501,
        64'h9b5fe0ef_8522e901,
        64'h2501f01f_f0ef842a,
        64'he406e022_11418082,
        64'h01416402_60a24505,
        64'hea3fe06f_014160a2,
        64'h640200f5_02234785,
        64'h00f40523_fdf7f793,
        64'h600800a4_47830007,
        64'h89a30007_892300e7,
        64'h8ca300d7_8da30460,
        64'h07130086_d69b00e7,
        64'h8c230210_07130106,
        64'hd69b00e7_8aa30087,
        64'h571b0107_571b0107,
        64'h171b00e7_8a230107,
        64'h571b0107_169b00e7,
        64'h8d230007_8ba30007,
        64'h8b234858_00e78fa3,
        64'h00d78f23_0187571b,
        64'h0107569b_00d78ea3,
        64'h00e78e23_0086d69b,
        64'h0106d69b_0107169b,
        64'h481800e7_85a30207,
        64'h671300b7_c703741c,
        64'he1552501_b5ffe0ef,
        64'h6008500c_00f40523,
        64'hfbf7f793_00a44783,
        64'hed4d2501_6ab040ef,
        64'h03040593_0017c503,
        64'h46854c50_601cc395,
        64'h0407f793_cf610207,
        64'hf71300a4_4783e16d,
        64'h2501ab7f_e0ef842a,
        64'he406e022_1141bd15,
        64'h499db5f1_c81cbf41,
        64'h00f40523_0407e793,
        64'h00a44783_9b5fe0ef,
        64'h952285d2_86260305,
        64'h05130007_049b0127,
        64'h746340ab_873b1ff5,
        64'h75130009_049b4448,
        64'h01b42e23_fd012501,
        64'h6ed040ef_85da4685,
        64'h0017c503_00d77a63,
        64'h44584814_00c70e63,
        64'h4c58bdc9_00faa023,
        64'h9fa5000a_a783c45c,
        64'h9fa54099_093b445c,
        64'h9a3e9381_02049793,
        64'h0094949b_00f40523,
        64'hfbf7f793_00a44783,
        64'ha29fe0ef_855a95d2,
        64'h20000613_91811582,
        64'h0097959b_0297f263,
        64'h41b587bb_4c4cf149,
        64'h25017890_40ef85d2,
        64'h86a60017_c50341a6,
        64'h84bb00e6_f4630104,
        64'h873b0099_549b0027,
        64'hc683072c_7a6367a2,
        64'h8db200a8_063b000d,
        64'h081bd159_2501964f,
        64'hf0efe43e_853e4c0c,
        64'h601c00f4_0523fbf7,
        64'hf79300a4_4783f969,
        64'h25017d90_40ef85da,
        64'h0017c503_46854c50,
        64'h601cc38d_0407f793,
        64'h00a44783_c85ce311,
        64'hcc1c4858_bf894985,
        64'h00f405a3_47850197,
        64'h9763b785_00f40523,
        64'h0207e793_00a44783,
        64'h12f76b63_4818445c,
        64'hf3fd0005_079bd6af,
        64'hf0ef4c0c_b7494989,
        64'h00f405a3_478902e7,
        64'h98634705_cb914581,
        64'h485cef01_040d1a63,
        64'h0ffd7d13_01a7fd33,
        64'h37fd0025_47830097,
        64'h5d1b6008_14079463,
        64'h1ff77793_04090463,
        64'h44585cfd_03040b13,
        64'h1ff00c13_20000b93,
        64'h04f76e63_0127873b,
        64'h445c1a07_82638b89,
        64'h00a44783_80826109,
        64'h6de27d02_7ca27c42,
        64'h7be26b06_6aa66a46,
        64'h69e67906_74a6854e,
        64'h744670e6_0007899b,
        64'hc39d00b4_47830009,
        64'h97630005_099bca3f,
        64'he0ef8ab6_89328a2e,
        64'h842a0006_a023ec6e,
        64'hf06af466_f862fc5e,
        64'he0daf4a6_fc86e4d6,
        64'he8d2ecce_f0caf8a2,
        64'h7119b585_499dbf9d,
        64'hbb1fe0ef_855295a2,
        64'h86260305_85930007,
        64'h049b0127_746340bb,
        64'h873b1ff5_f5930009,
        64'h049b444c_01b42e23,
        64'hf10d2501_0e8050ef,
        64'h85da0017_c5038642,
        64'h4685601c_00f40523,
        64'hfbf7f793_682200a4,
        64'h4783f131_250113c0,
        64'h50efe442_85da4685,
        64'h0017c503_c30d0407,
        64'h771300a4_47030506,
        64'h01634c50_bf3900fa,
        64'ha0239fa5_000aa783,
        64'hc45c9fa5_4099093b,
        64'h445c9a3e_93810204,
        64'h97930094_949bc3ff,
        64'he0ef9552_85da2000,
        64'h06139101_15020097,
        64'h951b0097_fc6341b5,
        64'h07bb4c48_c3850407,
        64'hf79300a4_4783f945,
        64'h25011760_50ef85d2,
        64'h864286a6_0017c503,
        64'h41a684bb_00e6f463,
        64'h00c4873b_0099549b,
        64'h0027c683_072c7a63,
        64'h67a28dc2_00a6083b,
        64'h000d061b_d5792501,
        64'hb86ff0ef_e43e853e,
        64'h4c0c601c_cc08b795,
        64'h498500f4_05a34785,
        64'h01951763_b7e52501,
        64'hbc6ff0ef_4c0cbfb5,
        64'h498900f4_05a34789,
        64'h00a7ec63_47854848,
        64'heb11020d_19630ffd,
        64'h7d1301a7_fd3337fd,
        64'h00254783_00975d1b,
        64'h60081207_91631ff7,
        64'h77934458_fa090ae3,
        64'h5cfd0304_0b131ff0,
        64'h0c132000_0b930006,
        64'h091b00f6_7463893e,
        64'h40f907bb_445c0104,
        64'h29031607_8c638b85,
        64'h00a44783_80826109,
        64'h6de27d02_7ca27c42,
        64'h7be26b06_6aa66a46,
        64'h69e67906_74a6854e,
        64'h744670e6_0007899b,
        64'hc39d6622_00b44783,
        64'h00099863_0005099b,
        64'he85fe0ef_8ab6e432,
        64'h8a2e842a_0006a023,
        64'hec6ef06a_f466f862,
        64'hfc5ee0da_f0caf4a6,
        64'hfc86e4d6_e8d2ecce,
        64'hf8a27119_bdd14525,
        64'hbf51ec07_9ee3451d,
        64'h8b85fa09_00e30029,
        64'h7913ee07_16e30107,
        64'hf7134511_00b44783,
        64'hee051de3_bdf54501,
        64'h00f49423_0124b023,
        64'h0004ae23_0004a623,
        64'hc8880069_5783daff,
        64'he0ef01c4_0513c8c8,
        64'hf35fe0ef_00094503,
        64'h000485a3_d09c0134,
        64'h8523f480_03092783,
        64'h85a27922_0209e993,
        64'hc3990089_f793f139,
        64'h250180cf_f0ef0125,
        64'h262385d6_397d7522,
        64'hfd212501_e1fff0ef,
        64'h030a2a83_855285ca,
        64'h02090363_00fa0223,
        64'h0005091b_00040aa3,
        64'h00040a23_00040da3,
        64'h00040d23_4785f9bf,
        64'he0ef85a2_000a4503,
        64'h00040fa3_00040f23,
        64'h00040ea3_00040e23,
        64'h000405a3_00e40c23,
        64'h00040ba3_00040b23,
        64'h00e40823_000407a3,
        64'h00040723_00f40ca3,
        64'h00f408a3_02100713,
        64'h04600793_7a220089,
        64'he9936406_a0210809,
        64'h0a630089_7913fff9,
        64'h45210049_7793f3fd,
        64'h8bc5451d_00b44783,
        64'h80826149_6ae67a06,
        64'h79a67946_74e6640a,
        64'h60aac905_2501e7df,
        64'hf0ef1028_00f51763,
        64'h4791c115_10078e63,
        64'h01f97993_01c97793,
        64'h4519e011_e1196406,
        64'h2501b61f_f0efe4be,
        64'h1028083c_65a2e91d,
        64'h25019cef_f0ef1028,
        64'h002c8a79_84aa8932,
        64'h00053023_16050c63,
        64'he42eecd6_f0d2f4ce,
        64'hf8cafca6_e122e506,
        64'h7175bfe5_452d8082,
        64'h612170e2_2501a02f,
        64'hf0ef0828_080c4601,
        64'h00f61863_4785cb11,
        64'h4501e398_97aa0007,
        64'h0023c319_67620007,
        64'h0023c319_66226318,
        64'h00a78733_050eb067,
        64'h87930000_97970405,
        64'h4263832f_f0eff42e,
        64'he432e82e_fc061028,
        64'hec2a7139_80824509,
        64'hbf4d4505_bf5d4509,
        64'hbf65faf4_e7e30004,
        64'h891b4c1c_00f402a3,
        64'h0017e793_00544783,
        64'hc81c2785_01378a63,
        64'h481cfd71_25018abf,
        64'hf0ef8522_85ca4601,
        64'h03348c63_03448c63,
        64'h80826145_6a0269a2,
        64'h694264e2_740270a2,
        64'h4501e891_0005049b,
        64'hed6ff0ef_852285ca,
        64'h59fd4a05_06f5f063,
        64'h892e842a_e052e44e,
        64'hec26f406_e84af022,
        64'h71794d1c_08b7f063,
        64'h47858082_610564a2,
        64'h85266442_60e200e7,
        64'h82234705_601c80ef,
        64'hf0ef462d_6c08700c,
        64'h838ff0ef_45810200,
        64'h06136c08_e0850005,
        64'h049ba34f_f0ef6008,
        64'h484ce49d_0005049b,
        64'hfa9ff0ef_842aec06,
        64'he426e822_11018082,
        64'h610564a2_644260e2,
        64'h451d00f5_13634791,
        64'hdd792501_bb7ff0ef,
        64'h85224585_cb990097,
        64'h8d630007_c7836c1c,
        64'hed092501_a7eff0ef,
        64'h6008484c_0e500493,
        64'he50d2501_87dff0ef,
        64'h842ae426_ec06e822,
        64'h45811101_bfe54511,
        64'hb7cd0004_2a23d945,
        64'h2501bfdf_f0ef8522,
        64'h45818082_614569a2,
        64'h694264e2_740270a2,
        64'h45010097_9a630017,
        64'hb79317e1_8bfd0337,
        64'h80630327_026303f7,
        64'hf79300b7_c783c321,
        64'h0007c703_6c1ce129,
        64'h2501aecf_f0ef6008,
        64'ha0b1c90d_e199484c,
        64'h49bd0e50_09134511,
        64'h84aef406_842ae44e,
        64'he84aec26_f0227179,
        64'hbdc10ff7_77130017,
        64'he7933701_eca8efe3,
        64'h0ff57513_f9f7051b,
        64'heea8f3e3_0ff57513,
        64'hfbf7051b_b5754519,
        64'hef0719e3_00080663,
        64'h00054803_f1450513,
        64'h00008517_00054c63,
        64'h4185551b_0187151b,
        64'h02b6f263_fd370ae3,
        64'hf35709e3_f3470be3,
        64'hf2e37de3_00074703,
        64'h97229301_17020017,
        64'h061b8732_45ad46a1,
        64'h0ff7f793_0027979b,
        64'h05659a63_b5a1c4c8,
        64'hae4ff0ef_0007c503,
        64'h609cdbe5_8bc100b5,
        64'hc7836c8c_fbe58b91,
        64'hb7054515_f315bfd9,
        64'h4511b72d_4501e607,
        64'h0ae30004_bc230004,
        64'ha623cb99_0207f793,
        64'h0047f713_f4e513e3,
        64'h4711c515_00b7c783,
        64'h709cf127_9de3b7c5,
        64'h01066613_fed714e3,
        64'h46850037_f713bded,
        64'h00c905a3_00866613,
        64'h00e79463_47118bb1,
        64'h0ff7f793_0027979b,
        64'h01659f63_00e90023,
        64'h471500e6_95630e50,
        64'h07130009_4683c6e5,
        64'h460100e5_73634611,
        64'h94320200_05139201,
        64'h1602a865_268500e5,
        64'h0023954a_91010206,
        64'h95130027_e793a211,
        64'h0505a8c9_48e50200,
        64'h03134781_45a14701,
        64'h4681b78d_02400793,
        64'h943a12f6_e7630200,
        64'h0693f757_87e3b7b5,
        64'h4709b73d_04058082,
        64'h61216b02_6aa26a42,
        64'h69e27902_74a27442,
        64'h70e20004_bc232501,
        64'ha81ff0ef_85264581,
        64'hbf35c55c_4bdc611c,
        64'ha0e1dd5d_2501df9f,
        64'hf0ef8526_45810cd6,
        64'h0a63fff6_46030006,
        64'hc68300f5_86330785,
        64'h00f706b3_708cef89,
        64'h8ba100b7_47831207,
        64'h80630007_47836c98,
        64'h10051163_2501ce0f,
        64'hf0ef6088_48cc492d,
        64'h10051963_2501adff,
        64'hf0ef8526_458100f9,
        64'h05a30200_0793943a,
        64'h09479b63_470d1d37,
        64'h89630024_478300f9,
        64'h00a302e0_07930b37,
        64'h94630014_47830139,
        64'h00230d37_96630004,
        64'h4783b42f_f0ef854a,
        64'h02000593_462d0204,
        64'hb9030d57_84630d47,
        64'h86630004_47834b21,
        64'h02e00993_05c00a93,
        64'h02f00a13_0ce7f063,
        64'h47fd0004_47030004,
        64'ha6230405_0ce79463,
        64'h05c00713_00e78663,
        64'h842e84aa_02f00713,
        64'h0005c783_e05ae456,
        64'he852ec4e_f04afc06,
        64'hf426f822_7139b7e9,
        64'hdb1c2785_5b1c2a85,
        64'h6018f141_2501d24f,
        64'hf0ef0145_0223b7b9,
        64'hc848a89f_f0ef85a6,
        64'hc8046008_d91c4157,
        64'h87bb591c_00faed63,
        64'h00254783_60084a05,
        64'h02aa2823_aabff0ef,
        64'h855285a6_00043a03,
        64'hbf0ff0ef_03450513,
        64'h45812000_06136008,
        64'hf5792501_de0ff0ef,
        64'h6008fcf4_8de357fd,
        64'hfcf48be3_4785d4bd,
        64'h451d0005_049be83f,
        64'hf0ef480c_f60a0ee3,
        64'h06f4e063_4d1c6008,
        64'hb7614505_00f49463,
        64'h57fdbf49_45090097,
        64'he4634785_0005049b,
        64'hb2fff0ef_fc0a9fe3,
        64'h0157fab3_37fd0049,
        64'h5a9b0025_4783bf5d,
        64'h4501ec1c_97ce0347,
        64'h87930124_15230996,
        64'h601cfcf7_75e30009,
        64'h071b0085_5783e18d,
        64'hc85c6108_2785480c,
        64'h00099d63_842a8a2e,
        64'h00f97993_d7ed495c,
        64'h80826121_6aa26a42,
        64'h69e27902_74a27442,
        64'h70e24511_eb9993c1,
        64'he456e852_ec4ef426,
        64'h03091793_2905f822,
        64'hfc0600a5_5903f04a,
        64'h7139b795_547df6f5,
        64'h14e34785_dd612501,
        64'hdbdff0ef_852685ce,
        64'h8622bfb5_00f482a3,
        64'h0017e793_0054c783,
        64'hc89c37fd_f8e788e3,
        64'h577dc4c0_489c0209,
        64'h9063e905_2501debf,
        64'hf0ef8526_85a2167d,
        64'h10000637_b7cdfd24,
        64'h1de3fb45_0ae30555,
        64'h0a63c901_2501c0df,
        64'hf0ef8526_85a24409,
        64'hb7e94401_012a6463,
        64'h00f46763_24054c9c,
        64'h5afd4a05_844afef4,
        64'h61e3894e_4c9c08f4,
        64'h026357fd_80826121,
        64'h6aa26a42_69e27902,
        64'h74a27442_70e28522,
        64'h44050087_ed634785,
        64'h0005041b_c5bff0ef,
        64'ha8154905_02f96d63,
        64'h4d1c0009_056300c5,
        64'h2903e991_89ae84aa,
        64'he456e852_f04af822,
        64'hfc06ec4e_f4267139,
        64'hbf79012a_81a300fa,
        64'h81230189_591b0109,
        64'h579b00fa_80a30087,
        64'hd79b0324_0a230107,
        64'hd79b9426_0109179b,
        64'h29010125_69338d71,
        64'hf0000637_2501d96f,
        64'hf0ef8556_9aa60344,
        64'h0a931fc4_74130024,
        64'h141bf80a_16e30005,
        64'h0a1bfdcf_f0ef9dbd,
        64'h0075d59b_515cbf79,
        64'h01348223_03240aa3,
        64'h0089591b_0109591b,
        64'h0109191b_03240a23,
        64'h94261fe4_74130014,
        64'h141bfc0a_12e30005,
        64'h0a1b815f_f0ef9dbd,
        64'h0085d59b_515cb7e9,
        64'h0127e933_9bc100f9,
        64'h79130089_591b0347,
        64'hc7830154_87b38082,
        64'h61216aa2_6a4269e2,
        64'h790274a2_85527442,
        64'h70e200f4_82234785,
        64'h032a8a23_9aa60ff9,
        64'h79130049_591bc40d,
        64'h1ffafa93_000a1f63,
        64'h00050a1b_86fff0ef,
        64'h9dbd8526_009ad59b,
        64'h50dc00f4_82234785,
        64'h02f98a23_99a60ff7,
        64'hf7938fd9_8ff50049,
        64'h179b00f7_f71316c1,
        64'h66850347_c7830134,
        64'h87b3cc19_1ff9f993,
        64'h0ff97793_00198a9b,
        64'h8805060a_16630005,
        64'h0a1b8bdf_f0ef9dbd,
        64'h0099d59b_00b989bb,
        64'h515c0015_d99b0937,
        64'h94630ee7_8863470d,
        64'h0ae78f63_842e8932,
        64'h47090005_47830af5,
        64'hf0634a09_84aa4d1c,
        64'h0ab9f563_4a094985,
        64'he456f04a_f426f822,
        64'hfc06e852_ec4e7139,
        64'h80826105_64a28526,
        64'h644260e2_00e78223,
        64'h4705601c_00e78023,
        64'h57156c1c_f3cff0ef,
        64'h45810200_06136c08,
        64'hec990005_049b939f,
        64'hf0ef6008_484ce495,
        64'h0005049b_f35ff0ef,
        64'h842aec06_e426e822,
        64'h110100a5_5583b795,
        64'h4505bfc1_4134043b,
        64'hf6f4f7e3_4f9c0009,
        64'h3783f69a_fce30144,
        64'h8c630005_049be75f,
        64'hf0efbf7d_2501e5df,
        64'hf0ef0134_766385a6,
        64'h00093503_09924a85,
        64'h5a7d0027_c98384ba,
        64'hb75d4501_00893c23,
        64'h943e0347_87930416,
        64'h883d0009_378300f9,
        64'h2a239fa9_0044579b,
        64'hd1710099_28235788,
        64'hfce477e3_0087d703,
        64'heb0d5798_00e69463,
        64'h470d0007_c683e0a9,
        64'h842efee4_f4e34f98,
        64'h611c8082_61216aa2,
        64'h6a4269e2_790274a2,
        64'h744270e2_450900f4,
        64'h9c63892a_478500b5,
        64'h1523e456_e852ec4e,
        64'hf822fc06_f04a4544,
        64'hf4267139_8082853e,
        64'h4785bfb9_02455793,
        64'h1512ffaf_f0ef954a,
        64'h03450513_1fc57513,
        64'h0024151b_f93d2501,
        64'ha3bff0ef_9dbd0075,
        64'hd59b515c_b7618fc9,
        64'h0087979b_03494503,
        64'h03594783_99221fe4,
        64'h74130014_141bf145,
        64'h2501a65f_f0ef9dbd,
        64'h0085d59b_515cbf4d,
        64'h93d117d2_bf658391,
        64'hc0198fc5_0087979b,
        64'h88050349_4783994e,
        64'h1ff9f993_f5792501,
        64'ha93ff0ef_0344c483,
        64'h854a9dbd_94ca1ff4,
        64'hf4930099_d59b0014,
        64'h899b0249_27838082,
        64'h6145853e_69a26942,
        64'h64e27402_70a257fd,
        64'hc9112501_ac7ff0ef,
        64'h9dbd0094_d59b9cad,
        64'h515c0015_d49b00f7,
        64'h1e6308d7_0d63468d,
        64'h06d70b63_842e4689,
        64'h00054703_02e5f963,
        64'h892ae44e_ec26f022,
        64'hf406e84a_71794d18,
        64'h0eb7f563_47858082,
        64'h45018082_9d3d02b7,
        64'h87bb5548_00254783,
        64'h00e7f963_377985be,
        64'hffe5879b_4d188082,
        64'h610564a2_644260e2,
        64'h00a03533_25016710,
        64'h50ef4581_46010014,
        64'h45030004_02a367d0,
        64'h50ef85a6_4685d810,
        64'h22f401a3_22e40123,
        64'h20d40ca3_20d40c23,
        64'h0187d79b_0107d71b,
        64'h260522e4_00a322f4,
        64'h00230720_06930014,
        64'h45030087_571b0107,
        64'h571b0107_971b5010,
        64'h20e40f23_445c20f4,
        64'h0fa30187_d79b0107,
        64'hd71b20e4_0ea320f4,
        64'h0e230087_571b0107,
        64'h571b0107_971b20e4,
        64'h0d2302e4_0ba30410,
        64'h0713481c_20f40da3,
        64'h02f40b23_06100793,
        64'h02f40aa3_02f40a23,
        64'h05200793_22f409a3,
        64'hfaa00793_22f40923,
        64'h05500793_9fdff0ef,
        64'h85264581_20000613,
        64'h03440493_0af71b63,
        64'h47850054_47030cf7,
        64'h1063478d_00044703,
        64'hed692501_c01ff0ef,
        64'h842ae426_ec06e822,
        64'h1101bdcd_9cbd0017,
        64'hd79b8885_029787bb,
        64'h478db709_0014949b,
        64'h00f91563_4789d41c,
        64'h9fb5e00a_84e3b545,
        64'ha19ff0ef_05440513,
        64'hb5b10005_099ba27f,
        64'hf0ef0584_0513b351,
        64'h47810004_2a230124,
        64'h002300f4_132362f7,
        64'h10230000_971793c1,
        64'h17c22785_62e7d783,
        64'h00009797_c448a57f,
        64'hf0ef2204_0513c808,
        64'ha61ff0ef_21c40513,
        64'h00f51c63_27278793,
        64'h25016141_77b7a77f,
        64'hf0ef2184_051302f5,
        64'h17632527_87932501,
        64'h416157b7_a8dff0ef,
        64'h03440513_04e79263,
        64'ha5570713_4107d79b,
        64'h776d0107_979b8fd9,
        64'h0087979b_000402a3,
        64'h23244703_23344783,
        64'he13d2501_ce7ff0ef,
        64'h8522001a_059b06e7,
        64'h9b634705_4107d79b,
        64'h0107979b_8fd90087,
        64'h979b0644_47030654,
        64'h478308f9_1963478d,
        64'h00f402a3_f8000793,
        64'hc45cc81c_57fdee99,
        64'he6e30094_d49b1ff4,
        64'h849b0024_949bd408,
        64'hb09ff0ef_06040513,
        64'hf00a93e3_10e91163,
        64'h470dd05c_03442023,
        64'hcc04d458_014787bb,
        64'h24890147_073b0909,
        64'h00b93933_19556941,
        64'h00b67763_49051655,
        64'h6605f326_6ce384ae,
        64'h032655bb_40c5063b,
        64'hf4c563e3_873200d7,
        64'h063b9f3d_004ad71b,
        64'h27810334_86bbdfa9,
        64'h8fd90087_979b2501,
        64'h04244703_04344783,
        64'h14050e63_8d5d0085,
        64'h151b0474_47830484,
        64'h4503ffbd_00faf793,
        64'h01541423_00faeab3,
        64'h008a9a9b_04544783,
        64'h04644a83_ffc100f9,
        64'h77b3fff9_079b2901,
        64'hfa0903e3_01240123,
        64'h04144903_faf769e3,
        64'h0ff7f793_009401a3,
        64'hfff4879b_47050134,
        64'h2e230444_44832981,
        64'h1a098763_00f9e9b3,
        64'h0089999b_04a44783,
        64'h04b44983_fee791e3,
        64'h20000713_4107d79b,
        64'h0107979b_8fd90087,
        64'h979b03f4_47030404,
        64'h4783b785_47b5c119,
        64'h4a01f6e5_05e34785,
        64'h470dbf85_00e51963,
        64'h4785470d_fe9915e3,
        64'h0491c10d_ea1ff0ef,
        64'h852285d2_000a0763,
        64'h45090004_aa030104,
        64'h8913ff2a_14e30991,
        64'h094100a9_a0232501,
        64'hc51ff0ef_854ac789,
        64'h4501ffc9_478389a6,
        64'h23a40a13_1fa40913,
        64'h848a04f5_1a634785,
        64'hee5ff0ef_85224581,
        64'hf5718911_00090463,
        64'hfb79478d_00157713,
        64'h136060ef_00a400a3,
        64'h00040023_0ff4f513,
        64'h80826161_853e6ae2,
        64'h7a0279a2_794274e2,
        64'h640660a6_47a9c111,
        64'h89110009_0563e385,
        64'h00157793_222060ef,
        64'h00144503_c79d0004,
        64'h47830089_b023c015,
        64'h47b184aa_638097ba,
        64'h8a878793_0000a797,
        64'h00351713_02054e63,
        64'h47adddbf_f0ef8932,
        64'h852e89aa_00053023,
        64'hec56f052_fc26e0a2,
        64'he486f44e_f84a715d,
        64'hbfcd450d_80826105,
        64'h690264a2_644260e2,
        64'h00a03533_8d050125,
        64'h75332501_d25ff0ef,
        64'h08640513_00978c63,
        64'h45010127_f7b31465,
        64'h04930054_4537fff5,
        64'h09130100_05370005,
        64'h079bd4bf_f0ef06a4,
        64'h051302e7_9f63a557,
        64'h07134107_d79b776d,
        64'h0107979b_8fd90087,
        64'h979b4509_23244703,
        64'h23344783_e52d2501,
        64'hfa3ff0ef_842ad91c,
        64'h00050223_57fde04a,
        64'he426ec06_e8221101,
        64'h80826105_690264a2,
        64'h644260e2_85220324,
        64'ha823597d_4405c119,
        64'h25012d60_60ef0344,
        64'h8593864a_46850014,
        64'hc503ec19_0005041b,
        64'hfddff0ef_892e84aa,
        64'h02b78763_4401e04a,
        64'he426ec06_e8221101,
        64'h591c8082_4501f8df,
        64'hf06fc399_00454783,
        64'hb7f94505_b7e5397d,
        64'h34e060ef_85ce8626,
        64'h9cbd4685_00144503,
        64'h4c5cff2a_74e34a05,
        64'h00344903_80826145,
        64'h6a0269a2_694264e2,
        64'h740270a2_450100e7,
        64'heb6340f4_87bb0004,
        64'h02234c58_505ce131,
        64'h25013900_60ef85ce,
        64'h86264685_00154503,
        64'h842a0345_0993e052,
        64'he84af406_5904e44e,
        64'hec26f022_71798082,
        64'h853e2781_8fd50107,
        64'h979b8fd1_0087179b,
        64'h0145c603_0155c703,
        64'h00e51d63_0006879b,
        64'h8edd0087_979b470d,
        64'h01a5c683_01b5c783,
        64'h80824525_80820141,
        64'h60a24525_c3914501,
        64'h00157793_402060ef,
        64'h0017c503_e4061141,
        64'h02e69063_00855703,
        64'h0067d683_c70d0007,
        64'hc703cb85_611cc915,
        64'hbfd5aa27_47030000,
        64'ha7178082_853ae11c,
        64'h0006871b_078900b6,
        64'h66630ff6_f593fd06,
        64'h869b577d_46050007,
        64'hc683b7dd_0705a00d,
        64'h577d00d7_06630017,
        64'h869300c6_986302d5,
        64'hfc630007_468303a0,
        64'h06130200_0593cf99,
        64'h873e611c_80826105,
        64'h690264a2_644260e2,
        64'h00040023_00f49323,
        64'h8fd90087_979b0169,
        64'h47030179_478300f4,
        64'h92238fd9_0087979b,
        64'h01894703_01994783,
        64'hc088f4bf_f0ef00f5,
        64'h842384ae_01c90513,
        64'h00b94783_fcd79be3,
        64'h07850405_00e40023,
        64'h04050114_00230103,
        64'h15630007_831b0e50,
        64'h071300a7_146302c7,
        64'h00630007_470300f9,
        64'h073346ad_02e00893,
        64'h48214515_02000613,
        64'h47810185_3903cfb5,
        64'h00958413_e04ae426,
        64'hec06e822_1101495c,
        64'hbfc5feb5_0fa30505,
        64'h808200f6_13630005,
        64'h079b9e29_b7d500d7,
        64'h00230785_00f50733,
        64'h00074683_00f58733,
        64'h808200e6_13630007,
        64'h871b4781_80822501,
        64'h8d5d0562_8fd907c2,
        64'h00354503_00254783,
        64'h8f5d07a2_00054703,
        64'h00154783_b7d914fd,
        64'hb7e9bf9f_f0efbfc1,
        64'h710a8493_7c9050ef,
        64'h4501dff1_54fd000a,
        64'h2783bfc5_c13ff0ef,
        64'hfc075de3_03379713,
        64'h83093783_02074563,
        64'h03379713_83093783,
        64'h5a0b0493_f23fe0ef,
        64'h8522e78d_0009a783,
        64'he4a9be07_a5230000,
        64'ha797be07_ab230000,
        64'ha797c007_a1230000,
        64'ha797be07_ad230000,
        64'ha797c007_93230000,
        64'ha797c2f7_07a30000,
        64'ha7170054_4783c2f7,
        64'h0d230000_a7170044,
        64'h4783c4f7_02a30000,
        64'ha7170034_4783c4f7,
        64'h08230000_a7173000,
        64'h19370026_2b370024,
        64'h4783c6f7_01a30000,
        64'ha7176a89_c54a0a13,
        64'h0000aa17_00144783,
        64'hc6f70c23_0000a717,
        64'hc6098993_0000a997,
        64'h44810004_4783c864,
        64'h04130000_a41709b0,
        64'h30efeb25_05130000,
        64'h9517c9a5_c5830000,
        64'ha597ca36_46030000,
        64'ha617cac6_c6830000,
        64'ha697cb78_48030000,
        64'ha817cbe7_c7830000,
        64'ha797cc57_47030000,
        64'ha7170d70_30efede5,
        64'h05130000_951780e7,
        64'hb423e05a_e456e852,
        64'hec4ef04a_f426f822,
        64'hfc068f4d_91c115c2,
        64'h00800737_71398087,
        64'hb5838007_b6033000,
        64'h17b78082_61616ae2,
        64'h7a0279a2_794274e2,
        64'h82f6b423_47a16406,
        64'h60a68086_b7838006,
        64'hb78380f6_b42393c1,
        64'h80a6b023_17c29101,
        64'h300016b7_8fd91502,
        64'h0ff77713_8ff18321,
        64'h0087179b_f0060613,
        64'h01000637_4722f43f,
        64'hf0ef4512_7ce050ef,
        64'h0028d5a5_85930000,
        64'ha5974609_7de050ef,
        64'h0048d6c5_85930000,
        64'ha5974611_fc941ee3,
        64'h185030ef_00c78023,
        64'h0ff67613_00ca5633,
        64'h0286061b_0405854a,
        64'h0004059b_013407b3,
        64'h028a863b_4499f969,
        64'h09130000_9917da69,
        64'h89930000_a9975ae1,
        64'h44011bf0_30eff9e5,
        64'h05130000_95178a2a,
        64'h047070ef_c63eec56,
        64'hf052f44e_f84afc26,
        64'he0a2e486_04b00513,
        64'h45854601_00740207,
        64'h879b0700_07b7715d,
        64'h80822501_8d5d8d79,
        64'h00ff0737_0085151b,
        64'h8fd98f75_0085571b,
        64'hf0068693_8fd966c1,
        64'h0185579b_0185171b,
        64'h80829141_15428d5d,
        64'h05220085_579b8082,
        64'h614564e2_740270a2,
        64'h85228e0f_f0efe2e5,
        64'h05130000_a5170450,
        64'h0693e267_57030000,
        64'ha717e228_88930000,
        64'ha89785a6_862247b2,
        64'h0007a803_e3c78793,
        64'h0000a797_0d7050ef,
        64'hf4060068_e8458593,
        64'h0000a597_461184ae,
        64'h8432ec26_f0227179,
        64'hbfc14785_ec3ff0ef,
        64'h80826105_64a26442,
        64'h60e2c3c0_0c2007b7,
        64'h29d030ef_06450513,
        64'h00009517_e7990206,
        64'hc1630337_16938304,
        64'hb7033000_14b74781,
        64'h2401ec06_e42643c0,
        64'he8220c20_07b71101,
        64'h80826101_01135f81,
        64'h34838526_60013403,
        64'h60813083_8287b823,
        64'h300017b7_0405a9bf,
        64'hf0ef8626_fef845e3,
        64'h0006881b_ff063c23,
        64'h06210685_00083803,
        64'h983a0036_98139742,
        64'h85b24681_4037d79b,
        64'h30000837_860a2785,
        64'h0077e793_37ed02d5,
        64'h1e638066_86936685,
        64'hc6918005_069b0001,
        64'h550300d1_00230086,
        64'hd69b0106_d69b0106,
        64'h969b00d1_00a345d4,
        64'h95ba070e_9f318006,
        64'h871b7007_76130084,
        64'h171beb3d_4318f4e7,
        64'h07130000_a717c349,
        64'h27018f71_fff74713,
        64'h00c5163b_10100513,
        64'h8a1d0905_6c63ffc7,
        64'h849b5f20_0513fee7,
        64'h881b2781_60113423,
        64'h5e913c23_639c97ae,
        64'h300005b7_9fad8406,
        64'h879b0387_f5930034,
        64'h179b6685_8387b703,
        64'h00f67413_26016081,
        64'h30239f01_01138307,
        64'hb6033000_17b7bba5,
        64'h46013cf0_30ef17e5,
        64'h05130000_951785aa,
        64'hb36900f4_16236080,
        64'h079300f4_1f230024,
        64'hd78300f4_1e230004,
        64'hd78302f4_142301e4,
        64'h578302f4_132302a0,
        64'h061301c4_57832790,
        64'h50ef8522_85ca4619,
        64'h283050ef_00640513,
        64'h01858593_0000a597,
        64'h46192950_50ef854e,
        64'h02858593_0000a597,
        64'h46192a50_50ef854a,
        64'h85ce4619_00f59a23,
        64'h01658993_02058913,
        64'h20000793_eaf719e3,
        64'h06a7d783_0000a797,
        64'h0285d703_ecf711e3,
        64'h07848493_0000a497,
        64'h0807d783_0000a797,
        64'h0265d703_b1e91f65,
        64'h05130000_9517b9d1,
        64'h1e850513_00009517,
        64'hb9f91c25_05130000,
        64'h9517b1e5_1ac50513,
        64'h00009517_b9cd19e5,
        64'h05130000_9517b9f5,
        64'h18050513_00009517,
        64'hb31917a5_05130000,
        64'h9517bb01_16450513,
        64'h00009517_bb291565,
        64'h05130000_9517b315,
        64'h14050513_00009517,
        64'hb33d13a5_05130000,
        64'h9517b799_357050ef,
        64'h08681025_85930000,
        64'ha5974611_f4f70de3,
        64'h02045703_f6f701e3,
        64'h17fd67c1_01e45703,
        64'hf6e787e3_5fe00713,
        64'hbf95cb4f_f0ef02a4,
        64'h051385ca_521030ef,
        64'h16050513_00009517,
        64'hccaff0ef_852285a6,
        64'h535030ef_16450513,
        64'h00009517_02e79863,
        64'h4d200713_b765d73f,
        64'he0ef02a4_05131465,
        64'h85930000_a5971426,
        64'h06130000_a6171466,
        64'h86930000_a697f7e9,
        64'h439c1527_87930000,
        64'ha797c799_439c1627,
        64'h87930000_a79714f7,
        64'h2f230000_a71747e2,
        64'h04e69463_04300713,
        64'h80826161_79a27942,
        64'h74e26406_60a654e0,
        64'h60ef4501_02a40593,
        64'hff89061b_17478793,
        64'h0000a797_66a24762,
        64'h42b050ef_e43618f7,
        64'h2f230000_a71719e5,
        64'h05130000_a5171965,
        64'h85930000_a5974619,
        64'h47e21ad7_9f230000,
        64'ha79704e7_9b6301c1,
        64'h56830450_071300e1,
        64'h0e230234_470300e1,
        64'h0ea301c1_19030224,
        64'h470300e1_0e232781,
        64'h02744703_00e10ea3,
        64'h01c11783_00f10e23,
        64'h02544783_00f10ea3,
        64'h02644703_02444783,
        64'hbdbd24a5_05130000,
        64'h9517b561_23c50513,
        64'h00009517_bd4922e5,
        64'h05130000_9517a06d,
        64'hdcdfe0ef_450185a2,
        64'h862602a4_122300a1,
        64'h1e238d5d_05220085,
        64'h579bdb3f_f0ef00f4,
        64'h1e230029_d78300f4,
        64'h1d230009_d78302f4,
        64'h10230224_0513fde4,
        64'h859b01c4_578300f4,
        64'h1f230204_12230204,
        64'h012301a4_57835090,
        64'h50ef854a_29c58593,
        64'h0000a597_46195190,
        64'h50ef8522_85ca4619,
        64'h10f71b63_2ce7d783,
        64'h0000a797_02045703,
        64'h12f71363_2dc98993,
        64'h0000a997_2e47d783,
        64'h0000a797_01e45703,
        64'hb73d42a5_05130000,
        64'h9517f0f5_9ce30880,
        64'h079326f5_88630ff0,
        64'h079326f5_87630890,
        64'h0793b73d_f4f58ae3,
        64'h42050513_00009517,
        64'h06c00793_26f58a63,
        64'h06700793_00b7ef63,
        64'h28f58563_08400793,
        64'hbf91f6f5_8de340e5,
        64'h05130000_951705e0,
        64'h079328f5_836305c0,
        64'h0793b7bd_f8f58ae3,
        64'h3f850513_00009517,
        64'h03200793_28f58663,
        64'h02f00793_00b7ef63,
        64'h2af58163_03300793,
        64'h04b7e263_2cf58163,
        64'h06200793_b7c93f65,
        64'h05130000_9517faf5,
        64'h96e30290_07932af5,
        64'h85630210_0793bf6d,
        64'hfef580e3_3dc50513,
        64'h00009517_47d916f5,
        64'h896347c5_00b7ed63,
        64'h2cf58163_47f5a429,
        64'h7ad030ef_fef591e3,
        64'h3c050513_00009517,
        64'h47a118f5_81634799,
        64'ha4157c70_30ef5565,
        64'h05130000_951702f5,
        64'h83633ba5_05130000,
        64'h95174789_10f58463,
        64'h478502b7_e3631af5,
        64'h82634791_04b7e563,
        64'h1cf58163_47b108b7,
        64'he76332f5_886302e0,
        64'h07930174_45836790,
        64'h50ef3d25_05130000,
        64'ha5174619_85ca0064,
        64'h091368d0_50ef4611,
        64'h082884b2_05e94407,
        64'h99638005_079b0af5,
        64'h0e636dd7_879367a1,
        64'h3cf50463_842e8067,
        64'h8793f44e_f84afc26,
        64'he486e0a2_6785715d,
        64'hbf45943e_93c117c2,
        64'h00f11723_8fd90087,
        64'h979b0087_d71b0489,
        64'h00c15783_6df050ef,
        64'h00684609_85a68082,
        64'h61459141_694264e2,
        64'h1542fff5_45137402,
        64'h70a29522_01045513,
        64'h942a9041_14420104,
        64'h551302f0_44634099,
        64'h07bb00a5_893b4401,
        64'h84aaf406_e84aec26,
        64'hf0227179_80824365,
        64'h05130000_9517bf75,
        64'h48050513_00009517,
        64'h84078793_fce608e3,
        64'h48050513_00009517,
        64'h83878713_bfe946e5,
        64'h05130000_95178287,
        64'h879300c7_4963fee6,
        64'h09e34925_05130000,
        64'h95178307_87138082,
        64'hfaf612e3_47450513,
        64'h00009517_81878793,
        64'h00e60a63_47450513,
        64'h00009517_81078713,
        64'h80820141_4d450513,
        64'h0000a517_60a210e0,
        64'h40efe406_4e450513,
        64'h0000a517_51458593,
        64'h00009597_9e3d1141,
        64'h7c07879b_77fd04c7,
        64'hc9635225_05130000,
        64'h951787f7_87936785,
        64'hc3ad4a25_05130000,
        64'h95178006_079b04c7,
        64'h496306e6_0b634c65,
        64'h05130000_95178087,
        64'h871308a7_4463862a,
        64'h0ce50763_82078713,
        64'h67858082_953e057e,
        64'h450597aa_20000537,
        64'he3089536_00178693,
        64'h00756513_157d631c,
        64'h58070713_0000a717,
        64'h80824000_05378082,
        64'h057e4505_bfb12405,
        64'h7ed050ef_854a4581,
        64'h86261d60_40ef855e,
        64'h85ca993e_86268c9d,
        64'h79020097_ff6377a2,
        64'h74c29982_85260009,
        64'h061b45c2_1f8040ef,
        64'h856a86ca_85a66642,
        64'h8082612d_6d0a6caa,
        64'h6c4a6bea_7b0a7aaa,
        64'h7a4a79ea_690e64ae,
        64'h644e60ee_55752220,
        64'h40ef51a5_05130000,
        64'h951785a6_0397e863,
        64'h018487b3_74820409,
        64'h08637922_240040ef,
        64'h855a85a2_cfbd77c2,
        64'h09579263_47a29982,
        64'h9dbd0028_03800613,
        64'h7786028a_05bba091,
        64'h656600f4_64630781,
        64'h578357ad_0d130000,
        64'h9d170800_0cb78000,
        64'h0c375a2b_8b930000,
        64'h9b9756ab_0b130000,
        64'h9b174a85_03800a13,
        64'h440106e7_9d635579,
        64'h83e107e2_631848e7,
        64'h07130000_a7176786,
        64'h9982e16a_e566e962,
        64'hed5ef15a_f556f952,
        64'he1cae5a6_e9a2ed86,
        64'h00884581_89aa0400,
        64'h0613fd4e_7115bfd5,
        64'h8f8d2505_8082e21c,
        64'h00b7f463_45019181,
        64'h87aa1582_b70d0705,
        64'h27850117_00230006,
        64'h54634186_561b0186,
        64'h161bc519_09757513,
        64'h00054503_00cc0533,
        64'h00074603_bfdd4781,
        64'hbf253cfd_fe97eae3,
        64'h27856782_0e4070ef,
        64'he03e855e_b76500c5,
        64'h80230ff6_761395be,
        64'h082c0007_4603bf6d,
        64'h00c59023_95aa9241,
        64'h16420828_00179593,
        64'h00075603_011d1d63,
        64'hbfd1e190_95aa0828,
        64'h00379593_6310010d,
        64'h1963bf9d_46914821,
        64'h07859752_488967a2,
        64'h67023760_40efe03a,
        64'he43e855a_85d69201,
        64'h1602c190_95aa2601,
        64'h08280027_95934310,
        64'h02dd1963_b79d557d,
        64'hd13d0b80_70ef9936,
        64'h92811682_41b4043b,
        64'h66823ae0_40effa07,
        64'h8c23e036_69450513,
        64'h00009517_97ba1098,
        64'h0b079c63_0006881b,
        64'h02e00893_85ba4781,
        64'h083803bd_06bb0d9d,
        64'he56399be_034787b3,
        64'h9381020d_979305b6,
        64'h6b630007_861b4889,
        64'h48214691_4781874e,
        64'h000c8d9b_008cf463,
        64'h00040d9b_408040ef,
        64'h6d850513_00009517,
        64'h85ca8082_61697da6,
        64'h7d467ce6_6c0a6baa,
        64'h6b4a6aea_7a0a79aa,
        64'h794a74ea_640e60ae,
        64'h4501e00d_5dcc0c13,
        64'h00008c17_684b8b93,
        64'h00009b97_71cb0b13,
        64'h00009b17_020a5a13,
        64'h001a849b_020d1a13,
        64'h001d1a9b_03acdcbb,
        64'h4cc1000c_956302cc,
        64'hdcbb0400_0c9300e7,
        64'hf6638436_8d3289ae,
        64'h892a0400_0793f4ee,
        64'he162e55e_e95aed56,
        64'hf152fd26_e586f8ea,
        64'hf54ef94a_e1a202c7,
        64'h073b8cba_fce67155,
        64'h4a40406f_610576e5,
        64'h05130000_951764a2,
        64'h690285a6_864a60e2,
        64'h64424be0_40ef7665,
        64'h05130000_951785a2,
        64'hc8014ce0_40ef8932,
        64'h77050513_00009517,
        64'h85be0785_14590087,
        64'h74630104_5433942a,
        64'h472500d4_14334405,
        64'h03b6869b_02e50533,
        64'h4729c10d_44018d79,
        64'hfff74713_01071733,
        64'h577db7f5_7c450513,
        64'h00009517_85aafab7,
        64'h1ce32705_5200406f,
        64'h61057da5_05130000,
        64'h951785aa_690264a2,
        64'h60e26442_e495e04a,
        64'he822ec06_00074483,
        64'he426972e_11017765,
        64'h85930000_a5979301,
        64'h1702cf85_00f557b3,
        64'h883e03c6_879b02e8,
        64'h86bb4599_58d94701,
        64'h862ebfa1_7fc50513,
        64'h00009517_85aabf55,
        64'h4401bf51_843a0086,
        64'hf46302f4_5733bf61,
        64'h02e45433_5900406f,
        64'h61058425_05130000,
        64'ha5176902_64a285ca,
        64'h862660e2_64425aa0,
        64'h40ef8525_05130000,
        64'ha51785a2_c8015ba0,
        64'h40ef84b2_85c50513,
        64'h0000a517_943e0014,
        64'h44130324_341302e4,
        64'h743302f4_57b30640,
        64'h07130087_7d630630,
        64'h0713cf39_02f47733,
        64'h46a547a9_0687e263,
        64'h47293e80_0793c815,
        64'h02f555b3_02f57433,
        64'hbf7d2407_87934685,
        64'hb7d9a007_87934681,
        64'h6140406f_61058a65,
        64'h05130000_a51785aa,
        64'h690264a2_60e26442,
        64'h02091663_e426e822,
        64'hec060007_4903e04a,
        64'h97361101_87470713,
        64'h0000b717_3e800793,
        64'h46890ca7_fc633e70,
        64'h079304a7_676323f7,
        64'h8713000f_47b704a7,
        64'h6963862e_9ff78713,
        64'h3b9ad7b7_8082612d,
        64'h450160ee_678040ef,
        64'h90050513_0000a517,
        64'h002cfebf_f0efed86,
        64'h45050c80_0613002c,
        64'h7115f73f_f06f4581,
        64'h862e86b2_80826145,
        64'h69a26942_64e2854a,
        64'h740270a2_26a060ef,
        64'h91858593_0000a597,
        64'h00890533_ffd4841b,
        64'h00f44463_ffe4879b,
        64'h9c2968e0_40ef954a,
        64'h94860613_0000a617,
        64'h86ce40a4_85bb0095,
        64'h5d630009_8f63842a,
        64'h6ac040ef_854a85a6,
        64'h96060613_0000a617,
        64'he1870713_00009717,
        64'h96868693_0000a697,
        64'hc5091ba6_86930000,
        64'ha6978932_89ae84b6,
        64'hf022f406_e44ee84a,
        64'hec267179_bfdd72a0,
        64'h40ef8562_b7f10905,
        64'h734040ef_856600fb,
        64'he7630ff7_f793fe05,
        64'h879b0007_c5830129,
        64'h87b3bf15_04857520,
        64'h40ef5325_05130000,
        64'ha51700f4_5a630009,
        64'h079b4124_093b76a0,
        64'h40ef00f4_f913855a,
        64'hff2dcce3_2d8577a0,
        64'h40ef8552_bfdd7820,
        64'h40ef8562_b75d0905,
        64'h78c040ef_856600fb,
        64'he7630ff7_f793fe05,
        64'h879b0007_c5830129,
        64'h87b3a805_00f97913,
        64'h4d81fffd_4913068d,
        64'h12637b60_40efa165,
        64'h05130000_a5170007,
        64'hc5830099_87b37ca0,
        64'h40ef8552_7d0040ef,
        64'h5b050513_0000a517,
        64'h02879d63_0009079b,
        64'hff048913_7e8040ef,
        64'h855ae39d_00f47793,
        64'hc01d8082_61656da2,
        64'h6d426ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h694664e6_740670a6,
        64'h03544163_0004841b,
        64'hfff58d1b_a6cc8c93,
        64'h0000ac97_a7cc0c13,
        64'h0000ac17_06000b93,
        64'ha70b0b13_0000ab17,
        64'h740a0a13_0000aa17,
        64'h44818aae_89aae46e,
        64'he8caf0a2_f486e86a,
        64'hec66f062_f45ef85a,
        64'hfc56e0d2_e4ceeca6,
        64'h7159b7cd_069040ef,
        64'hc007a823_0000b797,
        64'ha9850513_0000a517,
        64'h80826151_641260b2,
        64'h85220870_40efa7e5,
        64'h05130000_a517a565,
        64'h85930000_a597860a,
        64'hc10d842a_e01ff0ef,
        64'h85220a70_40efa765,
        64'h05130000_a517a765,
        64'h85930000_a597842a,
        64'h00054603_00154683,
        64'h00254703_00354783,
        64'h00454803_00554883,
        64'he222e606_716d8082,
        64'h616569a6_694664e6,
        64'h74064501_70a67f01,
        64'h01138ddf_f0ef86c6,
        64'h85a61808_56326882,
        64'hfc4ff0ef_03e10513,
        64'h863e86c2_85a267c2,
        64'h6822f94f_f0efd64e,
        64'h05210513_85a2864a,
        64'h86ba943e_7fc40413,
        64'h6762747d_97ba8107,
        64'h87931018_67857a00,
        64'h60efd602_e83eec3a,
        64'he4428936_89b2e046,
        64'h05a10513_84aa8101,
        64'h0113e4ce_e8caeca6,
        64'hf0a2f486_715915b0,
        64'h406fb125_05130000,
        64'ha51785aa_80826125,
        64'h7aa27a42_79e26906,
        64'h64a66446_450160e6,
        64'h911a6305_96fff0ef,
        64'h85ce86a6_10084652,
        64'h855ff0ef_460156fd,
        64'h02e10513_85a2821f,
        64'hf0ef0440_06130430,
        64'h06930421_051385a2,
        64'h943e1451_978a020a,
        64'h879312f1_1c233537,
        64'h87936799_12f11b23,
        64'h26378793_77e10390,
        64'h60ef04f1_06230661,
        64'h05134641_479985ce,
        64'h04f11523_10100793,
        64'h005060ef_ca3e04a1,
        64'h05134581_0f000613,
        64'h0fc00793_067060ef,
        64'h000107a3_15410223,
        64'h14f101a3_14510513,
        64'h460585ca_57fd0810,
        64'h60ef13f1_05134611,
        64'h95beff04_0593978a,
        64'h020a8793_12f10f23,
        64'h479112f1_0ea30370,
        64'h07930a50_60ef0141,
        64'h07a31a68_460585ca,
        64'h993e978a_020a8793,
        64'h12f11d23_13500793,
        64'hc83e4a05_fef40913,
        64'h439cc827_87930000,
        64'hb7970870_60ef8526,
        64'h55fd4619_94beff84,
        64'h0493978a_020a8793,
        64'h747d27f0_40efca02,
        64'h6a85c225_05130000,
        64'ha517911a_89aaf456,
        64'hf852fc4e_e0cae4a6,
        64'he8a2ec86_711d737d,
        64'hb34d2a70_40efc0e5,
        64'h05130000_a517bf45,
        64'hc0850513_0000a517,
        64'h95be978a_d0040593,
        64'h35078793_67852cb0,
        64'h40efc025_05130000,
        64'ha5172d70_40efbfe5,
        64'h05130000_a51700fa,
        64'h20234785_de0794e3,
        64'h000a2783_b3fd2f30,
        64'h40efc0a5_05130000,
        64'ha517bbf5_301040ef,
        64'hc0050513_0000a517,
        64'h95be978a_f0040593,
        64'h35048793_319040ef,
        64'hc0850513_0000a517,
        64'h95bee004_0593978a,
        64'h35048793_331040ef,
        64'h02f5d5bb_e107879b,
        64'h678502f6_763b02f5,
        64'hf6bb02f5_d63b03c0,
        64'h0793f4f7_1e230000,
        64'hb7170121_5783f6f7,
        64'h13230000_b717c2e5,
        64'h05130000_a51755c2,
        64'h01015783_371040ef,
        64'hc2050513_0000a517,
        64'h01014583_01114603,
        64'h01214683_01314703,
        64'h38d040ef_c1c50513,
        64'h0000a517_01814583,
        64'h01914603_01a14683,
        64'h01b14703_3a9040ef,
        64'h00b14703_fcf71323,
        64'h0000b717_c1c50513,
        64'h0000a517_00814583,
        64'h35215783_fcf71e23,
        64'h0000b717_00914603,
        64'h00a14683_35015783,
        64'h3dd040ef_c1c50513,
        64'h0000a517_35014583,
        64'h35114603_35214683,
        64'h35314703_267060ef,
        64'h01490593_4611953e,
        64'hcb840513_978a3504,
        64'h87936485_27f060ef,
        64'h0e880109_05934611,
        64'h41d040ef_c4c50513,
        64'h0000a517_00fa2023,
        64'h47851207_9a63000a,
        64'h2783b321_d00d0023,
        64'h2ab060ef_9d228562,
        64'h866ab749_cc048513,
        64'hbb39cef4_2023401c,
        64'h00f41023_8fd90087,
        64'h979b0087_d71bce24,
        64'h578300f4_11238fd9,
        64'h0087979b_0087d71b,
        64'hce045783_2e7060ef,
        64'h4611953e_ce048513,
        64'h978a3507_87936785,
        64'hbfdd855a_4611b395,
        64'h303060ef_85564611,
        64'hb3bdf00d_00233110,
        64'h60ef9d22_953e866a,
        64'hf0048513_978a3507,
        64'h87936785_a00d953e,
        64'h978a3507_87936785,
        64'h4611cd04_85138082,
        64'h3b010113_35013d03,
        64'h35813c83_36013c03,
        64'h36813b83_37013b03,
        64'h37813a83_38013a03,
        64'h38813983_39013903,
        64'h39813483_3a013403,
        64'h3a813083_911a6305,
        64'hcf3ff0ef_0e8885de,
        64'h86ca5672_bd9ff0ef,
        64'h35e10513_85a24601,
        64'h56fdba5f_f0ef3721,
        64'h051385a2_04400613,
        64'h04300693_943ecec4,
        64'h0413978a_350a8793,
        64'h46f11423_35378793,
        64'h679946f1_13232637,
        64'h879377e1_3bf060ef,
        64'h36f10e23_39610513,
        64'h85de4799_464136f1,
        64'h1d231010_079338b0,
        64'h60efde3e_37a10513,
        64'h45810f00_06131020,
        64'h07933ed0_60ef4731,
        64'h0d230001_03a346f1,
        64'h0ca347b1_051385a6,
        64'h460557fd_407060ef,
        64'h47410a23_47510513,
        64'h461195be_cf440593,
        64'h978a350a_879346f1,
        64'h09a30360_07934290,
        64'h60ef4741_072346f1,
        64'h05134611_4a1195be,
        64'hcf040593_978a350a,
        64'h879346f1_06a30320,
        64'h079344d0_60efc0d2,
        64'h46c10513_85a64605,
        64'h94becb74_0493c2a6,
        64'h978a350a_879346f1,
        64'h15231350_079300f1,
        64'h03a3478d_429060ef,
        64'h854a55fd_4619993e,
        64'hcf840913_978a350a,
        64'h879361f0_40efde02,
        64'h54e25a52_e3c50513,
        64'h0000a517_49f060ef,
        64'h953e4611_01490593,
        64'hce840513_978a350a,
        64'h87934b50_60ef013c,
        64'ha023953e_46110109,
        64'h0593ce44_05134985,
        64'h978a350a_87936a85,
        64'h16079263_000ca783,
        64'h3af59f63_478938f5,
        64'h83634799_24f58363,
        64'h747d4795_00614583,
        64'hf8e79ce3_0ff00713,
        64'h24e78563_03800713,
        64'haac94605_cb648513,
        64'hfae798e3_03500713,
        64'h20e78e63_03300713,
        64'h00f76e63_22e78163,
        64'h03600713_b769e00d,
        64'h002352d0_60ef9d22,
        64'h953e866a_e0048513,
        64'h978a3507_87936785,
        64'hfee794e3_473d22e7,
        64'h83634731_bf4d6e30,
        64'h40ef0625_05130000,
        64'ha51785be_22e78763,
        64'hcc848513_470d2ae7,
        64'h89634705_02f76263,
        64'h22e78f63_471904f7,
        64'h6b6326e7_8b6301a9,
        64'h89bb0589_02a00713,
        64'h29890f07_c7830015,
        64'hcd030139_07b395ca,
        64'h0f098593_9c3a9b3a,
        64'h49818a36_8cb28bae,
        64'hd0048c13_cb848b13,
        64'h970a3507_87139aba,
        64'hcd848a93_970a3507,
        64'h871374fd_678524f7,
        64'h1d634789_00054703,
        64'ha0017670_40eff5e5,
        64'h05130000_a51785aa,
        64'h00e7ea63_892a5800,
        64'h073797aa_d0040023,
        64'hf0040023_e0040023,
        64'hca040b23_ce042023,
        64'hd00007b7_943e747d,
        64'h978a911a_35078793,
        64'h35a13823_35913c23,
        64'h37813023_37713423,
        64'h37613823_37513c23,
        64'h39413023_39313423,
        64'h38913c23_3a113423,
        64'h39213823_3a813023,
        64'h6785737d_c5010113,
        64'hfadff06f_614564e2,
        64'h00e4859b_70a27402,
        64'h852200f4_162347a1,
        64'h663060ef_85b64619,
        64'h852266a2_66f060ef,
        64'he436f406_46190519,
        64'h84b2842a_ec26f022,
        64'h71798082_01416402,
        64'h60a28522_fa1ff0ef,
        64'he4064501_85aa8622,
        64'h0005841b_e0221141,
        64'hbfe10505_01173023,
        64'h97369742_0008b883,
        64'h00e588b3_00351713,
        64'h808280c6_b82396be,
        64'h678500f7_47630005,
        64'h071b6805_450102e7,
        64'hc7bb2785_0077e793,
        64'hfff6079b_8007bc23,
        64'h97b64721_67856394,
        64'h2b878793_0000b797,
        64'h80826145_740270a2,
        64'h00f41523_fff7c793,
        64'h9fb94107_d71b9fb9,
        64'h93411742_4107579b,
        64'hfed79ce3_9f31ffe7,
        64'hd6030789_470187a2,
        64'h01440693_727060ef,
        64'h01040513_002c4611,
        64'h733060ef_00c40513,
        64'h00041523_006c4611,
        64'h00f404a3_47c57490,
        64'h60efec3e_00840513,
        64'h00041323_082c4621,
        64'h47c175d0_60ef0044,
        64'h05130161_05934609,
        64'h76b060ef_00f11b23,
        64'hc4360509_084c57fd,
        64'h460900f1_1a238fd9,
        64'h0087979b_0ff77713,
        64'h0087d713_c632842a,
        64'h419c00f5_10230457,
        64'h879b6785_c19c27d1,
        64'hf022f406_7179419c,
        64'h80820005_132300f5,
        64'h122300d5_112300c5,
        64'h10238fd9_0087979b,
        64'h0ff77713_c19c0087,
        64'hd7138ed9_06a20086,
        64'hd71b8e59_27a10622,
        64'h0086571b_419cc19c,
        64'h2785c319_0017f713,
        64'h419cbfcd_fda00513,
        64'h80826121_74a27442,
        64'h70e29782_85a66562,
        64'h701ce509_c39ff0ef,
        64'h842a0830_65a2c105,
        64'hc7dff0ef_84b2e42e,
        64'hf822fc06_f4267139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2655c,
        64'h862686ca_6562e519,
        64'hc75ff0ef_083065a2,
        64'hc115cb7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2615c,
        64'h862686ca_6562e519,
        64'hcb5ff0ef_083065a2,
        64'hc115cf7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hb7e16522_f569cdbf,
        64'hf0ef8526_85ce0030,
        64'hbfc90284_8493c501,
        64'h681060ef_854a608c,
        64'h254050ef_855285ca,
        64'h60908082_61216a42,
        64'h69e27902_74a27442,
        64'h70e24501_00849b63,
        64'h942602f4_043325ea,
        64'h0a130000_aa1789ae,
        64'h892afc06_e852ec4e,
        64'hf04a0280_079302f4,
        64'h043b840d_8c0554e4,
        64'h84930000_b4975564,
        64'h04130000_b417f426,
        64'hf822639c_49478793,
        64'h0000b797_7139bfdd,
        64'h45018082_61056442,
        64'h60e2fda0_05138302,
        64'h610560e2_65a26442,
        64'h85220003_0e630205,
        64'h3303c919_db9ff0ef,
        64'he42eec06_4108842a,
        64'he8221101_bfc56562,
        64'hf96dd97f_f0ef0830,
        64'h80826145_70a24501,
        64'he50965a2_de1ff0ef,
        64'hf406e42e_7179bfc1,
        64'h5479fcf7_1be30ff0,
        64'h079300c7_c70367a2,
        64'h0de080ef_6522f565,
        64'h842adcff_f0ef85a6,
        64'h00308522_80826145,
        64'h64e27402_70a28522,
        64'h543510a0_80ef31e5,
        64'h05130000_a51700f4,
        64'hcf63445c_358050ef,
        64'h32050513_0000a517,
        64'h85a6842a_c11dfda0,
        64'h0413e47f_f0ef84ae,
        64'hf406ec26_f0227179,
        64'h80826145_694264e2,
        64'h740270a2_85221440,
        64'h80ef6522_390050ef,
        64'h34850513_0000a517,
        64'h864a608c_ed01842a,
        64'he45ff0ef_84aa85ca,
        64'h0030c11d_fda00413,
        64'he8dff0ef_892eec26,
        64'hf406e84a_f0227179,
        64'hb7d92405_182080ef,
        64'h65223ce0_50ef854e,
        64'h85a20127_896300c7,
        64'hc78367a2_ed09e83f,
        64'hf0ef8526_85a20030,
        64'h80826121_69e27902,
        64'h74a27442_70e200f4,
        64'h496344dc_3a498993,
        64'h0000a997_0ff00913,
        64'h440184aa_cd01eebf,
        64'hf0efec4e_f04af426,
        64'hf822fc06_7139bfd5,
        64'h54798082_61457402,
        64'h70a28522_1e8080ef,
        64'h00f70963_00c54703,
        64'h0ff00793_6562e911,
        64'h842aee7f_f0ef0830,
        64'h65a2c105_fda00413,
        64'hf2dff0ef_e42ef406,
        64'hf0227179_b7c1fda0,
        64'h0513bf65_24052220,
        64'h80ef4981_65224720,
        64'h50ef8552_00099563,
        64'h2485cb99_0087c783,
        64'h67a2ed19_f29ff0ef,
        64'h854a85a2_00308082,
        64'h61216a42_69e27902,
        64'h74a27442_70e25535,
        64'he0914501_00f44d63,
        64'h00c92783_28ca0a13,
        64'h0000ba17_44014481,
        64'h4985892a_cd31f9bf,
        64'hf0efe852_ec4ef04a,
        64'hf426f822_fc067139,
        64'hbfe54501_80820141,
        64'h60a26108_c509fbbf,
        64'hf0efe406_1141b7f5,
        64'h02870713_fea68de3,
        64'h47148082_853a4701,
        64'h00e79563_97ba02d7,
        64'h87b30280_069302d7,
        64'h87bb878d_8f997c67,
        64'h87930000_b7976294,
        64'h7d070713_0000b717,
        64'h70868693_0000b697,
        64'hb7edfda0_07138302,
        64'h853e85b2_00030563,
        64'h01853303_8082853a,
        64'he21c97b6_470102a7,
        64'h87b30a00_051300b7,
        64'hd963454c_0005cc63,
        64'h5735c285_87ae6914,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h000a2e2e_2e746e65,
        64'h6d6f6d20_61207469,
        64'h61772065_7361656c,
        64'h50202165_6e616972,
        64'h41206d6f_7266206f,
        64'h6c6c6548_ffdff06f,
        64'h10500073_34102373,
        64'h342022f3_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_67a090ef,
        64'hfec5c6e3_02058593,
        64'h0005bc23_0005b823,
        64'h0005b423_0005b023,
        64'h1c860613_0000c617,
        64'ha3058593_0000c597,
        64'h30579073_09078793,
        64'h00000797_00078067,
        64'h40b787b3_00d787b3,
        64'h01478793_00000797,
        64'hfcc5cce3_02068693,
        64'h02058593_00e6bc23,
        64'h0185b703_00e6b823,
        64'h0105b703_00e6b423,
        64'h0085b703_00e6b023,
        64'h0005b703_0006b703,
        64'hff810113_01b11113,
        64'h0110011b_fe0e9ae3,
        64'h0085b703_fffe8e93,
        64'h0005b703_240e8e9b,
        64'h000f4eb7_01169693,
        64'hfff6869b_000066b7,
        64'h9c560613_0000c617,
        64'hfc058593_00000597,
        64'h000280e7_13050513,
        64'h00000517_0b228293,
        64'h00008297_000280e7,
        64'h08c28293_00008297,
        64'h01111113_fff1011b,
        64'h00006137_11249463,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
