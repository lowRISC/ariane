/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module etherboot (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 5906;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'hbffe7060_00000000,
        64'hbffe709e_00000000,
        64'h00000000_ffffffff,
        64'h00000006_00000000,
        64'hbffeb1e0_cc33aa55,
        64'h00000000_2f7c5c2d,
        64'h00000000_bffeb028,
        64'h00000000_ffffffff,
        64'h00006772_615f6473,
        64'h0000646d_635f6473,
        64'h00000000_0c000000,
        64'h00000000_ffffffff,
        64'h00000000_00000000,
        64'h00000000_30000000,
        64'h00000000_004b4d47,
        64'h00004b4d_47545045,
        64'h00000003_0f060301,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'haaaaaaaa_aaaaaaaa,
        64'h55555555_55555555,
        64'h5851f42d_4c957f2d,
        64'h10000000_20000000,
        64'h10325476_98badcfe,
        64'hefcdab89_67452301,
        64'hcccccccc_cccccccd,
        64'h00000a0d_70617274,
        64'h00000000_000a7473,
        64'h65742065_68636143,
        64'h00000000_00000a74,
        64'h6f6f6220_50544654,
        64'h00000000_00000a74,
        64'h73657420_4d415244,
        64'h00000000_00000000,
        64'h0a746f6f_62204453,
        64'h00000000_0000000a,
        64'h5825203d_20646565,
        64'h73206d6f_646e6152,
        64'h000a5825_2c582520,
        64'h3d20676e_69747465,
        64'h73206863_74697753,
        64'h00000000_00000a78,
        64'h25203d20_5d64255b,
        64'h4d454f20_49505351,
        64'h0000000a_5825203d,
        64'h205d6425_5b707773,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00000000,
        64'h0a646c25_2e646c25,
        64'h203d2049_5043202c,
        64'h73656c63_79632064,
        64'h6c25202c_736e6f69,
        64'h74637572_74736e69,
        64'h20646c25_202c424b,
        64'h6425203d_20746573,
        64'h5f676e69_6b726f77,
        64'h00000000_00000000,
        64'h0a2e2979_6c6e6f28,
        64'h2032206e_6f697372,
        64'h65762065_736e6563,
        64'h694c2063_696c6275,
        64'h50206c61_72656e65,
        64'h4720554e_47206568,
        64'h74207265_646e7520,
        64'h6465736e_6563694c,
        64'h00000000_0000000a,
        64'h2e6e6f62_617a6143,
        64'h2073656c_72616843,
        64'h20323130_322d3130,
        64'h30322029_43282074,
        64'h68676972_79706f43,
        64'h00000000_0000000a,
        64'h29746962_2d642528,
        64'h20302e33_2e34206e,
        64'h6f697372_65762072,
        64'h65747365_746d656d,
        64'h00000a74_73657420,
        64'h4d415244_206c6174,
        64'h656d2065_7261420a,
        64'h00000a2e_656e6f44,
        64'h00000000_000a6b6f,
        64'h0000203a_73252020,
        64'h00000073_73657264,
        64'h6441206b_63757453,
        64'h00000000_00000a3a,
        64'h00000000_0075252f,
        64'h00752520_706f6f4c,
        64'h00000000_000a7025,
        64'h7830206f_74207025,
        64'h78302073_69206567,
        64'h6e617220_74736574,
        64'h00000000_00082008,
        64'h00000000_00000008,
        64'h08080808_08080808,
        64'h08082020_20202020,
        64'h20202020_20080808,
        64'h08080808_08080808,
        64'h00000000_0000000a,
        64'h2e2e2e74_73657420,
        64'h7478656e_206f7420,
        64'h676e6970_70696b53,
        64'h00000000_000a2e78,
        64'h25783020_74657366,
        64'h666f2074_6120656e,
        64'h696c2073_73657264,
        64'h64612064_61622065,
        64'h6c626973_736f7020,
        64'h3a455255_4c494146,
        64'h00000000_00007525,
        64'h20676e69_74736574,
        64'h00000000_00007525,
        64'h20676e69_74746573,
        64'h00000000_00080808,
        64'h08080808_08080808,
        64'h00000000_00202020,
        64'h20202020_20202020,
        64'h00000000_0000000a,
        64'h7025203d_20327020,
        64'h2c702520_3d203170,
        64'h00000a2e_78257830,
        64'h20746573_66666f20,
        64'h74612078_25783020,
        64'h3d212078_25783020,
        64'h3a455255_4c494146,
        64'h00000000_000a7325,
        64'h206e6f69_74636e75,
        64'h66202c64_2520656e,
        64'h696c202c_73252065,
        64'h6c696620_2c64656c,
        64'h69616620_7325206e,
        64'h6f697472_65737361,
        64'h00000a72_6564616f,
        64'h6c20746f_6f622065,
        64'h67617473_20747372,
        64'h69662064_65736162,
        64'h20746f6f_622d750a,
        64'h00000000_5c2d2f7c,
        64'h00000000_64252065,
        64'h646f6320_68746977,
        64'h2064656c_69616620,
        64'h64616572_20666c65,
        64'h000a7972_6f6d656d,
        64'h20524444_206f7420,
        64'h666c6520_64616f6c,
        64'h00000000_00000000,
        64'h0a2e7365_74796220,
        64'h64252066_6f206e69,
        64'h622e746f_6f62206d,
        64'h6f726620_78252073,
        64'h73657264_64612079,
        64'h726f6d65_6d206f74,
        64'h20736574_79622064,
        64'h25206465_64616f4c,
        64'h00000000_216b7369,
        64'h6420746e_756f6d75,
        64'h206f7420_6c696166,
        64'h00000000_0021656c,
        64'h69662065_736f6c63,
        64'h206f7420_6c696166,
        64'h0000000a_21746f6f,
        64'h62206e65_706f206f,
        64'h74206465_6c696146,
        64'h00000000_00000000,
        64'h6e69622e_746f6f62,
        64'h00000000_00000a79,
        64'h726f6d65_6d206f74,
        64'h6e69206e_69622e74,
        64'h6f6f6220_64616f4c,
        64'h00000000_0000000a,
        64'h21726576_69726420,
        64'h44532074_6e756f6d,
        64'h206f7420_6c696146,
        64'h00000000_00000000,
        64'h0a2e6e6f_69746172,
        64'h65706f20_50544654,
        64'h206c6167_656c6c49,
        64'h00000000_000a2e64,
        64'h656c6c61_63207172,
        64'h775f656c_646e6168,
        64'h00000000_00000a2e,
        64'h646e6520_656c6966,
        64'h20657669_65636552,
        64'h00000000_00000000,
        64'h0a64253d_657a6973,
        64'h6b636f6c_62202c22,
        64'h73252220_3a717277,
        64'h00000000_0000002f,
        64'h00000000_000a646c,
        64'h25202e67_6e6f6c20,
        64'h6f6f7420_68746170,
        64'h20747365_75716552,
        64'h00000000_00000000,
        64'h0a732520_3d202964,
        64'h252c7025_2835646d,
        64'h00000000_0000000a,
        64'h6425203d_20687467,
        64'h6e656c20_656c6946,
        64'h00000000_00636d6d,
        64'h00000029_73252820,
        64'h00006425_203a7325,
        64'h00000000_00004453,
        64'h00000000_434d4d65,
        64'h00000000_00000000,
        64'h0a646e75_6f662074,
        64'h6f6e2064_25206563,
        64'h69766544_20434d4d,
        64'h0000297a_484d3030,
        64'h32282030_30325348,
        64'h00000000_00297a48,
        64'h4d383032_28203430,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282030,
        64'h35524444_20534855,
        64'h00000000_0000297a,
        64'h484d3030_31282030,
        64'h35524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282035,
        64'h32524453_20534855,
        64'h00000000_00000029,
        64'h7a484d35_32282032,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d32_35282032,
        64'h35524444_20434d4d,
        64'h0000297a_484d3235,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000029_7a484d30,
        64'h35282064_65657053,
        64'h20686769_48204453,
        64'h0000297a_484d3632,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000000_00000079,
        64'h63616765_4c204453,
        64'h00000000_00007963,
        64'h6167656c_20434d4d,
        64'h00000064_252e6425,
        64'h00000000_63256325,
        64'h63256325_63256325,
        64'h00000078_34302578,
        64'h34302520_726e5320,
        64'h78363025_206e614d,
        64'h00000000_00000a21,
        64'h646e756f_66206473,
        64'h635f7478_65206f4e,
        64'h00000000_00000000,
        64'h0a65646f_6d206120,
        64'h7463656c_6573206f,
        64'h7420656c_62616e75,
        64'h00000000_00000000,
        64'h0a217463_656c6573,
        64'h20656761_746c6f76,
        64'h206f7420_646e6f70,
        64'h73657220_746f6e20,
        64'h64696420_64726143,
        64'h0000000a_746e6573,
        64'h65727020_64726163,
        64'h206f6e20_3a434d4d,
        64'h00000000_0000000a,
        64'h64656e6f_69746974,
        64'h72617020_79646165,
        64'h726c6120_64726143,
        64'h00000000_000a7367,
        64'h6e697474_65732079,
        64'h74696c69_6261696c,
        64'h65722065_74697277,
        64'h206e6f69_74697472,
        64'h61702064_656c6c6f,
        64'h72746e6f_63207473,
        64'h6f682074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000a29_7525203e,
        64'h20752528_206d756d,
        64'h6978616d_20736465,
        64'h65637865_20657a69,
        64'h73206465_636e6168,
        64'h6e65206c_61746f54,
        64'h00000000_0000000a,
        64'h65747562_69727474,
        64'h61206465_636e6168,
        64'h6e652074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0a64656e,
        64'h67696c61_20657a69,
        64'h73207075_6f726720,
        64'h50572043_4820746f,
        64'h6e206e6f_69746974,
        64'h72617020_69255047,
        64'h0000000a_64656e67,
        64'h696c6120_657a6973,
        64'h2070756f_72672050,
        64'h57204348_20746f6e,
        64'h20616572_61206465,
        64'h636e6168_6e652061,
        64'h74616420_72657355,
        64'h00000a65_7a697320,
        64'h70756f72_67205057,
        64'h20434820_656e6966,
        64'h65642074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_000a676e,
        64'h696e6f69_74697472,
        64'h61702074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0000000a,
        64'h61657261_20617461,
        64'h64207265_73752064,
        64'h65636e61_686e6520,
        64'h726f6620_64657269,
        64'h75716572_20342e34,
        64'h203d3e20_434d4d65,
        64'h00000000_000a2978,
        64'h6c257830_2878616d,
        64'h20736465_65637865,
        64'h20786c25_78302072,
        64'h65626d75_6e206b63,
        64'h6f6c6220_3a434d4d,
        64'h00000000_00000a64,
        64'h6d632070_6f747320,
        64'h646e6573_206f7420,
        64'h6c696166_20636d6d,
        64'h00000000_000a7964,
        64'h61657220_64726163,
        64'h20676e69_74696177,
        64'h2074756f_656d6954,
        64'h0000000a_58383025,
        64'h7830203a_726f7272,
        64'h45207375_74617453,
        64'h00000000_65646f6d,
        64'h206e776f_6e6b6e55,
        64'h00000000_00006473,
        64'h5f637369_72776f6c,
        64'h00000078_25782520,
        64'h00000020_3a78250a,
        64'h00000000_0a732574,
        64'h69622d64_25203a68,
        64'h74646957_20737542,
        64'h00000000_0000203a,
        64'h79746963_61706143,
        64'h00000000_00000a73,
        64'h25203a79_74696361,
        64'h70614320_68676948,
        64'h00000a64_25203a64,
        64'h65657053_20737542,
        64'h00000000_00000a20,
        64'h63256325_63256325,
        64'h6325203a_656d614e,
        64'h00000000_00000000,
        64'h0a782520_3a4d454f,
        64'h00000000_0a782520,
        64'h3a444920_72657275,
        64'h74636166_756e614d,
        64'h00000000_000a7325,
        64'h203a6563_69766544,
        64'h00202020_3a434d4d,
        64'h00000000_52444420,
        64'h00000000_00006f4e,
        64'h00000000_00736559,
        64'h0000000a_7825203d,
        64'h2074736f_68202c78,
        64'h25207461_20646574,
        64'h61657263_20636d6d,
        64'h00000000_00000a64,
        64'h25206f74_20646567,
        64'h6e616863_206b7361,
        64'h6d202c64_65747265,
        64'h736e6920_64726143,
        64'h00000000_0000000a,
        64'h6425206f_74206465,
        64'h676e6168_63206b73,
        64'h616d202c_6465766f,
        64'h6d657220_64726143,
        64'h000a7475_6f656d69,
        64'h74207325_203a6473,
        64'h5f637369_72776f6c,
        64'h00726464_615f6573,
        64'h61625f64_73203d3d,
        64'h20657361_625f6473,
        64'h00000000_00000063,
        64'h2e636d6d_5f637369,
        64'h72776f6c_2f637273,
        64'h00000000_00000000,
        64'h66656463_62613938,
        64'h37363534_33323130,
        64'h007f7c5d_5b3f3e3d,
        64'h3c3b3a2e_2c2b2a22,
        64'h00007f7c_5d5b3f3e,
        64'h3d3c3b3a_2c2b2a22,
        64'h00000000_0a2e2e2e,
        64'h20726574_6f6f6220,
        64'h2c657962_646f6f47,
        64'h00000000_000a2e2e,
        64'h2e6d6172_676f7270,
        64'h20646564_616f6c20,
        64'h65687420_746f6f42,
        64'h00000000_00000000,
        64'h0a646c25_203d2073,
        64'h75746174_73207470,
        64'h75727265_746e6920,
        64'h74656e72_65687445,
        64'h0000000a_2e783230,
        64'h253a7832_30253a78,
        64'h3230253a_78323025,
        64'h3a783230_253a7832,
        64'h3025203d_20737365,
        64'h72646461_2043414d,
        64'h00000a78_6c253a78,
        64'h6c25203d_2043414d,
        64'h000a7264_64612043,
        64'h414d2070_75746553,
        64'h0000000a_21747075,
        64'h72726574_6e692064,
        64'h656c646e_61686e75,
        64'h00000000_00000a78,
        64'h25783020_3d206570,
        64'h79745f6f_746f7270,
        64'h00000000_0a297825,
        64'h28206465_74726f70,
        64'h7075736e_75203d20,
        64'h6f746f72_70205049,
        64'h000a5741_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a534c50_4d203d20,
        64'h6f746f72_50205049,
        64'h00000000_000a4554,
        64'h494c5044_55203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505443_53203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a504d4f_43203d20,
        64'h6f746f72_50205049,
        64'h00000000_0000004d,
        64'h00000000_0000000a,
        64'h5041434e_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000a48,
        64'h50544545_42203d20,
        64'h6f746f72_50205049,
        64'h000a5054_4d203d20,
        64'h6f746f72_50205049,
        64'h00000a48_41203d20,
        64'h6f746f72_50205049,
        64'h000a5053_45203d20,
        64'h6f746f72_50205049,
        64'h000a4552_47203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505653_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000036,
        64'h00000000_00000000,
        64'h0a504343_44203d20,
        64'h6f746f72_50205049,
        64'h00000a50_54203d20,
        64'h6f746f72_50205049,
        64'h000a5044_49203d20,
        64'h6f746f72_50205049,
        64'h000a3a73_746e6574,
        64'h6e6f6320_74736574,
        64'h0000000a_3a726564,
        64'h61656820_74736574,
        64'h000a5055_50203d20,
        64'h6f746f72_50205049,
        64'h000a5047_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000054,
        64'h00000000_00000000,
        64'h0a504950_49203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000047,
        64'h00006425_2b544553,
        64'h46464f5f_524c5052,
        64'h00000000_3f3f3f3f,
        64'h00000000_00544553,
        64'h46464f5f_524c5052,
        64'h00000000_00544553,
        64'h46464f5f_44414252,
        64'h00000000_00005445,
        64'h5346464f_5f525352,
        64'h00000000_00544553,
        64'h46464f5f_53434652,
        64'h00544553_46464f5f,
        64'h4c525443_4f49444d,
        64'h00000000_00544553,
        64'h46464f5f_53434654,
        64'h00000000_00544553,
        64'h46464f5f_524c5054,
        64'h00000000_54455346,
        64'h464f5f49_4843414d,
        64'h00000000_54455346,
        64'h464f5f4f_4c43414d,
        64'h00000000_000a3b29,
        64'h78257830_2c302c78,
        64'h25287465_736d656d,
        64'h00000a3b_29782578,
        64'h302c7825_78302c78,
        64'h25287970_636d656d,
        64'h000a7825_203d206c,
        64'h61757463_61202c58,
        64'h25203d20_64657269,
        64'h75716572_206e656c,
        64'h00000020_3a5d6425,
        64'h5b6e6f69_74636553,
        64'h000a7325_20202020,
        64'h00786c6c_2a302520,
        64'h00003a78_6c383025,
        64'h00732542_69632520,
        64'h00000000_00732573,
        64'h65747942_20756c25,
        64'h0073257a_48632520,
        64'h00000000_646c252e,
        64'h00000000_00756c25,
        64'h00000000_00000000,
        64'h73257a48_20756c25,
        64'h00000000_00007325,
        64'h00000000_00732520,
        64'h3a646c69_7542202c,
        64'h00000000_73257325,
        64'h00000000_00000a0a,
        64'h00000058_32302520,
        64'h00000000_0000002e,
        64'h00000000_00006325,
        64'h00000000_00000020,
        64'h20202020_20202020,
        64'h000a5245_46464f5f,
        64'h50434844_20726f66,
        64'h20676e69_74696157,
        64'h00000a73_25203a73,
        64'h25206563_69766564,
        64'h206e6f20_59524556,
        64'h4f435349_44205043,
        64'h48442064_6e657320,
        64'h74276e64_6c756f43,
        64'h000a5832_30253a58,
        64'h3230253a_58323025,
        64'h3a583230_253a5832,
        64'h30253a58_32302520,
        64'h3a204341_4d207325,
        64'h00000000_30687465,
        64'h00000000_000a2973,
        64'h2528726f_72726570,
        64'h000a5952_45564f43,
        64'h5349445f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_0000000a,
        64'h64252065_646f6370,
        64'h6f205043_48442064,
        64'h656c646e_61686e55,
        64'h00000000_0a642520,
        64'h6e6f6974_706f2064,
        64'h656c646e_61686e75,
        64'h00000000_0000000a,
        64'h73252072_6f727245,
        64'h00000000_00000a64,
        64'h65737566_65722073,
        64'h73657264_64612064,
        64'h65747365_75716552,
        64'h00000000_0000000a,
        64'h4b414e20_50434844,
        64'h00000000_0a444550,
        64'h50494b53_204b4341,
        64'h000a2273_2522203d,
        64'h20656d61_6e74736f,
        64'h4820746e_65696c43,
        64'h00000a22_73252220,
        64'h3d206e69_616d6f44,
        64'h00000000_0000000a,
        64'h7364253a_6d64253a,
        64'h68642520_3d20656d,
        64'h69742065_7361654c,
        64'h000a6425_2e64252e,
        64'h64252e64_2520203a,
        64'h73736572_64646120,
        64'h6b73616d_2074654e,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h61207265_74756f52,
        64'h00000000_00000000,
        64'h0a64252e_64252e64,
        64'h252e6425_20203a73,
        64'h73657264_64412050,
        64'h49207265_76726553,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h41205049_20746e65,
        64'h696c4320_50434844,
        64'h00000000_0000000a,
        64'h4b434120_50434844,
        64'h0000000a_54534555,
        64'h5145525f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_00000000,
        64'h0a702520_2c726f72,
        64'h7265206c_616e7265,
        64'h746e6920_70636864,
        64'h00000a29_73252c73,
        64'h25287075_6b6f6f6c,
        64'h000a6563_69766564,
        64'h206e776f_6e6b6e75,
        64'h00000000_203a6425,
        64'h20656369_7665440a,
        64'h00203a64_25206563,
        64'h69766564_2073250a,
        64'h00000000_00203a64,
        64'h25206563_69766544,
        64'h00000000_00000000,
        64'h73736572_6464612d,
        64'h63616d2d_6c61636f,
        64'h6c006874_6469772d,
        64'h6f692d67_65720074,
        64'h66696873_2d676572,
        64'h00737470_75727265,
        64'h746e6900_746e6572,
        64'h61702d74_70757272,
        64'h65746e69_00646565,
        64'h70732d74_6e657272,
        64'h75630076_65646e2c,
        64'h76637369_72007974,
        64'h69726f69_72702d78,
        64'h616d2c76_63736972,
        64'h0073656d_616e2d67,
        64'h65720064_65646e65,
        64'h7478652d_73747075,
        64'h72726574_6e690073,
        64'h65676e61_7200656c,
        64'h646e6168_702c7875,
        64'h6e696c00_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h00100000_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_00000064,
        64'h6e727768_2d637369,
        64'h72776f6c_1b000000,
        64'h0e000000_03000000,
        64'h00003030_30303030,
        64'h30344064_6e727768,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h00800000_00000000,
        64'h00000030_00000000,
        64'h67000000_10000000,
        64'h03000000_00007fe3,
        64'h023e1800_47010000,
        64'h06000000_03000000,
        64'h03000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_00636d6d,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_02000000,
        64'h25010000_04000000,
        64'h03000000_02000000,
        64'h14010000_04000000,
        64'h03000000_00000100,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40636d6d,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h04000000_3a010000,
        64'h04000000_03000000,
        64'h02000000_30010000,
        64'h04000000_03000000,
        64'h01000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h00c20100_06010000,
        64'h04000000_03000000,
        64'h80f0fa02_4b000000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000010_00000000,
        64'h67000000_10000000,
        64'h03000000_00303537,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000000,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'hffff0000_01000000,
        64'hca000000_08000000,
        64'h03000000_00333130,
        64'h2d677562_65642c76,
        64'h63736972_1b000000,
        64'h10000000_03000000,
        64'h00003040_72656c6c,
        64'h6f72746e_6f632d67,
        64'h75626564_01000000,
        64'h02000000_02000000,
        64'hbb000000_04000000,
        64'h03000000_02000000,
        64'hb5000000_04000000,
        64'h03000000_03000000,
        64'hfb000000_04000000,
        64'h03000000_07000000,
        64'he8000000_04000000,
        64'h03000000_00000004,
        64'h00000000_0000000c,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h09000000_01000000,
        64'h0b000000_01000000,
        64'hca000000_10000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00000c00,
        64'h00000000_00000002,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_01000000,
        64'h03000000_01000000,
        64'hca000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6e696c63,
        64'h01000000_c3000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h01000000_bb000000,
        64'h04000000_03000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00007663_73697200,
        64'h656e6169_7261202c,
        64'h7a687465_1b000000,
        64'h13000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha8060000_59010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'he0060000_38000000,
        64'h39080000_edfe0dd0,
        64'h00000000_64726143,
        64'h2d445320_726f6620,
        64'h746f6f62_2d752064,
        64'h6573696d_696e696d,
        64'h20435349_52776f4c,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00020000_00010000,
        64'h0000c000_00008000,
        64'h00006000_00004000,
        64'h00002000_00001000,
        64'h00000800_00000400,
        64'h00000200_00000100,
        64'h00000080_00000040,
        64'h00000020_00000000,
        64'h0bebc200_0c65d400,
        64'h02faf080_05f5e100,
        64'h02faf080_017d7840,
        64'h03197500_03197500,
        64'h02faf080_018cba80,
        64'h017d7840_017d7840,
        64'h00989680_000f4240,
        64'h000186a0_00002710,
        64'h50463c37_322d2823,
        64'h1e19140f_0d0c0a00,
        64'h00000000_00000000,
        64'h00000000_10000000,
        64'h00000001_00000000,
        64'h20000000_00000002,
        64'h00000000_40000000,
        64'h00000005_00000001,
        64'h20000000_00000006,
        64'h00000001_40000000,
        64'h70000000_00000000,
        64'h70000000_00000002,
        64'h70000000_00000004,
        64'h60000000_00000005,
        64'h30000000_00000001,
        64'h30000000_00000003,
        64'h00000000_40050100,
        64'h40050000_40040500,
        64'h40040401_40040400,
        64'h40040300_40040200,
        64'h40040100_40040000,
        64'h00000000_bffeb190,
        64'h00000000_bffeb178,
        64'h00000000_bffeb160,
        64'h00000000_bffeb148,
        64'h00000000_bffeb130,
        64'h00000000_bffeb118,
        64'h00000000_bffeb100,
        64'h00000000_bffeb0e8,
        64'h00000000_bffeb0d0,
        64'h00000000_bffeb0b8,
        64'h00000000_bffeb0a8,
        64'h00000000_bffeb098,
        64'hffffbd8c_ffffbd8c,
        64'hffffbd8c_ffffbd8c,
        64'hffffbd88_ffffbd84,
        64'hffffbd84_ffffbd5e,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_bffe4d12,
        64'h00000000_bffe4ab4,
        64'h00000000_bffe4ea6,
        64'h00646374_65675f63,
        64'h6d6d5f64_72616f62,
        64'h00000002_0000ffff,
        64'h004c4b40_004c4b40,
        64'h00300000_20000000,
        64'h00000000_bffe9a88,
        64'h00000000_bffead80,
        64'h00717269_5f646e65,
        64'h5f617461_645f6473,
        64'h5f637369_72776f6c,
        64'h00000000_00007172,
        64'h695f646d_635f6473,
        64'h5f637369_72776f6c,
        64'h00007172_695f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0067616c,
        64'h665f7470_75727265,
        64'h746e695f_74696177,
        64'h5f637369_72776f6c,
        64'h00000000_646d635f,
        64'h74726174_735f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0000006e,
        64'h655f7172_695f6473,
        64'h00000000_00007475,
        64'h6f656d69_745f6473,
        64'h00000000_0000657a,
        64'h69736b6c_625f6473,
        64'h00000000_00000074,
        64'h6e636b6c_625f6473,
        64'h00000000_00000000,
        64'h74657365_725f6473,
        64'h00000000_74726174,
        64'h735f646d_635f6473,
        64'h00000000_0000676e,
        64'h69747465_735f6473,
        64'h00000000_00007669,
        64'h645f6b6c_635f6473,
        64'h00000000_00000000,
        64'h6e67696c_615f6473,
        64'h00000000_00006465,
        64'h6c5f7465_735f6473,
        64'h5f637369_72776f6c,
        64'h09020b04_0d060f08,
        64'h010a030c_050e0700,
        64'h020f0c09_0603000d,
        64'h0a070401_0e0b0805,
        64'h0c07020d_08030e09,
        64'h040f0a05_000b0601,
        64'heb86d391_2ad7d2bb,
        64'hbd3af235_f7537e82,
        64'h4e0811a1_a3014314,
        64'hfe2ce6e0_6fa87e4f,
        64'h85845dd1_ffeff47d,
        64'h8f0ccc92_655b59c3,
        64'hfc93a039_ab9423a7,
        64'h432aff97_f4292244,
        64'hc4ac5665_1fa27cf8,
        64'he6db99e5_d9d4d039,
        64'h04881d05_d4ef3085,
        64'heaa127fa_289b7ec6,
        64'hbebfbc70_f6bb4b60,
        64'h4bdecfa9_a4beea44,
        64'hfde5380c_6d9d6122,
        64'h8771f681_fffa3942,
        64'h8d2a4c8a_676f02d9,
        64'hfcefa3f8_a9e3e905,
        64'h455a14ed_f4d50d87,
        64'hc33707d6_21e1cde6,
        64'he7d3fbc8_d8a1e681,
        64'h02441453_d62f105d,
        64'he9b6c7aa_265e5a51,
        64'hc040b340_f61e2562,
        64'h49b40821_a679438e,
        64'hfd987193_6b901122,
        64'h895cd7be_ffff5bb1,
        64'h8b44f7af_698098d8,
        64'hfd469501_a8304613,
        64'h4787c62a_f57c0faf,
        64'hc1bdceee_242070db,
        64'he8c7b756_d76aa478,
        64'h02020202_02020202,
        64'h10020202_02020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02010101_01010101,
        64'h10010101_01010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h08101010_10020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02424242_42424210,
        64'h10101010_10010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h01414141_41414110,
        64'h10101010_10100404,
        64'h04040404_04040404,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h08080808_08080808,
        64'h08080808_08080808,
        64'h08082828_28282808,
        64'h08080808_08080808,
        64'h00000000_0000b7e9,
        64'he2bff0ef_8b2fc0ef,
        64'h04850513_00002517,
        64'hbff1ec0f_80ef8c4f,
        64'hc0ef04a5_05130000,
        64'h2517b7fd_d53ff0ef,
        64'h8d6fc0ef_04c50513,
        64'h00002517_a001b43f,
        64'he0ef8522_8eafc0ef,
        64'h05050513_00002517,
        64'h00e78c63_470504e7,
        64'h8163470d_02e78b63,
        64'h47090064_57930ff4,
        64'h7413fd39_1be3914f,
        64'hc0ef2581_8552688c,
        64'h0004b823_922fc0ef,
        64'h86222401_25816080,
        64'h608ce09c_09058556,
        64'h0007c783_016907b3,
        64'h499108aa_0a130000,
        64'h2a1707aa_8a930000,
        64'h2a974000_04b7216b,
        64'h0b130000_2b174901,
        64'hfc941ee3_962fc0ef,
        64'h2405854a_85a2862a,
        64'hf43ff0ef_c03e04b0,
        64'h05134585_4601868a,
        64'h0137e7b3_0204079b,
        64'h44990a29_09130000,
        64'h29170200_09b74401,
        64'hfe9416e3_99afc0ef,
        64'h0405854a_0004059b,
        64'h6390078e_013407b3,
        64'h44950ba9_09130000,
        64'h29170800_09b74401,
        64'haddfe0ef_0bc50513,
        64'h00002517_ab7fe0ef,
        64'he15ae556_e952ed4e,
        64'hf14af526_f922fd06,
        64'h7131afff_e06f1865,
        64'h05130000_2517bfe1,
        64'hf7100691_27850006,
        64'he6038082_73884000,
        64'h07b7ffe5_37fdc319,
        64'h8b097a98_400006b7,
        64'h3e800793_00b7ef63,
        64'h40000737_47812581,
        64'hf7888d51_400007b7,
        64'h0106161b_8d5d0085,
        64'h979b8082_25017b88,
        64'h400007b7_80822501,
        64'h6b880007_b8234000,
        64'h07b78082_25016388,
        64'h400007b7_8082e388,
        64'h400007b7_91011502,
        64'hbff1f5df_f0ef4541,
        64'hf63ff0ef_4521f69f,
        64'hf0ef4511_f6fff0ef,
        64'h4509f75f_f0ef4505,
        64'hf7bff0ef_4501e406,
        64'h1141bf51_c00028f3,
        64'hc02026f3_fac710e3,
        64'ha96fc06f_14c50513,
        64'h00002517_02a74733,
        64'h02a767b3_02b345bb,
        64'h02c74733_40000593,
        64'h02a68733_411686b3,
        64'h3e800513_c00026f3,
        64'h8e15c020_267302b7,
        64'h1d632705_fe0813e3,
        64'h97aa387d_00078023,
        64'h97aa0007_802397aa,
        64'h00078023_97aa0007,
        64'h80234000_081387f2,
        64'h45a901f6_1e134681,
        64'h48814701_00c5131b,
        64'h46058082_80826145,
        64'h69a26942_64e27402,
        64'h70a2ff24_17e3e6df,
        64'hf0ef2405_01358533,
        64'h46054685_008495b3,
        64'h497901f4_99934441,
        64'hb36fc0ef_4485e665,
        64'h05130000_2517b44f,
        64'hc0ef1b25_05130000,
        64'h2517b50f_c0ef18e5,
        64'h05130000_2517b5cf,
        64'hc0ef1725_05130000,
        64'h25170400_0593c8bf,
        64'he0efe44e_e84aec26,
        64'hf022f406_17450513,
        64'h00002517_7179bfa1,
        64'h0485b88f_c0efeb65,
        64'h05130000_2517b7e9,
        64'h4a89b98f_c0ef1865,
        64'h05130000_25179782,
        64'h852285ce_6642008a,
        64'h3783bb0f_c0ef1965,
        64'h05130000_2517c58d,
        64'h000a3583_02f74963,
        64'h6762010a_2783bccf,
        64'hc0ef856e_ed15920f,
        64'hf0ef8522_65a2bdcf,
        64'hc0ef856a_85e6be4f,
        64'hc0ef8562_beafc0ef,
        64'h855e85ca_00090663,
        64'hbf6fc0ef_855a85a6,
        64'h80826149_7da27d42,
        64'h7ce26c06_6ba66b46,
        64'h6ae67a06_79a67946,
        64'h74e68556_640a60aa,
        64'hc1efc0ef_21450513,
        64'h00002517_02997863,
        64'had0a0a13_00003a17,
        64'h220d8d93_00002d97,
        64'h220d0d13_00002d17,
        64'h218c8c93_00002c97,
        64'h218c0c13_00002c17,
        64'h218b8b93_00002b97,
        64'h218b0b13_00002b17,
        64'h44854a81_e43e99a2,
        64'h0034d793_e83e0014,
        64'hd9930044_d793c7cf,
        64'hc0efec36_e506f46e,
        64'hf86afc66_e0e2e4de,
        64'he8daecd6_f0d2f4ce,
        64'h23050513_00002517,
        64'h85aa962a_84ae842a,
        64'hfca6e122_fff58613,
        64'h8932f8ca_71758082,
        64'h6505b789_547dbf29,
        64'h0d85ee5f_e0ef0007,
        64'hc50397ea_8b8d0007,
        64'h8b1b001b_079bef9f,
        64'he0ef4521_ef91034d,
        64'hf7b300f6_932393c1,
        64'h17c20064_d78300f6,
        64'h922393c1_17c20044,
        64'hd78300f6_912393c1,
        64'h17c20024_d78300f6,
        64'h902393c1_17c20004,
        64'hd783e388_66c267e2,
        64'hbca7bc23_00003797,
        64'h8d419101_14021502,
        64'h8c518d59_0106161b,
        64'h0105151b_67026622,
        64'h87efe0ef_e02a884f,
        64'he0efe42a_88afe0ef,
        64'h842a890f_e0efe836,
        64'hec3eb775_8c4a8bce,
        64'h4a858082_61497da2,
        64'h7d427ce2_6c066ba6,
        64'h6b466ae6_7a0679a6,
        64'h794674e6_640a60aa,
        64'h8522d78f_c0ef30e5,
        64'h05130000_2517020a,
        64'h8863e579_842aa82f,
        64'hf0ef854a_85ce866e,
        64'h059d9563_97de00fc,
        64'h06b3003d_97934d81,
        64'h8c4e8bca_664d0d13,
        64'h00002d17_9c4a0a13,
        64'hc7848493_00003497,
        64'h4a81fe5f_e0ef4b01,
        64'h8cb2f46e_e122e506,
        64'hf86afc66_e0e2e4de,
        64'he8daecd6_fca66a05,
        64'h02000513_89ae892a,
        64'hf0d2f4ce_f8ca7175,
        64'hbfa1547d_bf0d0d85,
        64'h81aff0ef_0007c503,
        64'h97e68b8d_00078a9b,
        64'h001a879b_82eff0ef,
        64'h4521ef91_0ba1033d,
        64'hf7b3ffa7_95e300d6,
        64'h00230ff6_f6930785,
        64'h00fb8633_0006c683,
        64'h018786b3_4781e288,
        64'hcea7b823_00003797,
        64'h8d4166e2_91011402,
        64'h15028c51_0106161b,
        64'h8d5d0105_151b6642,
        64'h67a29a0f_e0efe42a,
        64'h9a6fe0ef_e82a9acf,
        64'he0ef842a_9b2fe0ef,
        64'hec36b775_8ba68b4a,
        64'h4a058082_61497da2,
        64'h7d427ce2_6c066ba6,
        64'h6b466ae6_7a0679a6,
        64'h794674e6_640a60aa,
        64'h8522e98f_c0ef42e5,
        64'h05130000_2517020a,
        64'h0863ed45_842aba2f,
        64'hf0ef8526_85ca866e,
        64'h04fd9563_96da003d,
        64'h96936782_4d214d81,
        64'h8bca8b26_784c8c93,
        64'h00002c97_9c498993,
        64'hd90c0c13_00003c17,
        64'h4a01904f_f0ef4a81,
        64'he032f46e_f86ae122,
        64'he506fc66_e0e2e4de,
        64'he8daecd6_f0d26985,
        64'h02000513_892e84aa,
        64'hf4cef8ca_fca67175,
        64'hb7e95b7d_b7490605,
        64'h00b83023_e30c85d6,
        64'he11185e2_00167513,
        64'h80826109_6de27d02,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e67906,
        64'h74a6855a_744670e6,
        64'hf46fc0ef_4b450513,
        64'h00002517_fafb90e3,
        64'h04000793_2b85fbb4,
        64'h1be38c56_2405e931,
        64'h8b2ac5ef_f0ef854a,
        64'h85ce6622_f72fc0ef,
        64'h856a85da_f7afc0ef,
        64'he4328552_06f61063,
        64'h974e00e9_08330036,
        64'h17136782_4601fffc,
        64'h4a93f98f_c0ef8566,
        64'h85da0084_8b3bfa4f,
        64'hc0ef8552_4401003b,
        64'h949b0177_9c334785,
        64'h4da14bad_0d130000,
        64'h2d174b2c_8c930000,
        64'h2c974aaa_0a130000,
        64'h2a17fd0f_c0ef4b81,
        64'he03289ae_f862e0da,
        64'he4d6f4a6_f8a2fc86,
        64'hec6ef06a_f466fc5e,
        64'he8d2ecce_4c450513,
        64'h00002517_892af0ca,
        64'h7119bf75_5dfdbfc5,
        64'h85bafe08_1be385c6,
        64'hb7610605_e10ce28c,
        64'h85be0008_1363859a,
        64'h008bea63_00167813,
        64'h80826109_6de27d02,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e67906,
        64'h74a6856e_744670e6,
        64'h847fc0ef_5b450513,
        64'h00002517_f8f41be3,
        64'h08000793_2405ed29,
        64'h8daad56f_f0ef8526,
        64'h85ca6622_86bfc0ef,
        64'h856685a2_873fc0ef,
        64'he432854e_05461c63,
        64'h96ca00d4_85330036,
        64'h16934601_fff7c313,
        64'hfff74893_8fd5008d,
        64'h16b300fd_17b30024,
        64'h079b8f5d_00ed1733,
        64'h00fd17b3_408b07bb,
        64'h408a873b_8b3fc0ef,
        64'h856285a2_8bbfc0ef,
        64'h854e5c2c_8c930000,
        64'h2c9703f0_0b930810,
        64'h0b134d05_07f00a93,
        64'h5c8c0c13_00002c17,
        64'h5c098993_00002997,
        64'h8e7fc0ef_44018a32,
        64'h892eec6e_fc86f06a,
        64'hf466f862_fc5ee0da,
        64'he4d6e8d2_eccef0ca,
        64'hf8a25da5_05130000,
        64'h251784aa_f4a67119,
        64'hb7f15dfd_bfe5e19c,
        64'he31cbf61_0605e194,
        64'he314008c_66638082,
        64'h61096de2_7d027ca2,
        64'h7c427be2_6b066aa6,
        64'h6a4669e6_790674a6,
        64'h856e7446_70e694df,
        64'hc0ef6ba5_05130000,
        64'h2517fb54_17e32405,
        64'he1398daa_e58ff0ef,
        64'h852685ca_662296df,
        64'hc0ef856a_85a2975f,
        64'hc0efe432_85520566,
        64'h1a63974a_00e485b3,
        64'h00361713_4601fff6,
        64'hc693fff7_c7930089,
        64'h96b300f9_97b3408b,
        64'h87bb9a1f_c0ef8566,
        64'h85a29a9f_c0ef8552,
        64'h08000a93_6b4d0d13,
        64'h00002d17_03f00c13,
        64'h498507f0_0b936b6c,
        64'h8c930000_2c976aea,
        64'h0a130000_2a179d5f,
        64'hc0ef4401_8b32892e,
        64'hec6efc86_f06af466,
        64'hf862fc5e_e0dae4d6,
        64'he8d2ecce_f0caf8a2,
        64'h6c850513_00002517,
        64'h84aaf4a6_7119b7f1,
        64'h5dfdbfe5_e298e398,
        64'hbf610605_e28ce38c,
        64'h008c6663_80826109,
        64'h6de27d02_7ca27c42,
        64'h7be26b06_6aa66a46,
        64'h69e67906_74a6856e,
        64'h744670e6_a3bfc0ef,
        64'h7a850513_00002517,
        64'hfb541be3_2405e139,
        64'h8daaf46f_f0ef8526,
        64'h85ca6622_a5bfc0ef,
        64'h856a85a2_a63fc0ef,
        64'he4328552_05661a63,
        64'h97ca00f4_86b30036,
        64'h17934601_008995b3,
        64'h00e99733_408b873b,
        64'ha87fc0ef_856685a2,
        64'ha8ffc0ef_85520800,
        64'h0a9379ad_0d130000,
        64'h2d1703f0_0c134985,
        64'h07f00b93_79cc8c93,
        64'h00002c97_794a0a13,
        64'h00002a17_abbfc0ef,
        64'h44018b32_892eec6e,
        64'hfc86f06a_f466f862,
        64'hfc5ee0da_e4d6e8d2,
        64'heccef0ca_f8a27ae5,
        64'h05130000_251784aa,
        64'hf4a67119_bff159fd,
        64'hb74d0605_e29ce31c,
        64'h80826125_6c426be2,
        64'h7b027aa2_7a4279e2,
        64'h690664a6_854e6446,
        64'h60e6b11f_c0ef87e5,
        64'h05130000_3517f94c,
        64'h19e30c05_e91d89aa,
        64'h81dff0ef_852285a6,
        64'h6622b31f_c0ef855e,
        64'h85ceb39f_c0efe432,
        64'h854a0556_17639726,
        64'h00e406b3_00361713,
        64'h46018fd9_038c1713,
        64'h8fd9030c_17138fd9,
        64'h028c1713_8fd9020c,
        64'h17138fd9_018c1713,
        64'h0187e7b3_8fd9010c,
        64'h1793008c_1713b7df,
        64'hc0ef855a_85ce000c,
        64'h099bb89f_c0ef854a,
        64'h10000a13_894b8b93,
        64'h00003b97_88cb0b13,
        64'h00003b17_88490913,
        64'h00003917_babfc0ef,
        64'h4c018ab2_84aefc4e,
        64'hec86e862_ec5ef05a,
        64'hf456f852_e0cae4a6,
        64'h89850513_00003517,
        64'h842ae8a2_711db7e1,
        64'h5d7db779_0605e198,
        64'he398872a_c291876a,
        64'h00167693_bf49000b,
        64'h3d038082_61656d42,
        64'h6ce27c02_7ba27b42,
        64'h7ae26a06_69a66946,
        64'h64e6856a_740670a6,
        64'hc0ffc0ef_97c50513,
        64'h00003517_fb441ae3,
        64'h2405e529_8d2a91bf,
        64'hf0ef8526_85ca6622,
        64'hc2ffc0ef_856685a2,
        64'hc37fc0ef_e432854e,
        64'h05561c63_97ca00f4,
        64'h85b30036_1793fffd,
        64'h45134601_c53fc0ef,
        64'h856285a2_000bbd03,
        64'hcba50014_7793c65f,
        64'hc0ef854e_04000a13,
        64'h970c8c93_00003c97,
        64'h968c0c13_00003c17,
        64'hc58b8b93_00003b97,
        64'hc58b0b13_00003b17,
        64'h97098993_00003997,
        64'hc97fc0ef_44018ab2,
        64'h892ee86a_f486ec66,
        64'hf062f45e_f85afc56,
        64'he0d2e4ce_e8caf0a2,
        64'h98850513_00003517,
        64'h84aaeca6_7159bfc1,
        64'h54fdbf59_0605e198,
        64'he3988726_c2918766,
        64'h00167693_80826165,
        64'h6ce27c02_7ba27b42,
        64'h7ae26a06_69a664e6,
        64'h69468526_740670a6,
        64'hcf7fc0ef_a6450513,
        64'h00003517_fb541be3,
        64'h2405e129_84aaa03f,
        64'hf0ef854a_85ce6622,
        64'hd17fc0ef_856285a2,
        64'hd1ffc0ef_e4328552,
        64'h05661863_97ce00f9,
        64'h05b30036_179314fd,
        64'h46014090_0cb3d3df,
        64'hc0ef8885_855e85a2,
        64'hfff44493_d4bfc0ef,
        64'h85520400_0a93a56c,
        64'h0c130000_3c17a4eb,
        64'h8b930000_3b97a46a,
        64'h0a130000_3a17d6df,
        64'hc0ef4401_8b3289ae,
        64'hec66eca6_f486f062,
        64'hf45ef85a_fc56e0d2,
        64'he4cef0a2_a5c50513,
        64'h00003517_892ae8ca,
        64'h7159bfc9_070500a8,
        64'h3023e288_00f70533,
        64'ha9dff06f_6121863a,
        64'h69e2854e_790274a2,
        64'h70e27442_00c71c63,
        64'h96ae00d9_88330037,
        64'h16934701_8fc59081,
        64'h178265a2_66021482,
        64'h8fc18cc9_0109179b,
        64'h0105151b_92bfe0ef,
        64'h84aa931f_e0ef892a,
        64'h937fe0ef_842a93df,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7f100e8,
        64'h30238f69_00083703,
        64'he3148ee9_07856314,
        64'hb15ff06f_6121863e,
        64'h69e2854e_790274a2,
        64'h70e27442_00c79c63,
        64'h974e00e5_88330037,
        64'h97134781_8d5d9101,
        64'h178265a2_66021502,
        64'h8fc18d45_0109179b,
        64'h0105151b_9a3fe0ef,
        64'h84aa9a9f_e0ef892a,
        64'h9affe0ef_842a9b5f,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7f100e8,
        64'h30238f49_00083703,
        64'he3148ec9_07856314,
        64'hb8dff06f_6121863e,
        64'h69e2854e_790274a2,
        64'h70e27442_00c79c63,
        64'h974e00e5_88330037,
        64'h97134781_8d5d9101,
        64'h178265a2_66021502,
        64'h8fc18d45_0109179b,
        64'h0105151b_a1bfe0ef,
        64'h84aaa21f_e0ef892a,
        64'ha27fe0ef_842aa2df,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7d100e8,
        64'h302302a7_57330008,
        64'h3703e314_02a6d6b3,
        64'h07856314_4505e111,
        64'hc0dff06f_6121863e,
        64'h69e2854e_790274a2,
        64'h70e27442_00c79c63,
        64'h974e00e5_88330037,
        64'h97134781_8d5d9101,
        64'h178265a2_66021502,
        64'h8fc18d45_0109179b,
        64'h0105151b_a9bfe0ef,
        64'h84aaaa1f_e0ef892a,
        64'haa7fe0ef_842aaadf,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7e100e8,
        64'h302302a7_07330008,
        64'h3703e314_02a686b3,
        64'h07856314_c89ff06f,
        64'h6121863e_69e2854e,
        64'h790274a2_70e27442,
        64'h00c79c63_974e00e5,
        64'h88330037_97134781,
        64'h8d5d9101_178265a2,
        64'h66021502_8fc18d45,
        64'h0109179b_0105151b,
        64'hb17fe0ef_84aab1df,
        64'he0ef892a_b23fe0ef,
        64'h842ab29f_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7f100e8_30238f09,
        64'h00083703_e3148e89,
        64'h07856314_d01ff06f,
        64'h6121863e_69e2854e,
        64'h790274a2_70e27442,
        64'h00c79c63_974e00e5,
        64'h88330037_97134781,
        64'h8d5d9101_178265a2,
        64'h66021502_8fc18d45,
        64'h0109179b_0105151b,
        64'hb8ffe0ef_84aab95f,
        64'he0ef892a_b9bfe0ef,
        64'h842aba1f_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7f100e8_30238f29,
        64'h00083703_e3148ea9,
        64'h07856314_d79ff06f,
        64'h6121863e_69e2854e,
        64'h790274a2_70e27442,
        64'h00c79c63_974e00e5,
        64'h88330037_97134781,
        64'h8d5d9101_178265a2,
        64'h66021502_8fc18d45,
        64'h0109179b_0105151b,
        64'hc07fe0ef_84aac0df,
        64'he0ef892a_c13fe0ef,
        64'h842ac19f_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7ad0485_b0fff0ef,
        64'h0007c503_97e20039,
        64'hf7930985_b1fff0ef,
        64'h4521ef81_00adb023,
        64'h00acb023_8d419101,
        64'h14021502_01a46433,
        64'h00a96533_010d1d1b,
        64'h0105151b_0344f7b3,
        64'hc6ffe0ef_892ac75f,
        64'he0ef8d2a_c7bfe0ef,
        64'h842ac81f_e0efe33f,
        64'hf06f6165_7ae28556,
        64'h7b4264e6_85da8626,
        64'h6da26d42_6ce27c02,
        64'h7ba26a06_69a66946,
        64'h70a67406_962fd0ef,
        64'hef850513_00003517,
        64'h03749b63_00fb0cb3,
        64'h00fa8db3_00349793,
        64'h238c0c13_00003c17,
        64'h9c4a0a13_4981bb1f,
        64'hf0ef4481_8bb28b2e,
        64'he46ee86a_ec66e8ca,
        64'hf0a2f486_f062f45e,
        64'hf85ae4ce_eca60200,
        64'h05138aaa_6a05fc56,
        64'he0d27159_bfa507a1,
        64'h05858082_61256ca2,
        64'h6c426be2_7b027aa2,
        64'h7a4279e2_690664a6,
        64'h644660e6_557d9dcf,
        64'hd0eff2a5_05130000,
        64'h35179e8f_d0efefe5,
        64'h05130000_3517058e,
        64'h02e60d63_40e98733,
        64'h00359713_c689873e,
        64'h8a856390_008586b3,
        64'hbf5d07a1_04856398,
        64'he39840e9_87330034,
        64'h9713c689_873e8a85,
        64'h008486b3_a8894501,
        64'ha2efd0ef_f9c50513,
        64'h00003517_fd5417e3,
        64'h040502b4_9b634581,
        64'h87caa48f_d0ef8562,
        64'h85e6a50f_d0ef8552,
        64'h03649863_448187ca,
        64'ha5efd0ef_855e85e6,
        64'h00040c9b_a6afd0ef,
        64'h85524ac1_f74c0c13,
        64'h00003c17_fff94993,
        64'hf70b8b93_00003b97,
        64'hf68a0a13_00003a17,
        64'ha8efd0ef_44018b2e,
        64'he466e4a6_ec86e862,
        64'hec5ef05a_f456f852,
        64'hfc4ee8a2_f7c50513,
        64'h00003517_892ae0ca,
        64'h711dbf5d_0785a001,
        64'habefd0ef_f7c50513,
        64'h00003517_85a28626,
        64'hacefd0ef_f6450513,
        64'h00003517_6090600c,
        64'h02e80363_60980004,
        64'h38038082_61054501,
        64'h64a26442_60e200c7,
        64'h986300d5_043300d5,
        64'h84b30037_96934781,
        64'he426e822_ec061101,
        64'hc2dff06f_80824501,
        64'h80824501_80828082,
        64'h80828082_45098082,
        64'h45098082_4509bff9,
        64'h26052004_04136622,
        64'hedbfc0ef_e4328522,
        64'h85b28082_61454501,
        64'h64e27402_70a20096,
        64'h186300c6_84bb842e,
        64'hf406ec26_f0227179,
        64'h80824505_80824505,
        64'h80824505_80820141,
        64'h8d7d6402_60a29522,
        64'h408007b3_f57ff0ef,
        64'he406952e_842ae022,
        64'h1141a001_d2dff0ef,
        64'h4505b90f_d0efe406,
        64'hff050513_00003517,
        64'h85aa862e_86b28736,
        64'h11418082_02f55533,
        64'h47a9b000_25738082,
        64'h45018082_45018082,
        64'h01414501_60a2f89f,
        64'hc0ef2000_0537bccf,
        64'hd0efe406_00450513,
        64'h00003517_11418082,
        64'h80826105_644260e2,
        64'h85229e8f_f0ef4581,
        64'h6622c509_842afd1f,
        64'hf0efe432_8532ec06,
        64'he8221101_02b50633,
        64'h8082953e_055e10d0,
        64'h0513e308_95360017,
        64'h86930075_6513157d,
        64'h631c8827_07130000,
        64'h47178082_45018082,
        64'h24050513_000f4537,
        64'ha001ddbf_f0efe406,
        64'h25011141_90020000,
        64'h0023e8df_f0efc4cf,
        64'hd0ef83a5_05130000,
        64'h3517bddd_c5afd0ef,
        64'h06850513_00003517,
        64'hc981c62e_0005059b,
        64'h962f90ef_01849513,
        64'h85a2c78f_d0ef06e5,
        64'h05130000_3517c84f,
        64'hd0ef0325_05130000,
        64'h351785a2_01849613,
        64'h86a20bf0_0493bf1d,
        64'h03050513_00003517,
        64'hc5112501_dabfa0ef,
        64'h4501d3a5_85930000,
        64'h35974605_bf9101e5,
        64'h05130000_3517bfb9,
        64'h04050513_00003517,
        64'hc9192501_c96fb0ef,
        64'h54020808_f3f99cbd,
        64'h47b22860_10ef854e,
        64'hdbfff0ef_00044503,
        64'h9452dc9f_f0ef880d,
        64'h45210004_099b00c4,
        64'hd41be505_2501fedf,
        64'ha0ef0808_95ca6605,
        64'h00749181_02049593,
        64'h140a0a13_00003a17,
        64'h09620bf0_0913e12d,
        64'h44812501_e85fa0ef,
        64'h08080825_85930000,
        64'h35974605_d3afd0ef,
        64'h07050513_00003517,
        64'h80822701_01132401,
        64'h3a032481_39832501,
        64'h39032581_34832601,
        64'h34032681_3083d64f,
        64'hd0ef07a5_05130000,
        64'h3517c515_2501e75f,
        64'ha0ef2541_30232531,
        64'h34232521_38232491,
        64'h3c232681_30232611,
        64'h34239fa5_05130000,
        64'h4517e225_85930000,
        64'h35974605_d9010113,
        64'h8302037e_a9c58593,
        64'h00002597_4305f140,
        64'h25730ff0_000f0000,
        64'h100f8082_610560e2,
        64'he9fff0ef_00914503,
        64'hea7ff0ef_00814503,
        64'hf13ff0ef_ec06002c,
        64'h11018082_61456942,
        64'h64e27402_70a2fe94,
        64'h10e3ec9f_f0ef0091,
        64'h4503ed1f_f0ef3461,
        64'h00814503_f3fff0ef,
        64'h0ff57513_002c0089,
        64'h553354e1_03800413,
        64'h892af406_e84aec26,
        64'hf0227179_80826145,
        64'h694264e2_740270a2,
        64'hfe9410e3_f0bff0ef,
        64'h00914503_f13ff0ef,
        64'h34610081_4503f81f,
        64'hf0ef0ff5_7513002c,
        64'h0089553b_54e14461,
        64'h892af406_e84aec26,
        64'hf0227179_80826105,
        64'h644260e2_f43ff0ef,
        64'h00914503_f4bff0ef,
        64'h00814503_fb7ff0ef,
        64'h0ff47513_002cf5df,
        64'hf0ef0091_4503f65f,
        64'hf0ef0081_4503fd1f,
        64'hf0efec06_8121842a,
        64'h002ce822_11018082,
        64'h00f58023_00e580a3,
        64'h0007c783_00074703,
        64'h97aa973e_811100f5,
        64'h7713b7a7_87930000,
        64'h2797b7f5_0405fa5f,
        64'hf0ef8082_01416402,
        64'h60a2e509_00044503,
        64'h842ae406_e0221141,
        64'h808200e7_88230200,
        64'h071300e7_8423fc70,
        64'h071300e7_8623470d,
        64'h00078223_00e78023,
        64'h476d00e7_8623f800,
        64'h07130007_82231000,
        64'h07b78082_00a70023,
        64'hdfe50207_f7930147,
        64'h47831000_07378082,
        64'h02057513_0147c503,
        64'h100007b7_80820005,
        64'h45038082_00b50023,
        64'h80826105_690264a2,
        64'h644260e2_f47dfa1f,
        64'hf0ef4124_0433854a,
        64'h89260084_f3638922,
        64'h68048493_842ae04a,
        64'hec06e822_009894b7,
        64'he4261101_80826105,
        64'h690264a2_644260e2,
        64'hfe856ee3_f45ff0ef,
        64'h0405944a_02855433,
        64'h24040413_000f4437,
        64'h02a48533_370000ef,
        64'h892af63f_f0ef84aa,
        64'he04ae426_e822ec06,
        64'h11018082_02a7d533,
        64'h01419101_15026402,
        64'h60a202f4_07b32407,
        64'h8793000f_47b73a20,
        64'h00ef842a_f95ff0ef,
        64'he022e406_11418082,
        64'h610564a2_8d0502a7,
        64'hd5336442_60e29101,
        64'h150202f4_07b33e80,
        64'h07933ce0_00ef842a,
        64'hfc1ff0ef_84aae426,
        64'he822ec06_11018082,
        64'h45018082_01418d5d,
        64'h91011782_150260a2,
        64'h1007e783_10a7a223,
        64'h10e1a023_27051001,
        64'ha70300e5_7763878e,
        64'h1041e703_492000ef,
        64'he4061141_8082cf5f,
        64'hf06fa925_85930000,
        64'h45974611_cb81caa7,
        64'hd7830000_47978082,
        64'h24010113_22013903,
        64'h22813483_23013403,
        64'h23813083_f63ff0ef,
        64'h8522002c_ed4ff0ef,
        64'he802c44a_08282040,
        64'h061385a6_e92ff0ef,
        64'h22113c23_00282180,
        64'h06134581_893284ae,
        64'h842a2321_30232291,
        64'h34232281_3823dc01,
        64'h0113ebff_f06f6145,
        64'h05c170a2_41907402,
        64'hd8dff06f_614570a2,
        64'h65a27402_85228d5f,
        64'hd0efe42e_3b450513,
        64'h00003517_842a8e5f,
        64'hd06f6145_3dc50513,
        64'h00003517_70a27402,
        64'h02e78a63_470d00e7,
        64'h8e6301e1_578300f1,
        64'h0f230115_c78300f1,
        64'h0fa34709_0105c783,
        64'hf022f406_71798082,
        64'h61056902_64a26442,
        64'h60e2d61f_f06f6105,
        64'h690264a2_60e26442,
        64'h937fd0ef_3fc50513,
        64'h00003517_0087cf63,
        64'h278d439c_d9478793,
        64'h00004797_daf71023,
        64'h00004717_27850007,
        64'hd783dae7_87930000,
        64'h47972400_00ef0200,
        64'h0513d35f_f0ef4515,
        64'hdc45d583_00004597,
        64'h256000ef_4535e2df,
        64'hf0ef854a_bcc58593,
        64'h00004597_bca79b23,
        64'h00004797_4611d23f,
        64'hf0efdee5_55030000,
        64'h4517bea7_95230000,
        64'h4797d37f_f0ef4511,
        64'hdc3ff0ef_00448513,
        64'hffc4059b_06a79a63,
        64'h25010024_d783d53f,
        64'hf0efe1e5_55030000,
        64'h451708a7_95632501,
        64'h0004d783_d69ff0ef,
        64'h84ae450d_892a08c7,
        64'hdf638432_478de04a,
        64'he426ec06_e8221101,
        64'hb799e487_97230000,
        64'h4797eb1f_f0ef854e,
        64'hc5058593_00004597,
        64'h4611c4a7_9e230000,
        64'h4797da7f_f0ef4501,
        64'hc6a79423_00004797,
        64'hdb5ff0ef_e8f73623,
        64'h00004717_e8f73623,
        64'h00004717_451101f4,
        64'h17934405_a4bfd0ef,
        64'h4f050513_00003517,
        64'h858a4390_ea478793,
        64'h00004797_e22ff0ef,
        64'h850a85a2_e2aff0ef,
        64'h850a50a5_85930000,
        64'h359700f7_096302f0,
        64'h07930129_4703e1af,
        64'hf0ef850a_31458593,
        64'h00003597_893ff0ef,
        64'h850a4581_10000613,
        64'hb755eef7_25230000,
        64'h47172000_07938082,
        64'h615569b2_695264f2,
        64'h741270b2_abbfd0ef,
        64'h53850513_00003517,
        64'h00a405b3_f54ff0ef,
        64'h35850513_00003517,
        64'h842af62f_f0ef8522,
        64'h04a7f263_0ff00793,
        64'h9526f72f_f0ef3765,
        64'h05130000_351784aa,
        64'hf80ff0ef_8522f4a7,
        64'ha3230000_479704e7,
        64'hee631ff0_0793fff5,
        64'h071beabf_f0ef9526,
        64'h0505fa2f_f0ef8526,
        64'h00a404b3_0505faef,
        64'hf0ef892e_ea4aee26,
        64'hf6068522_89aae64e,
        64'h01258413_f2227169,
        64'h80824501_80820141,
        64'h640260a2_557d0085,
        64'h03638c0f_a0ef8432,
        64'he406e022_11418302,
        64'h61052501_05458593,
        64'h00002597_6902834a,
        64'h64a260e2_6442f140,
        64'h25730ff0_000f0000,
        64'h100fb81f_d0ef5e65,
        64'h05130000_35178622,
        64'h86aa608c_e77fc0ef,
        64'h85a26088_b9bfd0ef,
        64'h85a24124_043bec06,
        64'h5f050513_00003517,
        64'h0004b903_6380e04a,
        64'he82200a4_84930000,
        64'h449701a7_87930000,
        64'h4797e426_11018082,
        64'h610564a2_6442e00c,
        64'h95a660e2_600ca2ff,
        64'hf0efec06_600885aa,
        64'h84ae862e_e4260464,
        64'h04130000_4417e822,
        64'h11018082_04f73a23,
        64'h00004717_04f73a23,
        64'h00004717_07fe4785,
        64'h4e60006f_03050513,
        64'h014160a2_640202a4,
        64'h753b4529_fe7ff0ef,
        64'h357d02b4_55bb45a9,
        64'h00b7f863_47a500a0,
        64'h4563842e_e406e022,
        64'h1141bff9_0505fd07,
        64'h879b9fb9_02f587bb,
        64'h00d66763_0ff6f693,
        64'hfd07069b_8082853e,
        64'he3190005_470345a9,
        64'h46254781_80820141,
        64'h00e15503_00a10723,
        64'h812100a1_07a31141,
        64'hfa5ff06f_4581d7df,
        64'hf06f0141_05054581,
        64'h462960a2_6402f77d,
        64'h8b110007_4703973e,
        64'h00054703_fea47ae3,
        64'h157d8082_0141557d,
        64'h640260a2_e7198b11,
        64'h00074703_973efff5,
        64'h8513c227_87930000,
        64'h2797fff5_c70300a4,
        64'h05b395bf_f0efe589,
        64'h842ae406_e0221141,
        64'hbfd50789_bff1052a,
        64'h052ab7e9_e01c078d,
        64'h00e69863_04200713,
        64'h0027c683_fce69fe3,
        64'h052a0690_07130017,
        64'hc683fed7_16e306b0,
        64'h069302d7_076304d0,
        64'h06938082_01416402,
        64'h60a202d7_0e630470,
        64'h069300e6_ea6302d7,
        64'h04630007_c70304b0,
        64'h0693601c_f87ff0ef,
        64'h842ee406_e0221141,
        64'hb7e1e008_b7cdfc97,
        64'h879b0ff7_f793fe07,
        64'h079bc609_8a09b7d1,
        64'h96be0505_02d586b3,
        64'hfeb7f4e3_fd07879b,
        64'h00088b63_00467893,
        64'h80826105_85366442,
        64'h60e2ec05_00089863,
        64'h04467893_00064603,
        64'h00f80633_0007079b,
        64'h00054703_cfc80813,
        64'h00002817_468100c1,
        64'h6583e0ff_f0efc632,
        64'hec06006c_842ee822,
        64'h1101bfd5_0789bff1,
        64'h052a052a_b7e9e01c,
        64'h078d00e6_98630420,
        64'h07130027_c683fce6,
        64'h9fe3052a_06900713,
        64'h0017c683_fed716e3,
        64'h06b00693_02d70763,
        64'h04d00693_80820141,
        64'h640260a2_02d70e63,
        64'h04700693_00e6ea63,
        64'h02d70463_0007c703,
        64'h04b00693_601cf0df,
        64'hf0ef842e_e406e022,
        64'h11418082_014140a0,
        64'h053360a2_f23ff0ef,
        64'he4060505_1141f2df,
        64'hf06f00e6_846302d0,
        64'h07130005_4683b7e9,
        64'h4501e088_fcf718e3,
        64'h47a9fd27_9be30785,
        64'h8f81cb01_0007c703,
        64'hfe8782e3_67e2f5df,
        64'hf0ef8522_082c892a,
        64'h862e8082_61217902,
        64'h74a27442_70e25529,
        64'he90165a2_b0dff0ef,
        64'h84b2842a_e42e0006,
        64'h3023f04a_fc06f426,
        64'hf8227139_b7e1e008,
        64'hb7cdfc97_879b0ff7,
        64'hf793fe07_079bc609,
        64'h8a09b7d1_96be0505,
        64'h02d586b3_feb7f4e3,
        64'hfd07879b_00088b63,
        64'h00467893_80826105,
        64'h85366442_60e2ec05,
        64'h00089863_04467893,
        64'h00064603_00f80633,
        64'h0007079b_00054703,
        64'he5080813_00002817,
        64'h468100c1_6583f63f,
        64'hf0efc632_ec06006c,
        64'h842ee822_1101bf6d,
        64'h47a9bf7d_47a18082,
        64'h050900e7_93630780,
        64'h07130ff7_f7930207,
        64'h879bc709_8b050007,
        64'h4703973e_e9470713,
        64'h00002717_00154783,
        64'h02f71663_03000793,
        64'h00054703_02f71c63,
        64'h47c14198_c19c47c1,
        64'hc3b10447_f7930007,
        64'hc78397ba_00254703,
        64'h04d71b63_07800693,
        64'h0ff77713_0207071b,
        64'hc6898a85_0006c683,
        64'h00e786b3_ee478793,
        64'h00002797_00154703,
        64'h08f71163_03000793,
        64'h00054703_e7a9419c,
        64'hb7f1377d_87aabfa5,
        64'hfef51be3_0785f8b7,
        64'h12e30007_c70300d8,
        64'h0a630087_85130007,
        64'hb803bfcd_367d0785,
        64'hf8b71fe3_0007c703,
        64'hd24d8a1d_eb1187aa,
        64'h27018edd_00365713,
        64'h02079693_8fd90107,
        64'h179300b7_e7330085,
        64'h97938e1d_953e9381,
        64'h02071793_faf50785,
        64'h36fdfcb8_1ce30007,
        64'hc80387aa_0007069b,
        64'h40e7873b_47a1c31d,
        64'h00757713_b7f5367d,
        64'h0785feb7_1ce30007,
        64'hc7038082_853e4781,
        64'he60187aa_260100c7,
        64'hef630ff5_f59347c1,
        64'hb7ed853e_feb70be3,
        64'h00150793_00054703,
        64'h80824501_00c51463,
        64'h0ff5f593_962abfe9,
        64'h0405d175_f8bff0ef,
        64'h397d8522_85ce8626,
        64'h80826145_69a26942,
        64'h64e27402_70a28522,
        64'h44010099_5b630005,
        64'h091bd13f_f0ef8522,
        64'hc8890005_049bd1ff,
        64'hf0ef89ae_e84af406,
        64'he44eec26_852e842a,
        64'hf0227179_bfc50505,
        64'hfeb78de3_00054783,
        64'h808200c5_1363962a,
        64'hb7dd0585_0505fbed,
        64'h9f990005_c7030005,
        64'h47838082_853e4781,
        64'h00c51563_962ab7fd,
        64'h00f68023_16fd0005,
        64'hc78315fd_d7e500e5,
        64'h87b340b6_073300c5,
        64'h06b395b2_80820141,
        64'h640260a2_8522f57f,
        64'hf0ef00a5_e963842a,
        64'he406e022_11418082,
        64'h614564e2_69428526,
        64'h740270a2_00040023,
        64'hf79ff0ef_944a864a,
        64'h8522fff6_091300c5,
        64'h64636582_892ace11,
        64'h84aa6622_dcdff0ef,
        64'he02ee84a_f406e432,
        64'hec26852e_842af022,
        64'h7179bf65_fee78fa3,
        64'h0785fff5_c7030585,
        64'hbfe1469d_00c508b3,
        64'h87aa872e_bfc100e5,
        64'h07b3963e_95ba070e,
        64'h02f707b3_57e10036,
        64'h5713ff06_e8e340f8,
        64'h8833ff07_bc2307a1,
        64'hff873803_07218082,
        64'h02c79e63_963e87aa,
        64'hcb9d8b9d_00a5e7b3,
        64'h00b50a63_bf6dfeb7,
        64'h8fa30785_bfe1fef7,
        64'h3c230721_bfd10ff5,
        64'hf6934725_bfc1963a,
        64'h97aa078e_02e78733,
        64'h57610036_57930106,
        64'hef6340e8_8833469d,
        64'h00c508b3_872aff6d,
        64'h377d8fd5_07a28082,
        64'h04c79063_963e87aa,
        64'hcb9d0075_77938082,
        64'h4501b7e5_078900d7,
        64'h80a300e7_80238082,
        64'he3110017_c703ce81,
        64'h0007c683_87aacf99,
        64'h00054783_c11d8082,
        64'h610564a2_85266442,
        64'h60e2e008_05050005,
        64'h0023c501_f73ff0ef,
        64'h8526842a_c891e822,
        64'hec066104_e4261101,
        64'hbfd948a7_b9230000,
        64'h47970505_00050023,
        64'hc7810005_4783c519,
        64'hf9fff0ef_852285a6,
        64'h80826105_64a26442,
        64'h60e28522_44014a07,
        64'hbf230000_4797ef81,
        64'h00044783_942af9df,
        64'hf0ef85a6_8522cc11,
        64'h63804da7_87930000,
        64'h4797e519_842a84ae,
        64'hec06e426_e8221101,
        64'hbfd587ae_b7e50505,
        64'hfafd0007_c6830785,
        64'hfee68fe3_80824501,
        64'heb190005_4703bff9,
        64'h0785bfd5_872e8082,
        64'hfe081be3_00074803,
        64'h070500c8_0a638082,
        64'hea1140d7_85330007,
        64'hc60387aa_86aabfcd,
        64'h872eb7d5_0785fe08,
        64'h1be30007_48030705,
        64'hfed80fe3_8082ea99,
        64'h40c78533_0007c683,
        64'h87aa862a_b7fd0785,
        64'h808240a7_8533e701,
        64'h0007c703_00b78563,
        64'h87aa95aa_80826105,
        64'h644260e2_4501fe85,
        64'h7be3157d_00b78663,
        64'h00054783_0ff5f593,
        64'h952265a2_fe5ff0ef,
        64'hec06842a_e42ee822,
        64'h1101bfcd_07858082,
        64'h40a78533_e7010007,
        64'hc70387aa_bfcd0505,
        64'hdffd8082_00b79363,
        64'h00054783_0ff5f593,
        64'h80824501_bfcd0505,
        64'hc3998082_00b79363,
        64'h00054783_0ff5f593,
        64'h8082853e_ff790505,
        64'he3994187_d79b0187,
        64'h979b40f7_07bbfff5,
        64'hc7830005_47030585,
        64'ha8394781_00c59463,
        64'h962e8082_853ef37d,
        64'h0505e399_4187d79b,
        64'h0187979b_40f707bb,
        64'hfff5c783_00054703,
        64'h0585b7cd_87ba8082,
        64'h000780a3_00c71563,
        64'h8082e291_fed70fa3,
        64'h00178713_fff5c683,
        64'h0585963e_fb7d0017,
        64'h86930007_c70387b6,
        64'h8082e219_87aab7d5,
        64'h87b68082_fb75fee7,
        64'h8fa30785_fff5c703,
        64'h0585eb09_00178693,
        64'h0007c703_87aa8082,
        64'hfb65fee7_8fa30785,
        64'hfff5c703_058500c7,
        64'h896387aa_962a8082,
        64'hfb75fee7_8fa30785,
        64'hfff5c703_058587aa,
        64'h80820141_640260a2,
        64'h8d411502_9001fd1f,
        64'hf0ef1402_0005041b,
        64'hfdbff0ef_e022e406,
        64'h11418082_01412501,
        64'h640260a2_8d410105,
        64'h151bfe9f_f0ef842a,
        64'hfefff0ef_e022e406,
        64'h1141fc3f_f06f6de5,
        64'h05130000_45178082,
        64'h25018d5d_00f717bb,
        64'h40f007b3_00f7553b,
        64'h93ed836d_8f3d0127,
        64'hd713e118_97360017,
        64'h671302d7_86b36518,
        64'h6294611c_4b468693,
        64'h00004697_1180106f,
        64'h80826105_690264a2,
        64'h644260e2_8522e99f,
        64'hf0ef10f4_00230247,
        64'hc7838522_0ea42e23,
        64'h681c18f4_342320a7,
        64'h87930000_179718f4,
        64'h302321a7_87930000,
        64'h179716f4_3c2391c7,
        64'h8793ffff_f797e65f,
        64'hf0ef0405_28230325,
        64'h3023e904_10f502a3,
        64'h47850ef5_2c234799,
        64'hc57c57fd_cd21842a,
        64'h15c010ef_45051c00,
        64'h059384aa_892ec7ad,
        64'h639cc7bd_651ccbad,
        64'h511ccbbd_4d5ccfad,
        64'h44014d1c_c1414401,
        64'he04ae426_ec06e822,
        64'h1101b771_60002860,
        64'h10ef56a5_05130000,
        64'h351701a9_8863da4f,
        64'he0ef8566_85e20097,
        64'h8e63601c_db2fe0ef,
        64'h855e85ca_00090663,
        64'hdbefe0ef_638c855a,
        64'h0fc42603_681c8956,
        64'h0007c363_89524c1c,
        64'hc7914901_541cddcf,
        64'he06f6125_10c50513,
        64'h00004517_6d026ca2,
        64'h6c426be2_7b027aa2,
        64'h7a4279e2_690664a6,
        64'h60e66446_02941563,
        64'h4d295e2c_8c930000,
        64'h3c970005_0c1b04eb,
        64'h8b930000_4b9704eb,
        64'h0b130000_4b17046a,
        64'h8a930000_4a97056a,
        64'h0a130000_4a1789aa,
        64'he0caec86_e06ae466,
        64'he862ec5e_f05af456,
        64'hf852fc4e_6080e8a2,
        64'h86848493_00005497,
        64'he4a6711d_8082e308,
        64'he518e11c_e7886798,
        64'h88078793_00005797,
        64'he5088082_7007ae23,
        64'h00004797_e79ce39c,
        64'h89878793_00005797,
        64'hb7d56000_a9cff0ef,
        64'h8522c781_19a44783,
        64'h80826105_64a26442,
        64'h60e20094_176384be,
        64'hec06e426_6380e822,
        64'h8c878793_00005797,
        64'h11018082_43887667,
        64'h87930000_47978082,
        64'h0f850513_8082c398,
        64'h0015071b_438877e7,
        64'h87930000_4797bfd5,
        64'h55358082_610564a2,
        64'h644260e2_e0800f84,
        64'h0413e501_cf0ff0ef,
        64'h842acd09_f7dff0ef,
        64'h84aee822_ec06e426,
        64'h1101bfcd_f8400513,
        64'hbfe54501_80826105,
        64'h60e25535_eb3fe06f,
        64'h610560e2_00f70c63,
        64'h0ff00793_08154703,
        64'h02b70063_65a21035,
        64'h4703c105_fbdff0ef,
        64'he42eec06_11014148,
        64'h8082853e_bfd187b6,
        64'h00a60463_0fc7a603,
        64'h80820141_853e4781,
        64'h60a2f60f_e0efe406,
        64'h16850513_00004517,
        64'h85aa1141_02e79063,
        64'h6394631c_99470713,
        64'h00005717_80824501,
        64'h80820141_45016402,
        64'h60a20dc0_00ef13e0,
        64'h00ef02c0_0513fc5f,
        64'hf0ef8522_00055563,
        64'haeefe0ef_852212a0,
        64'h00ef9cf7_23230000,
        64'h5717842a_e406e022,
        64'h47851141_ef9d439c,
        64'h9dc78793_00005797,
        64'h808218b5_0d238082,
        64'h557d8082_557d8082,
        64'h4501c56c_e54ff06f,
        64'hfa100413_f0eff06f,
        64'h2006061b_40010637,
        64'hf0a60963_4505f0c5,
        64'h43638ca6_02e34509,
        64'h8a3d01a6_d61bf2c5,
        64'h1a634000_063706bb,
        64'ha42306eb_a22306fb,
        64'ha02304db_ae23018b,
        64'ha50345e6_475647c6,
        64'h46b6ea05_1163842a,
        64'h93bfe0ef_c4be855e,
        64'h0107979b_008c4601,
        64'h07cbd783_c2be479d,
        64'h04f11023_47a506fb,
        64'h9e2304e1_57830007,
        64'hd663018b_a783ec05,
        64'h1b63842a_96ffe0ef,
        64'hc2be47d5_855ec4be,
        64'h0107979b_008c4601,
        64'h07cbd783_04f11023,
        64'h478d6da0_00ef06cb,
        64'h851300ec_4641bf6d,
        64'h11872583_974e8379,
        64'h02079713_fcfc65e3,
        64'h4581b7c9_f521d31f,
        64'he0ef855e_45850b70,
        64'h06130ff6_f693bb91,
        64'hfd319fdf_e0ef855e,
        64'hcb0ff0ef_855e4601,
        64'h18fbae23_08bba223,
        64'h0017b793_17ed088b,
        64'ha583ef8d_1afba823,
        64'h409ce79d_0046f793,
        64'h00892683_f941808f,
        64'hf0ef855e_408c933f,
        64'he0ef855e_02ebaa23,
        64'h0017b713_41b787b3,
        64'h01a78663_471100d7,
        64'h89634721_400006b7,
        64'h00092783_bb6d925f,
        64'he0ef1ba5_05130000,
        64'h4517f764_9fe304a1,
        64'hfb9911e3_0931973f,
        64'he0ef855e_035baa23,
        64'h08fba223_180bae23,
        64'h1a0ba823_088ba783,
        64'hddbfe0ef_855e4585,
        64'h0b700613_4681c131,
        64'hdebfe0ef_855e0fb6,
        64'hf6934585_0b700613,
        64'h00894683_c3a18ff9,
        64'h00fa77b3_00092703,
        64'h40dc04f7_18630017,
        64'hb79317ed_00494703,
        64'h409c1000_0db72000,
        64'h0d37d8a9_09130000,
        64'h3917cbb5_278100fa,
        64'h77b300fa_97bb409c,
        64'hddcc8c93_00003c97,
        64'h4c2ddaab_0b130000,
        64'h3b174a85_db4ff0ef,
        64'hd9848493_00003497,
        64'h00fa7a33_855e4601,
        64'h088ba583_044ba783,
        64'h040baa03_04fba023,
        64'h00c7e793_040ba783,
        64'hc7998b85_04eba023,
        64'h01076713_040ba703,
        64'h04eba023_0217071b,
        64'hc68900c7_f693ce91,
        64'h0027f693_1adba423,
        64'h03f7f693_0c46c783,
        64'h04fba023_0017079b,
        64'h70000737_bb952e65,
        64'h05130000_4517e691,
        64'hecf76ce3_1a0bb683,
        64'h400407b7_04fba023,
        64'h27851000_07b7b8d1,
        64'h02fba423_47857400,
        64'h10ef8526_a3ffe0ef,
        64'h8a3d8abd_0146561b,
        64'h0106569b_06248513,
        64'h36858593_00004597,
        64'h074ba603_a5ffe0ef,
        64'h04d48513_36c58593,
        64'h00004597_26810ff7,
        64'h77130ff8_78130ff7,
        64'hf7930188_569b0108,
        64'h571b0088_579b06cb,
        64'hc603077b_c883070b,
        64'ha803a95f_e0effef5,
        64'h36230245_051338e5,
        64'h85930000_459784aa,
        64'h06fbc603_074bd683,
        64'h07abd703_02c7d7b3,
        64'hed109201_0a8bb783,
        64'hd11c9fb9_071200e0,
        64'h37338f75_02071613,
        64'h76c19fb5_068e00d0,
        64'h36b38ef9_f0068693,
        64'hff0106b7_9fb5068a,
        64'h00d036b3_8ef90f06,
        64'h8693f0f0_f6b79fb5,
        64'h00f037b3_068600d0,
        64'h36b32781_8ef98ff9,
        64'hccc68693_aaa78793,
        64'hccccd6b7_aaaab7b7,
        64'h08cba703_00050623,
        64'h00051523_484000ef,
        64'h855e08fb_a82308fb,
        64'ha6232000_0793c799,
        64'h19cba783_1afbaa23,
        64'h1b0ba783_0adba223,
        64'h0afba023_02d606bb,
        64'h02f757bb_8a8d0106,
        64'hd69b02e6_073b3e80,
        64'h0613c305_c38d03f7,
        64'h77132781_0126d71b,
        64'h8fd10186_d61b8ff9,
        64'h17fd67c1_00cca683,
        64'h08fbae23_0087171b,
        64'h1487a783_97b6078a,
        64'hee868693_00003697,
        64'h04d61c63_800306b7,
        64'h018ba603_00f6f863,
        64'h8bbd00c7_579b46a5,
        64'h008ca703_fdb59ee3,
        64'hfefdae23_8fd98ff5,
        64'h8f510087_d79b8e69,
        64'h0087961b_8f510187,
        64'h971b0187_d61b0d91,
        64'h000da783_f0068693,
        64'h00ff0537_040d8593,
        64'h66c1b545_11872583,
        64'h974e8379_02079713,
        64'heaf768e3_4581472d,
        64'hb35d04fb_a0230087,
        64'h6793da06_d9e3040b,
        64'ha70302e7_96938fd1,
        64'h8ff50087_d79b0087,
        64'h961bf006_869366c1,
        64'h44dcfbe1_8b8583a5,
        64'h4cdcd005_1ce3d61f,
        64'he0efdc3e_f84af426,
        64'hc556855e_010c0400,
        64'h07931030_c33e47d5,
        64'h08f11023_4799020a,
        64'h08633a7d_09053ac5,
        64'h4a159881_19020100,
        64'h0ab70ff1_04934905,
        64'hbbc58003_0737de07,
        64'h5ee30307_971300eb,
        64'hac238002_0737b519,
        64'ha007071b_80011737,
        64'hb61ddf40_0413cbdf,
        64'he0ef5525_05130000,
        64'h4517e6f4_9fe30967,
        64'h87930000_379704a1,
        64'heafa94e3_47a10a91,
        64'h8c9ff0ef_855e8405,
        64'h85934601_180bae23,
        64'h096ba223_1afba823,
        64'h017d85b7_4785f3ed,
        64'h37fd6702_67a20e05,
        64'h0c63e0df_e0efe03a,
        64'hc93ae552_e16ee43e,
        64'h855e110c_01100400,
        64'h07134791_d502d33a,
        64'h0af11023_47b56702,
        64'he915e35f_e0efd53e,
        64'he03ad33a_8cee855e,
        64'h110c0107_979b4601,
        64'h475507cb_d7830af1,
        64'h10230370_0793fe07,
        64'hfd930ff1_0793947f,
        64'hf0ef855e_460118fb,
        64'hae2308bb_a2230017,
        64'hb79317ed_088ba583,
        64'h14079a63_1afba823,
        64'h409c09b7_94638bbd,
        64'h010c4783_e941e91f,
        64'he0efc93e_e552e162,
        64'h855e110c_04000793,
        64'h0110d53e_00fde7b3,
        64'h17c12d81_810007b7,
        64'hd33e47d5_0af11023,
        64'h47994d85_0ce79163,
        64'h470d01a7_8663409c,
        64'hdfdfe0ef_855e02fb,
        64'haa23001c_b79340fc,
        64'h8cb31000_07b700ec,
        64'h88634791_20000737,
        64'h00ec8d63_47a14000,
        64'h07370e05_1c638daa,
        64'h971ff0ef_855e0015,
        64'hb59340bc_85b31000,
        64'h05b700fc_88634591,
        64'h200007b7_00fc8d63,
        64'h45a14000_07b71407,
        64'h81630197_f7b300f9,
        64'h77b340dc_0007ac83,
        64'h97d6109c_840b0b1b,
        64'h4a81017d_8b371607,
        64'h85632781_00f977b3,
        64'h00e797bb_47854098,
        64'h0a05fe07_fc1383f9,
        64'h79130ff1_079300f9,
        64'h793321a4_84930000,
        64'h3497020d_1a13044b,
        64'ha783f0be_4d05040b,
        64'ha903639c_e3c78793,
        64'h00005797_1ef71863,
        64'h800107b7_018ba703,
        64'h04fba023_8fd92000,
        64'h0737040b_a7830007,
        64'h596302d7_971300eb,
        64'hac238001_073720d7,
        64'h02634689_21270063,
        64'h8b3d0187_d71b04eb,
        64'hac238f55_8f718ecd,
        64'h0087571b_8de90087,
        64'h159b8ecd_0187169b,
        64'h0187559b_40d804fb,
        64'haa232781_8fd58ef1,
        64'hf0070613_8fd16741,
        64'h0087569b_8e698fd5,
        64'h0087161b_0187179b,
        64'h0187569b_00ff0537,
        64'h4098b555_8b1d9381,
        64'h00f7571b_17828fd5,
        64'h01e7569b_8ff50027,
        64'h979b16f1_6685b54d,
        64'h08bba823_00b515bb,
        64'h89bd0165_d59bbd99,
        64'h40030637_a7a94002,
        64'h0637bb45_842afe0a,
        64'h16e33a7d_c131850f,
        64'hf0efd05a_ec56e826,
        64'h855e108c_08104b21,
        64'h0a854a11_d48206f1,
        64'h10239881_02091a93,
        64'h03300793_0bf10493,
        64'h4905d2ca_ed05880f,
        64'hf0efd4be_d2ca855e,
        64'h0107979b_108c4601,
        64'h07cbd783_06f11023,
        64'h03700793_04fba023,
        64'h27891000_07b75407,
        64'h5a63018b_a703e005,
        64'h1fe3842a_ffbfe0ef,
        64'h855e00b5_45830f70,
        64'h00ef855e_e2051ae3,
        64'h842ac9af_f0ef855e,
        64'h08fb80a3_57fd08fb,
        64'haa234785_e40516e3,
        64'h842a8e4f_f0efc4be,
        64'hc2ca855e_008c0107,
        64'h979b4601_495507cb,
        64'hd78304f1_1023479d,
        64'h902ff0ef_c282c4be,
        64'h04e11023_855e008c,
        64'h46010107_979b4711,
        64'h00e78e63_577d04cb,
        64'ha783c215_08fba823,
        64'h00e7f463_20000793,
        64'h090ba703_08fba623,
        64'h0107d463_20000793,
        64'h0afbb823_0e0bb023,
        64'h0c0bbc23_0c0bb823,
        64'h0c0bb423_0c0bb023,
        64'h0a0bbc23_030787b3,
        64'h00e797b3_07090785,
        64'h47219381_17828fd9,
        64'h8ff50107_571b003f,
        64'h06b70107_979b1406,
        64'h8e6302cb_a683090b,
        64'ha8231408_dc63090b,
        64'ha62300d5_183b8abd,
        64'h0107d69b_08dba223,
        64'h08dba423_04cba823,
        64'h180bae23_1a0ba823,
        64'h8a0500c7_d61b02d6,
        64'h06bb018b_a8834505,
        64'h1086a683_0f864603,
        64'h96ce964e_068a8a3d,
        64'h40098993_00003997,
        64'h8a9d0036_d61b00cb,
        64'hac234006_061b4001,
        64'h0637a029_40040637,
        64'h0ea61ee3_45111aa6,
        64'h0f63450d_bf0506fb,
        64'h9e234785_02fba623,
        64'h8b8541e7_d79b048b,
        64'ha78300fb_ac234000,
        64'h07b7bfe9_1a5010ef,
        64'h06400513_12a96ee3,
        64'h117010ef_85260007,
        64'hcc63048b_a783f155,
        64'h842ab36f_f0ef855e,
        64'h45853e80_09139081,
        64'h02051493_13b010ef,
        64'h4501b16f_f0ef855e,
        64'h0407c163_180b8c23,
        64'h048ba783_8082615d,
        64'h6db66d56_6cf67c16,
        64'h7bb67b56_7af66a1a,
        64'h69ba695a_64fa741a,
        64'h70ba8522_d55d842a,
        64'hd99ff0ef_855ea031,
        64'h020ba423_f4fd34fd,
        64'h100503e3_842aaa0f,
        64'hf0ef855e_008c4601,
        64'h4495cf81_8b851b8b,
        64'ha7831205_00e3842a,
        64'habaff0ef_c482c2be,
        64'h855e008c_479d4601,
        64'h04f11023_4789e7b5,
        64'h180b8ca3_198bc783,
        64'hc7b1199b_c7831cd0,
        64'h10ef4501_8baae3b5,
        64'h4401e6ee_eaeaeee6,
        64'hf2e2f6de_fadafed6,
        64'he352e74e_eb4aef26,
        64'hf706f322_7161551c,
        64'hb58584aa_b595fa10,
        64'h0493a10f_f0efa765,
        64'h05130000_5517d965,
        64'hc1cff0ef_85224585,
        64'hbfd118f4_0c234785,
        64'h0007d663_443ced09,
        64'hc34ff0ef_85224581,
        64'hc04ff0ef_852202f5,
        64'h1f63f920_0793b55d,
        64'h18f40ca3_47850604,
        64'h1e23d45c_8b8541e7,
        64'hd79bc43c_cc188001,
        64'h073700e6_85638002,
        64'h07374c14_bf452ff0,
        64'h10ef3e80_05130609,
        64'h0863397d_0007ca63,
        64'h47b2ed1d_b8eff0ef,
        64'h8522858a_4601c43e,
        64'h0197e7b3_01871563,
        64'hc43e0177_f7b3c25a,
        64'h4bdc0151_10234c18,
        64'h681ce13d_bb6ff0ef,
        64'hc402c252_01311023,
        64'h8522858a_46014000,
        64'h0cb78002_0c3700ff,
        64'h8bb74b05_02900a93,
        64'h4a550370_09933e90,
        64'h0913cc1c_800207b7,
        64'h00f71563_0aa00793,
        64'h00c14703_e911bf8f,
        64'hf0efc23e_c43a8522,
        64'h858a4601_47d50aa0,
        64'h0713e399_1aa00713,
        64'h8ff94bdc_00ff8737,
        64'h681c00f1_102347a1,
        64'h000505a3_45d000ef,
        64'h8522f149_84aacf2f,
        64'hf0ef8522_f1dff0ef,
        64'h85224581_4601b72f,
        64'hf0ef8522_d85c4785,
        64'h08f42223_1a042823,
        64'h18042e23_08842783,
        64'hf94584aa_97826b9c,
        64'h679c8522_681c3ef0,
        64'h10ef7d00_0513ba2f,
        64'hf0ef8522_02042c23,
        64'h02f40823_47851af4,
        64'h2c23478d_f93ff0ef,
        64'hf3e54481_541c8082,
        64'h61097ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h74a67906_85267446,
        64'h70e6f850_0493bacf,
        64'hf0efbfa5_05130000,
        64'h55170204_2423eb8d,
        64'h6b9c679c_681cc509,
        64'hf11ff0ef_842ac17c,
        64'h8fd9f466_f862fc5e,
        64'he0dae4d6_e8d2ecce,
        64'hf0caf4a6_fc86f8a2,
        64'h070d4b9c_71191000,
        64'h0737691c_80828082,
        64'hc2cff06f_02c50823,
        64'hdd0c0007_059b00e7,
        64'hf46385be_27814f18,
        64'h87ae00f5_f3634f5c,
        64'h6918ee09_b7cdc402,
        64'hfef414e3_47858082,
        64'h61217902_74a27442,
        64'h70e2d34f_f0ef8526,
        64'h858a4601_c43e4789,
        64'h00f41f63_4791c24a,
        64'h00f11023_4799ed19,
        64'hd52ff0ef_c43ec24a,
        64'h8526858a_46010107,
        64'h979b4955_842e07c4,
        64'hd78300f1_10230370,
        64'h079304f5_92635529,
        64'h478500f5_866384aa,
        64'h4791f04a_f822fc06,
        64'hf4267139_80820141,
        64'h640260a2_45058302,
        64'h014160a2_64028522,
        64'h00030763_0187b303,
        64'h679c681c_00055e63,
        64'h810ff0ef_842ae406,
        64'he0221141_b32ddd79,
        64'h842a945f_f0ef854a,
        64'h45850a70_061386ce,
        64'hbb3d842a_957ff0ef,
        64'h854a4585_09b00613,
        64'h46850137_9b630a7a,
        64'h4783d4fb_0de34785,
        64'hed19975f_f0ef854a,
        64'h458509c0_061386de,
        64'hfdb498e3_0c110ff4,
        64'hf493248d_ffac90e3,
        64'h0ffafa93_2ca12a85,
        64'he13999df_f0ef854a,
        64'h0ff6f693_0196d6bb,
        64'h45858656_000c2683,
        64'h4c818aa6_09b00d93,
        64'h4d61ffa4_92e32ca1,
        64'h0ff4f493_2485e935,
        64'h9cbff0ef_854a4585,
        64'h86260ff6_f693019a,
        64'hd6bb08f0_0d134c81,
        64'hffb492e3_2d210ff4,
        64'hf4932485_ed499f1f,
        64'hf0ef854a_45858626,
        64'h0ff6f693_01acd6bb,
        64'h08c00d93_4d010880,
        64'h049308f9_2a2300a7,
        64'h979b0e0a_47830afa,
        64'h07a34785_e569a21f,
        64'hf0ef854a_45850af0,
        64'h06134685_e3958b85,
        64'h0afa4783_e20b02e3,
        64'hb51d547d_dbaff0ef,
        64'hde850513_00005517,
        64'hcb898b85_09ba4783,
        64'hbfd100f9_f9b3fff7,
        64'hc793b591_2cc020ef,
        64'hdb850513_00005517,
        64'hef898b85_0a6a4783,
        64'h02d98263_fcc592e3,
        64'h872e0ff9_f99300f9,
        64'he9b3c70d_4189d99b,
        64'h4187d79b_8b050189,
        64'h999b0187_979b0027,
        64'h571b00b5_17bb0208,
        64'h04630018_78130017,
        64'h581b4b18_9726070e,
        64'h0017059b_46114505,
        64'h47010016_e993c399,
        64'h0fe6f993_8b89c719,
        64'h89b60017_f7130a7a,
        64'h46830084_c783b5c1,
        64'he56ff0ef_e0450513,
        64'h00005517_85ce0136,
        64'h7a63963e_09da4783,
        64'h9e3d0087_979b0106,
        64'h161b09ea_478309fa,
        64'h4603ee05_19e3842a,
        64'hf94ff0ef_854a85d2,
        64'hfe0a7a13_02f10a13,
        64'hf00600e3_e1450513,
        64'h00005517_8a09000b,
        64'h8963fbc5_96e387ae,
        64'h05110821_013309bb,
        64'h0ffbfb93_00dbebb3,
        64'h00be96bb_cb898b85,
        64'h0107c783_97a6078e,
        64'h02088063_00652023,
        64'h02e8d33b_b7f14b81,
        64'h4a814c81_b7c1ee4f,
        64'hf0efe325_05130000,
        64'h55170003_0d6302e8,
        64'hf33b0017_859b0008,
        64'h28834e11_4e854781,
        64'h89d68562_00c48813,
        64'h8c0a009c_9c9be399,
        64'h4b8502ea_dabb02c9,
        64'h2783bf41_5429f24f,
        64'hf0efe3a5_05130000,
        64'h5517cb89_02ecf7bb,
        64'h0005ac83_e79102ea,
        64'hf7bb060a_81630045,
        64'haa83db45_e3450513,
        64'h00005517_09892703,
        64'h80822a01_01132381,
        64'h3d832401_3d032481,
        64'h3c832501_3c032581,
        64'h3b832601_3b032681,
        64'h3a832701_3a032781,
        64'h39832801_39032881,
        64'h34832901_34032981,
        64'h30838522_f8400413,
        64'hf96ff0ef_e5c50513,
        64'h00005517_e7b90016,
        64'h779307e9_460300e7,
        64'heb63e3a5_05130000,
        64'h551784ae_8b32892a,
        64'hbfe78793_3ffc07b7,
        64'h9f3dbff7_879bbffc,
        64'h07b74d18_0ac7e963,
        64'h478923b1_3c2325a1,
        64'h30232591_34232581,
        64'h38232571_3c232761,
        64'h30232751_34232741,
        64'h38232731_3c232921,
        64'h30232891_34232881,
        64'h38232811_3c23d601,
        64'h01138082_614569a2,
        64'h694264e2_740270a2,
        64'h85220135_05a315e0,
        64'h10ef8526_842a875f,
        64'hf0ef8526_85ca0009,
        64'h1c6300f5_1e63842a,
        64'h57b5c519_cc7ff0ef,
        64'h84aa4585_0b300613,
        64'h8edd892e_9be10079,
        64'hf6930ff5_f9930815,
        64'h4783f022_f406e44e,
        64'he84aec26_7179b74d,
        64'h84aab75d_df400493,
        64'hf7d50b94_4783e519,
        64'h98dff0ef_854a85a2,
        64'h980101f1_0413f1e9,
        64'h258199f5_ffe4059b,
        64'hf57184aa_d1fff0ef,
        64'h892a4585_0b900613,
        64'h842e4685_fef760e3,
        64'h4705ffc5_879b8082,
        64'h24010113_22813483,
        64'h22013903_85262301,
        64'h34032381_308354a9,
        64'hc5854681_02b7e163,
        64'h02f58863_47892321,
        64'h30232291_34232281,
        64'h38232211_3c23dc01,
        64'h0113bf45_5929bf55,
        64'h5951bf65_1a04b023,
        64'h524020ef_d1691a04,
        64'hb503892a_bf4d08f4,
        64'haa2302f7_07bb2785,
        64'h27058bfd_8b7d0057,
        64'hd79b00a7_d71b50fc,
        64'h80822501_01132281,
        64'h39832301_39032381,
        64'h3483854a_24013403,
        64'h24813083_08f48023,
        64'h0a744783_08d4ac23,
        64'h02f686bb_00a6969b,
        64'h0dd44783_f8dc07a6,
        64'h0d442783_00098663,
        64'hc79954dc_08f4aa23,
        64'h00a6979b_c7b98b85,
        64'h0e044683_0af44783,
        64'h0af407a3_4785ed35,
        64'he0bff0ef_85264585,
        64'h0af00613_4685ce81,
        64'he3918bfd_09c44783,
        64'hc7898b85_0a044783,
        64'hf4fc07a6_c319f4fc,
        64'h54d89fb9_08844703,
        64'h9fb90087_171b0894,
        64'h47039fb9_0107171b,
        64'h0187979b_08a44703,
        64'h08b44783_f8fc07ce,
        64'h02e787b3_0dd44783,
        64'h02f70733_0e044703,
        64'h97ba08c4_47039fb9,
        64'h0087171b_0107979b,
        64'h468508d4_470308e4,
        64'h47830409_8f63fca7,
        64'h14e30621_070de21c,
        64'h07ce02b7_87b30dd4,
        64'h478302f5_85b30e04,
        64'h45830009_8c634685,
        64'hc39197ae_ffe74583,
        64'h9fad0105_959b0087,
        64'h979b0007_4583fff7,
        64'h4783e0fc_07c64681,
        64'h09d40513_0a844783,
        64'hfcdc07c6_0c848613,
        64'h09140713_0e244783,
        64'h06f48fa3_09c44783,
        64'hc7898b89_0a044783,
        64'h00098a63_08f480a3,
        64'h0b344783_c7890e24,
        64'h4783e781_0019f993,
        64'h8b8506f4_8f2309b4,
        64'h49830a04_4783f8dc,
        64'h00d77363_0147d693,
        64'h07a68007_07136705,
        64'h0d442783_00e7fd63,
        64'hcc981ff7_87934004,
        64'h07b753b8_97ba078a,
        64'hdf070713_00004717,
        64'h1cf76b63_47210c04,
        64'h47831230_10ef85a2,
        64'h20000613_1e050363,
        64'h1a04b503_1aa4b023,
        64'h6c2020ef_20000513,
        64'he7991a04_b7831e05,
        64'h1863892a_c09ff0ef,
        64'h84aa85a2_980101f1,
        64'h04131ce7_f5634901,
        64'h3ffc0737_23313423,
        64'h22913c23_24813023,
        64'h24113423_9fb92321,
        64'h3823bffc_07b7db01,
        64'h01134d18_bfcdfc79,
        64'h347d8082_612174a2,
        64'h744270e2_d91ff0ef,
        64'h85263e80_0593e919,
        64'hc53ff0ef_8526858a,
        64'h4601440d_c43684aa,
        64'hfc06f426_f8228ed1,
        64'h0106161b_8edd0300,
        64'h07b70086_969bc23e,
        64'h47f500f1_10234799,
        64'h71398082_61216aa2,
        64'h6a4269e2_74a27902,
        64'h85267442_70e2fc09,
        64'h99e39aa2_02878433,
        64'h9a224089_89b308c9,
        64'h6783fc85_1ae3f01f,
        64'hf0ef854a_85d68652,
        64'h86a2844e_0089f363,
        64'h0207e403_01093783,
        64'h89a6f96d_ecdff0ef,
        64'h854a08c9_2583a089,
        64'h4481bd9f_f0ef2365,
        64'h05130000_551700b6,
        64'h7a630144_85b36810,
        64'h00054d63_8c5fa0ef,
        64'h852200b4_4583c11d,
        64'h892a4820_10ef8ab6,
        64'h84b28a2e_4148842a,
        64'hce05e456_e852ec4e,
        64'hf04af426_f822fc06,
        64'h7139b7c5_4401b7d5,
        64'h0004841b_b74d02f6,
        64'h063bbf61_47c58082,
        64'h61256906_64a66446,
        64'h60e68522_c43ff0ef,
        64'h28050513_00005517,
        64'hc11dd55f_f0efd23e,
        64'hd402854a_100c47f5,
        64'h460102f1_102347b1,
        64'h0497f063_4785e529,
        64'h842ad75f_f0efc83e,
        64'hca26d23a_854a100c,
        64'h47850030_cc3ee42e,
        64'h4755d432_cf3108c9,
        64'h27832601_02f11023,
        64'h02c92703_47c906d7,
        64'hf66384b6_892a4785,
        64'he8a2ec86_e0cae4a6,
        64'h711d8082_4501bfd5,
        64'h45018082_612174a2,
        64'h744270e2_f8ed34fd,
        64'hc901dcdf_f0ef8522,
        64'h858a4601_4495cb91,
        64'h8b891b84_2783c11d,
        64'hde3ff0ef_c23e842a,
        64'hf426fc06_f822858a,
        64'h460147d5_c42e00f1,
        64'h102347c1_7139e7a9,
        64'h19c52783_bf7df920,
        64'h0513d09f_f0ef3265,
        64'h05130000_5517fc80,
        64'h49e34501_b7555a60,
        64'h20ef3e80_051300f0,
        64'h57630014_079b347d,
        64'hfe04c6e3_34fd8082,
        64'h61257aa2_7a4279e2,
        64'h690664a6_644660e6,
        64'hfba00513_d4bff0ef,
        64'h35050513_00005517,
        64'hc78d0125_f7b30547,
        64'h93630135_f7b3c789,
        64'h1005f793_45b2ed0d,
        64'he73ff0ef_8556858a,
        64'h4601e00a_0a13e009,
        64'h89930809_09134495,
        64'hc43e842e_8aaaec86,
        64'hf456e4a6_e8a26a05,
        64'h6989fdf9_49370107,
        64'h979bf852_fc4ee0ca,
        64'h07c55783_c23e47d5,
        64'h00f11023_47b5711d,
        64'h80826145_740270a2,
        64'hc43c47b2_e119ec9f,
        64'hf0ef8522_858a4601,
        64'hc43e8fd9_8f554000,
        64'h06b78f75_600006b7,
        64'h8ff58ff9_f8078793,
        64'h4ad40080_07b74538,
        64'h6914c195_842ac402,
        64'hc23ef406_f0224785,
        64'h00f11023_47857179,
        64'h80826145_740270a2,
        64'h852269a0_20ef7d00,
        64'h0513e509_842af21f,
        64'hf0efc202_c4020001,
        64'h1023858a_46018522,
        64'h6b8020ef_f4063e80,
        64'h0513842a_f0227179,
        64'hb761fb60_0513d551,
        64'h56f010ef_0d448513,
        64'h0d440593_461100f7,
        64'h1a630e04_47830e04,
        64'hc70302f7_10630c04,
        64'h47830c04_c70302f7,
        64'h16630dd4_47830dd4,
        64'hc70302f7_1c630a04,
        64'h47830a04_c703f579,
        64'hf95ff0ef_1a053483,
        64'h22113c23_22913423,
        64'h85a29801_01f10413,
        64'h22813823_dc010113,
        64'h80822401_01132281,
        64'h34832301_34032381,
        64'h30834501_80824501,
        64'h00e6fe63_40040737,
        64'h4d148082_616160a6,
        64'hfd3ff0ef_cc3ed402,
        64'he486100c_20000793,
        64'h0030e83e_e42e0785,
        64'h17824785_d23e47d5,
        64'h02f11023_47a1715d,
        64'h83020007_b303679c,
        64'h691c8082_4f450513,
        64'h00005517_80826108,
        64'h953e8175_24478793,
        64'h00004797_150200a7,
        64'heb6347ad_8082557d,
        64'h80820141_640260a2,
        64'h45018302_014160a2,
        64'h64028522_00030763,
        64'h0207b303_679c681c,
        64'h00055e63_ff5ff0ef,
        64'h842ae406_e0221141,
        64'h8082557d_8082557d,
        64'hb7e9659c_95aa058e,
        64'h05e135f1_bfd9617c,
        64'hbfe97d5c_80826105,
        64'h4501e91c_64a26442,
        64'h60e202f4_57b39381,
        64'h02049793_0c5010ef,
        64'h7540f55c_08c52483,
        64'h795c8782_97bae426,
        64'he822ec06_1101439c,
        64'h97ba83f9_2bc70713,
        64'h00004717_02059793,
        64'h04b7ee63_479d8082,
        64'h45018302_00030363,
        64'h0087b303_679c691c,
        64'h80826135_645260f2,
        64'h85220f70_20ef0808,
        64'h842ae3ff_f0efe436,
        64'heec6eac2_e6bee2ba,
        64'hea22ee06_08081000,
        64'h05931234_862afe36,
        64'hfa32f62e_710d8082,
        64'h616160e2_e69ff0ef,
        64'he436e4c6_e0c2fc3e,
        64'hf83aec06_10000593,
        64'h1014862e_f436f032,
        64'h715d8082_616160e2,
        64'he8dff0ef_e436e4c6,
        64'he0c2fc3e_f83aec06,
        64'h1034f436_715db7f1,
        64'h85220201_03930005,
        64'h059b4db0_10ef8522,
        64'h01247433_60000084,
        64'h0b13b5fd_845ad93f,
        64'hf0ef0084_0b130201,
        64'h03930004_4503a809,
        64'hddbff0ef_00280201,
        64'h03930005_059be37f,
        64'hf0ef4008_45a94601,
        64'h0016b693_00380084,
        64'h0b13f8b5_0693a811,
        64'h45c10016_36134685,
        64'h00380084_0b13fa85,
        64'h0613f6e5_10e30780,
        64'h071302e5_00630750,
        64'h0713a00d_46014685,
        64'h00380084_0b13f6e5,
        64'h1ee30700_071300a7,
        64'h6c6306e5_0e630730,
        64'h0713b74d_048d0024,
        64'hc5038082_61090007,
        64'h051b6b06_6aa66a46,
        64'h69e67906_74a67446,
        64'h70e6f55d_08f50963,
        64'h06300793_04d50f63,
        64'h05800693_02a6eb63,
        64'h06d50f63_06400693,
        64'h04890014_c5034781,
        64'h00f6f363_46a50ff7,
        64'hf793fd07_879bcb9d,
        64'h0004c783_03551063,
        64'h47810489_05450f63,
        64'h0014c503_bfe1e7bf,
        64'hf0ef0201_03930485,
        64'h01350863_04d7ff63,
        64'h93811782_76820017,
        64'h079bc52d_8f1d0004,
        64'hc50377a2_77420209,
        64'h59130300_0a9306c0,
        64'h0a130250_0993f82a,
        64'hf02ef42a_fc3e8436,
        64'h84b2e0da_fc86e4d6,
        64'he8d2ecce_f4a6f8a2,
        64'h597d011c_f0ca7119,
        64'hb7f10685_01178023,
        64'h00668023_26050006,
        64'hc8830007_c30397ba,
        64'h93811782_40c807bb,
        64'hb7d92585_fea68fa3,
        64'h0685bf5d_00a8053b,
        64'h808200b6_1b63fff5,
        64'h081b86ba_25810006,
        64'h80230015_559b40e6,
        64'h853b0685_00f68023,
        64'h02d00793_00088763,
        64'h02f5e963_03000513,
        64'h40e685bb_fe718532,
        64'hfea68fa3_06850ff5,
        64'h751302b6_563b0305,
        64'h051b046e_67630ff3,
        64'h751302b6_733b0005,
        64'h061b3859_86ba4e25,
        64'h0ff6f813_04100693,
        64'hc2190610_06934885,
        64'h40a0053b_e6810005,
        64'h56634881_bfe900d7,
        64'h00230785_0007c683,
        64'h00d3b823_00170693,
        64'h8082852e_00070023,
        64'h00b6e663_0103b703,
        64'h40a786bb_87aa9d9d,
        64'hfff7059b_00c6f563,
        64'h8e9dfff7_06930003,
        64'hb7038f99_92010205,
        64'h96130103_b7830083,
        64'hb7038082_45018082,
        64'h00078023_45050103,
        64'hb78300a7_002300f3,
        64'hb8230017_079300d7,
        64'hfe639381_17822785,
        64'h40f707b3_0003b683,
        64'h0083b783_0103b703,
        64'h80826145_45016a02,
        64'h69a26942_64e27402,
        64'h70a22e80_00efe165,
        64'h05130000_6517fd24,
        64'h9fe30405_2fa000ef,
        64'h819100f5_f6132485,
        64'h854e0004_458330c0,
        64'h00ef8552_85a6e789,
        64'h01f4f793_20000913,
        64'h8f898993_00006997,
        64'h8f8a0a13_00006a17,
        64'h4481ed5f_f0ef8426,
        64'h45818526_33a000ef,
        64'h8f850513_00006517,
        64'hbd060613_00006617,
        64'he7898726_06130000,
        64'h6617584c_19c42783,
        64'hdb5fb0ef_e8c58593,
        64'h00006597_744805e0,
        64'h30ef91a5_05130000,
        64'h65173780_00ef90e5,
        64'h05130000_65178965,
        64'h85930000_6597c789,
        64'h8a858593_00006597,
        64'h545c3980_00ef91e5,
        64'h05130000_65175c0c,
        64'h3a6000ef_26010ff6,
        64'hf6930ff7_f7930ff7,
        64'h77130187_d61b0107,
        64'hd69b0087_d71b92e5,
        64'h05130000_651706c4,
        64'h4583583c_3d2000ef,
        64'h91c115c2_0085d59b,
        64'h93850513_00006517,
        64'h546c3e80_00ef92e5,
        64'h05130000_651706f4,
        64'h45833f80_00ef638c,
        64'h93050513_00006517,
        64'h681c2060_10ef842a,
        64'h491010ef_450144b0,
        64'h10ef0001_b50310e0,
        64'h30ef94a5_05130000,
        64'h651784aa_006030ef,
        64'he052e44e_e84aec26,
        64'hf022f406_20000513,
        64'h71797940_006f6105,
        64'h468560e2_66226442,
        64'h85a24d30_10efe42e,
        64'hec064501_842ae822,
        64'h11018082_01416402,
        64'h60a2557d_e3914505,
        64'h703c0cc0_30ef8e65,
        64'h05130000_65178d65,
        64'h85930000_659734c0,
        64'h06137626_86930000,
        64'h469702f4_02632000,
        64'h07b7e406_6380e022,
        64'h1141711c_80822501,
        64'h6108953e_050e2000,
        64'h07b7f73f_f06f2000,
        64'h05374581_46098082,
        64'hbff9557d_0e8030ef,
        64'h8522b7e5_c45c4785,
        64'hd4fd4501_88858082,
        64'h614569a2_694264e2,
        64'h740270a2_4501c45c,
        64'h4789cb99_0024f793,
        64'hf4040124_2423e01c,
        64'h200007b7_02098b63,
        64'h4fe000ef_9f450513,
        64'h00006517_862285aa,
        64'h89aa7850_10ef7c65,
        64'h05130000_451785a2,
        64'hcc1d5551_842a1000,
        64'h30ef892e_84b2e44e,
        64'hf406e84a_ec26f022,
        64'h04800513_717908b0,
        64'h41635535_b7dd87ca,
        64'h0ca139a0_20efe43e,
        64'h002c4621_8566639c,
        64'h00878913_fa978de3,
        64'h94be0009_3c830109,
        64'h648397a6_67a1bf41,
        64'hb1dff0ef_8522b771,
        64'h00f92623_000cb783,
        64'hdbd98b85_bd9560f0,
        64'h20ef4505_d80c8ee3,
        64'hc47ff0ef_8522484c,
        64'hc85c9bf5_4c85485c,
        64'hb4dff0ef_8522ef8d,
        64'h8b850089_27830009,
        64'h09630404_30232100,
        64'h30ef8556_85d20ca0,
        64'h061385a6_86930000,
        64'h56970174_8c630404,
        64'h39036004_cc9d4c85,
        64'h8889c85c_9bf9485c,
        64'hc85c0027_e793485c,
        64'hcbb5603c_feb690e3,
        64'h0791872a_2685c398,
        64'h8f518361_ff873703,
        64'h01068763_c3900086,
        64'h161bff87_05136310,
        64'h4591480d_468100c9,
        64'h0793018c_871308e6,
        64'h9f630037_f693470d,
        64'h02043c23_00492783,
        64'hcba97c1c_28e030ef,
        64'h855685d2_09c00613,
        64'h8c068693_00005697,
        64'h017c8c63_03843903,
        64'h00043c83_cfb50014,
        64'hf7936580_00efb265,
        64'h05130000_651785ca,
        64'hd1fff0ef_85ca0049,
        64'h6913ff39_79138522,
        64'h01442903_c3950084,
        64'hf7936800_00efb265,
        64'h05130000_651785ca,
        64'hd47ff0ef_85ca0089,
        64'h6913ff39_79138522,
        64'h01442903_c3950044,
        64'hf793b27f_f0ef8522,
        64'h4581b6ff_f0ef8522,
        64'h4581cc5c_f9200793,
        64'hc7817c1c_00f76f63,
        64'h0c893783_02093703,
        64'h12048e63_24818cfd,
        64'h4c81485c_07093483,
        64'h33a030ef_855685d2,
        64'h0f200613_86e20179,
        64'h09630004_3903b711,
        64'h6f6000ef_b8450513,
        64'h00006517_95458593,
        64'h00005597_000b1d63,
        64'h3b7d2000_0bb78b4e,
        64'hbd6100c4_e493bd85,
        64'h37a030ef_b9450513,
        64'h00006517_b8458593,
        64'h00006597_14900613,
        64'h97068693_00005697,
        64'hb7654701_47812585,
        64'he31c9746_93818375,
        64'h17821702_00be873b,
        64'h8fd98fe9_01076733,
        64'h0087d79b_01c87833,
        64'h0087981b_01076733,
        64'h0187971b_0187d81b,
        64'hf2e50067_036316fd,
        64'h06052781_0107e7b3,
        64'h01e8183b_07050037,
        64'h1f1b0006_4803ec06,
        64'h89e36e89_f0050513,
        64'h00ff0e37_43114701,
        64'h47814581_63900107,
        64'he6836541_00043883,
        64'h603cee07_9be38b85,
        64'h449cdf3f_f0ef8522,
        64'h488cdb7f_f0efe024,
        64'h852244cc_80826165,
        64'h45016ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h694664e6_740670a6,
        64'hefe9485c_c64a8a93,
        64'h00006a97_68198993,
        64'heb7ff0ef_25810015,
        64'he5930098_99b78522,
        64'h0d89b583_cd1ff0ef,
        64'h85224585_e93ff0ef,
        64'h85222405_8593000f,
        64'h45b7d27f_f0ef8522,
        64'h45814605_46854705,
        64'hcf5ff0ef_85224581,
        64'hcbdff0ef_852285a6,
        64'hc81ff0ef_ca4a0a13,
        64'h00006a17_85220009,
        64'h5583c4ff_f0efacec,
        64'h0c130000_5c178522,
        64'h00892583_be1ff0ef,
        64'h85224581_d71ff0ef,
        64'h85224581_46054681,
        64'h47050144_e4931607,
        64'h86638b85_008a2783,
        64'h000a0963_8cdd0324,
        64'h3c234c1c_4485e391,
        64'h448d8b89_c7090017,
        64'hf7134481_00492783,
        64'h16f99a63_04043a03,
        64'h200007b7_00043983,
        64'hbf5ff0ef_45856008,
        64'h0e049c63_6ca020ef,
        64'h00c90513_45814611,
        64'hd01ce030_84b2892e,
        64'h0005d783_020408a3,
        64'hec66f062_f45ef85a,
        64'hfc56e0d2_e4cef486,
        64'he8caeca6_7100f0a2,
        64'h71598082_61056902,
        64'h64a26442_60e2c844,
        64'h04993c23_56e030ef,
        64'hd8850513_00006517,
        64'hd7858593_00006597,
        64'h07600613_b5468693,
        64'h00005697_02f90263,
        64'h84ae842a_200007b7,
        64'hec06e426_e8220005,
        64'h3903e04a_11018082,
        64'h610564a2_644260e2,
        64'he4245b40_30efdce5,
        64'h05130000_6517dbe5,
        64'h85930000_659706f0,
        64'h0613b8a6_86930000,
        64'h569702f4_026384ae,
        64'h200007b7_ec06e426,
        64'h6100e822_11018082,
        64'h610564a2_644260e2,
        64'he0a08c7d_17fd6785,
        64'h5fa030ef_e1450513,
        64'h00006517_e0458593,
        64'h00006597_06800613,
        64'hbc068693_00005697,
        64'h02f48263_842e2000,
        64'h07b7ec06_e8226104,
        64'he4261101_80826105,
        64'h64a26442_60e2fc80,
        64'h90411442_63e030ef,
        64'he5850513_00006517,
        64'he4858593_00006597,
        64'h06100613_bf468693,
        64'h00005697_02f48263,
        64'h842e2000_07b7ec06,
        64'he8226104_e4261101,
        64'hd4dff06f_01414581,
        64'h60a26402_6008f23f,
        64'hf0ef4605_46854705,
        64'h45818522_ef1ff0ef,
        64'h45818522_f39ff0ef,
        64'h842a4581_04053023,
        64'h02053c23_46054681,
        64'h4705e022_e4061141,
        64'h80820141_45016402,
        64'h60a2d97f_f0ef4581,
        64'h6008f67f_f0ef4581,
        64'h46054685_47058522,
        64'hf35ff0ef_45818522,
        64'hf7dff0ef_e4064581,
        64'h85224605_46814705,
        64'h7100e022_11418082,
        64'h612169e2_790274a2,
        64'h02b9b823_8dc57442,
        64'h70e288a1_0125e5b3,
        64'h0034949b_8dd90049,
        64'h79130029_191b8b05,
        64'h89890014_159b6722,
        64'h722030ef_e43af3e5,
        64'h05130000_6517f2e5,
        64'h85930000_659705a0,
        64'h0613cca6_86930000,
        64'h569702f9_84638436,
        64'h893284ae_200007b7,
        64'hfc06f04a_f426f822,
        64'h00053983_ec4e7139,
        64'h80826105_64a26442,
        64'h60e2f404_76e030ef,
        64'hf8850513_00006517,
        64'hf7858593_00006597,
        64'h05300613_d0468693,
        64'h00005697_02f40263,
        64'h84ae2000_07b7ec06,
        64'he4266100_e8221101,
        64'h80826105_64a26442,
        64'h60e2f004_7ae030ef,
        64'hfc850513_00006517,
        64'hfb858593_00006597,
        64'h04c00613_d3468693,
        64'h00005697_02f40263,
        64'h84ae2000_07b7ec06,
        64'he4266100_e8221101,
        64'h80826105_64a26442,
        64'h60e2ec80_90011402,
        64'h7f2030ef_00c50513,
        64'h00006517_ffc58593,
        64'h00006597_04500613,
        64'hc4868693_00007697,
        64'h02f48263_842e2000,
        64'h07b7ec06_e8226104,
        64'he4261101_80826105,
        64'h64a26442_60e2e880,
        64'h90011402_037030ef,
        64'h05050513_00006517,
        64'h04058593_00006597,
        64'h03e00613_c9468693,
        64'h00007697_02f48263,
        64'h842e2000_07b7ec06,
        64'he8226104_e4261101,
        64'h80826105_64a26442,
        64'h60e2e404_077030ef,
        64'h09050513_00006517,
        64'h08058593_00006597,
        64'h03600613_dec68693,
        64'h00005697_02f40263,
        64'h84ae2000_07b7ec06,
        64'he4266100_e8221101,
        64'h80826105_64a26442,
        64'h60e2e004_0b7030ef,
        64'h0d050513_00006517,
        64'h0c058593_00006597,
        64'h02f00613_e1c68693,
        64'h00005697_02f40263,
        64'h84ae2000_07b7ec06,
        64'he4266100_e8221101,
        64'h80826105_64a26442,
        64'h60e2fc24_0f7030ef,
        64'h11050513_00006517,
        64'h10058593_00006597,
        64'h08800613_e4468693,
        64'h00005697_02f50263,
        64'h84ae842a_200007b7,
        64'hec06e426_e8221101,
        64'h8082556d_bfe50007,
        64'hac238082_4501cf98,
        64'h02000713_00d71763,
        64'h469100d7_0d63711c,
        64'h46a15958_80826149,
        64'h640a60aa_f83ff0ef,
        64'h0808f01f_f0ef0808,
        64'he85ff0ef_080885a2,
        64'h6622f71f_f0efe42e,
        64'he5060808_842ae122,
        64'h71758082_6105f165,
        64'h05130000_751760e2,
        64'hfca71de3_fef68fa3,
        64'hfec68f23_0007c783,
        64'h97ae0006_46038bbd,
        64'h962e0047_d6130705,
        64'h06890007_c78300e1,
        64'h07b34541_19c58593,
        64'h00006597_f5468693,
        64'h00007697_47013bf0,
        64'h20efec06_850a4641,
        64'h05050593_11018082,
        64'he13cb6c7_87930000,
        64'h0797ed3c_639cd467,
        64'h87930000_7797e93c,
        64'h04053423_639cd4e7,
        64'h87930000_77978082,
        64'h614569a2_694264e2,
        64'h740270a2_fd24fde3,
        64'h45019782_8522603c,
        64'hfc1c078e_643c0124,
        64'hf5633c90_20ef9522,
        64'h45819201_16020006,
        64'h091b40a9_863b449d,
        64'h04000993_00e78023,
        64'h97a2f800_07130017,
        64'h8513e84a_f406e44e,
        64'hec26842a_03f7f793,
        64'hf0227179_653c8082,
        64'h61616ba2_6b426ae2,
        64'h7a0279a2_794274e2,
        64'h640660a6_b7c99782,
        64'h44018526_60bc0174,
        64'h176399d6_41590933,
        64'h481020ef_0144043b,
        64'h86560084_853385ce,
        64'h020ada93_020a1a93,
        64'h00090a1b_00f97463,
        64'h93811782_00078a1b,
        64'h408b07bb_04000b93,
        64'h04000b13_e53c8932,
        64'h89ae84aa_97b203f7,
        64'hf413ec56_f052e486,
        64'he45ee85a_f44ef84a,
        64'hfc26e0a2_715d653c,
        64'h80826105_692264c2,
        64'hcd70cd34_c97c0505,
        64'h282300c8_863b00d3,
        64'h06bb00fe_07bb010e,
        64'h883b6462_f3ef9de3,
        64'h00e587bb_0005869b,
        64'h0003861b_0f118f5d,
        64'h0157171b_00b7579b,
        64'h9f3d0077_47339fa1,
        64'h8f4dfff7_47130007,
        64'h081b00b3_85bb4080,
        64'h9fa18dd5_0115d59b,
        64'h94aa00f5_969b048a,
        64'h9db5ffc2_a4038db9,
        64'h02c10075_e5b3fff7,
        64'hc593023f_44839ead,
        64'h00c703bb_00c3e633,
        64'h400c9ead_0166561b,
        64'h00a6139b_0082a583,
        64'h9e2d8e3d_8e59fff6,
        64'hc6139db1_00f8073b,
        64'h01076833_01a8581b,
        64'h0003a583_9e2d0068,
        64'h171b0107_083b0042,
        64'ha5839f2d_942a040a,
        64'h418c95aa_058a93aa,
        64'h038a020f_45839f2d,
        64'h022f4403_021f4383,
        64'h0002a703_00d745b3,
        64'h8f5dfff6_47130962,
        64'h82930000_5297f5f5,
        64'h92e300e4_07bb0004,
        64'h069b0002_861b0f91,
        64'h8f5d0177_171b0097,
        64'h579b9f3d_8f219fa5,
        64'h00574733_0007081b,
        64'h00d2843b_8ec10009,
        64'h24830106_d69b9fa5,
        64'h0106941b_992a9ea1,
        64'h090a0056_c6b300e7,
        64'hc6b3ffc3_a4839c35,
        64'h00c702bb_03c100c2,
        64'he6330156_561b013f,
        64'hc90300b6_129b4080,
        64'h00c2863b_9ea194aa,
        64'h00e2c2b3_048a00f8,
        64'h073b0083_a4039e21,
        64'h01076833_01c8581b,
        64'h0048171b_012fc483,
        64'h0107083b_40809e21,
        64'h94aa048a_0043a403,
        64'h9f21011f_c4839f25,
        64'h400000c2_c4b3942a,
        64'h040a00d7_c2b30003,
        64'ha703010f_c40311e3,
        64'h83930000_53978ffa,
        64'h1a8f0f13_00005f17,
        64'hf25599e3_00e407bb,
        64'h0004069b_0003861b,
        64'h000f081b_8f5d0147,
        64'h171b00c7_579b9f3d,
        64'h00774733_01e77733,
        64'h0083c733_9fb900d3,
        64'h843b8ec1_40980126,
        64'hd69b9fb9_00e6941b,
        64'h94aa048a_ffcfa703,
        64'h9eb90fc1_01e6c6b3,
        64'hfff5c483_8efd007f,
        64'h46b30591_9f3500cf,
        64'h03bb00c3_e6334018,
        64'h9eb90176_561b0096,
        64'h139b008f_a7039e39,
        64'h8e3d8e75_01e7c633,
        64'h9f3100f8_0f3b010f,
        64'h68330003_a70301b8,
        64'h581b9e39_00581f1b,
        64'h010f083b_004fa703,
        64'h00ef0f3b_942a040a,
        64'h4318972a_070a93aa,
        64'h038a0005_c70300ef,
        64'h0f3b0025_c4030015,
        64'hc383000f_af0301e6,
        64'hc73300cf_7f3300d7,
        64'hcf332922_82930000,
        64'h52971caf_8f930000,
        64'h5f972925_85930000,
        64'h5597f45f_17e300e3,
        64'h87bb0003_869b0005,
        64'h881b0f41_8f5d0167,
        64'h171b00a7_579b9f3d,
        64'h8f2d9fa1_00777733,
        64'h8f2d0007_061b00d7,
        64'h03bbffcf_a4039fa1,
        64'h00d3e6b3_0116969b,
        64'h00f6d39b_007686bb,
        64'h8ebd00cf_24038ef9,
        64'h00b7c6b3_00d383bb,
        64'h00c5873b_008383bb,
        64'h8e590146_561b00c6,
        64'h171b9e39_008f2383,
        64'h8e358e6d_00f6c633,
        64'h9f3100f8_05bb0077,
        64'h073b0105_e8330198,
        64'h581b0078_159b0105,
        64'h883b004f_2703ff4f,
        64'ha3839db9_007585bb,
        64'h0fc1008f_a403000f,
        64'h2583000f_a38300b6,
        64'h47338dfd_00c6c5b3,
        64'h250f8f93_00005f97,
        64'h887687f2_869a8646,
        64'h04050293_8f2ae44a,
        64'he826ec22_110105c5,
        64'h28830585_23030545,
        64'h2e030505_2e83bf89,
        64'heaf71de3_0e500793,
        64'h01814703_f8d771e3,
        64'h0007869b_02000613,
        64'h47299381_1782f4c7,
        64'he5e30585_068500e5,
        64'h8023f917_80e3b751,
        64'h842abf19_00e785a3,
        64'h47216786_ae5fd0ef,
        64'h082c462d_6506b07f,
        64'hd0ef4581_02000613,
        64'h6506f445_0005041b,
        64'ha55fe0ef_1028dbd5,
        64'h01814783_02f51b63,
        64'h4791b7c1_0005041b,
        64'h8fefe0ef_00f50223,
        64'h47857522_00f50023,
        64'h5795a885_078500c6,
        64'h802300fe_06b3b7cd,
        64'hffe81be3_06080563,
        64'h00054803_0505bfcd,
        64'hf36d8082_61256446,
        64'h60e68522_441900ee,
        64'hf863a821_00070f1b,
        64'h70850513_00006517,
        64'h93411742_370100a3,
        64'h6c639141_1542f9f7,
        64'h051b2785_0006c703,
        64'h48b107f0_0e934365,
        64'h8e2e4781_082cfeb7,
        64'h06e30007_47039736,
        64'h93010207_9713fff6,
        64'h079bbf45_863eb74d,
        64'h2605a061_00e78ca3,
        64'h00078ba3_00078b23,
        64'h04600713_00e78c23,
        64'h02100713_6786bc7f,
        64'hd0ef082c_462dc3dd,
        64'h65060181_4783e179,
        64'h2501abbf_e0ef1028,
        64'h4585e841_0005041b,
        64'hbd6fe0ef_da021028,
        64'h4581ea29_02000593,
        64'heba10007_c78397b6,
        64'h93810206_17934601,
        64'h00010c23_66a2ec55,
        64'h0005041b_ee3fd0ef,
        64'hec86e8a2_1028002c,
        64'h4605e42a_711db7d5,
        64'h842abf55_00048023,
        64'h00f51563_47918082,
        64'h61256906_64a66446,
        64'h60e68522_00a92023,
        64'hc29fd0ef_953e0347,
        64'h87930270_079300e6,
        64'h84630005_46830430,
        64'h0793470d_6562e015,
        64'h0005041b_e69fd0ef,
        64'h510c6562_02090a63,
        64'hfec783e3_177d0007,
        64'hc78397a6_93811782,
        64'h0007869b_fff6879b,
        64'hce890007_00230200,
        64'h061346ad_00b48713,
        64'hca1fd0ef_8526462d,
        64'h75c2e93d_2501b8ff,
        64'he0ef0828_4585e559,
        64'h2501ca8f_e0efd202,
        64'h08284581_c4b9e051,
        64'h0005041b_f9bfd0ef,
        64'hec86e8a2_08284601,
        64'h002c8932_84aee42a,
        64'he0cae4a6_711d8082,
        64'h61256446_60e62501,
        64'had6fe0ef_00f50223,
        64'h478500e7_8ca30087,
        64'h571b00e7_8c230044,
        64'h570300e7_8ba30087,
        64'h571b00e7_8b237522,
        64'h00645703_cb856786,
        64'heb950207_f79300b7,
        64'hc7834519_67a6e129,
        64'h25019abf_e0efe4be,
        64'h1028083c_65a2e929,
        64'h2501810f_e0efec86,
        64'h1028002c_4605842e,
        64'he42ae8a2_711dbfcd,
        64'h47a18082_614d853e,
        64'h64ea740a_70aa0005,
        64'h079bb50f_e0ef6506,
        64'he7910005_079be24f,
        64'he0ef0088_00f70223,
        64'h06d707a3_478506f7,
        64'h04a30086_d69b0106,
        64'hd69b0087_d79b0107,
        64'hd79b0107_979b06f7,
        64'h04232781_0107d79b,
        64'h06f70723_0107969b,
        64'h57d602f6_9d630557,
        64'h468302e0_07936706,
        64'hefb10005_079bfc3f,
        64'hd0ef8522_c5a54789,
        64'h0005059b_caefe0ef,
        64'h85220005_059bf2df,
        64'hd0ef85a6_00044503,
        64'h06f70863_57d64736,
        64'hcbbd8bc1_00b4c783,
        64'h00f40223_478500f4,
        64'h85a30207_e7936406,
        64'h02814783_e0dfd0ef,
        64'h00d48513_02a10593,
        64'h464d648a_efc50005,
        64'h079bdc5f_e0ef10a8,
        64'h0ce79363_4711cbf9,
        64'h0005079b_aadfe0ef,
        64'h10a86582_0c054d63,
        64'h47adf05f_d0ef850a,
        64'he49fd0ef_10a8008c,
        64'h02800613_e55fd0ef,
        64'h102805ad_46550e05,
        64'h8e634791_65e61007,
        64'h12630207_77134799,
        64'h00b7c703_77861007,
        64'h9a630005_079baf7f,
        64'he0eff0be_083cf4be,
        64'h008865a2_67861207,
        64'h96630005_079b964f,
        64'he0efed26_f122f506,
        64'h0088002c_4605e02e,
        64'he42a7171_80826165,
        64'h64e67406_70a62501,
        64'hc9efe0ef_00f50223,
        64'h47850087_05a38c3d,
        64'h02747413_8c658cbd,
        64'h752200b7_4783c30d,
        64'h6706e39d_0207f793,
        64'h00b7c783_451967a6,
        64'he9152501_b65fe0ef,
        64'he4be1028_083c65a2,
        64'he1312501_9cafe0ef,
        64'hf4861028_4605002c,
        64'h843284ae_e42aeca6,
        64'hf0a27159_b7c54421,
        64'h8082614d_6d466ce6,
        64'h7c067ba6_7b467ae6,
        64'h6a0a69aa_694a64ea,
        64'h740a70aa_8522f25f,
        64'he0ef85ca_7522441d,
        64'hb7498c6a_0ffbfb93,
        64'hf61fd0ef_3bfd8552,
        64'h45812000_0613ec09,
        64'h0005041b_8dcfe0ef,
        64'h01950223_03852823,
        64'h001c0d1b_7522a82d,
        64'h0005041b_d5afe0ef,
        64'h00f50223_47850097,
        64'h8aa30167_8a230137,
        64'h8da30157_8d2300e7,
        64'h8ca30007_8ba30007,
        64'h8b230460_071300e7,
        64'h8c230210_071300e7,
        64'h85a37522_47416786,
        64'he8350005_041bf59f,
        64'he0ef1028_040b9963,
        64'h4c850027_4b8306f4,
        64'h04a306d4_07a30087,
        64'hd79b0086_d69b0107,
        64'hd79b0106_d69b0107,
        64'h979b06f4_04232781,
        64'h0107d79b_0107969b,
        64'h06f40723_478100f6,
        64'h93635714_00d61663,
        64'h57d20007_4603468d,
        64'h05740aa3_772280ef,
        64'he0ef0544_051385d2,
        64'h049404a3_05640423,
        64'h053407a3_05540723,
        64'h040405a3_04040523,
        64'h03740a23_02000613,
        64'h04f406a3_0084d49b,
        64'h0089d99b_04600793,
        64'h0ff97a93_04f40623,
        64'h02e00b93_0104d49b,
        64'h02100793_0109d99b,
        64'h02f40fa3_0104949b,
        64'h0109199b_0ff4fb13,
        64'h47c12481_88cfe0ef,
        64'h85520200_0593462d,
        64'h898fe0ef_85520005,
        64'h0c1b4581_20000613,
        64'h03440a13_f6efe0ef,
        64'h85220109_549b85ca,
        64'h74221604_14630005,
        64'h041ba98f_e0ef7522,
        64'h16f90b63_440557fd,
        64'h16f90f63_44094785,
        64'h18090263_0005091b,
        64'hb45fe0ef_45817522,
        64'h18079f63_0207f793,
        64'h00b7c783_441967a6,
        64'h1af41763_47911c04,
        64'h09630005_041bd67f,
        64'he0efe4be_1028083c,
        64'h65a21c04_14630005,
        64'h041bbd0f_e0efe8ea,
        64'hece6f0e2_f4def8da,
        64'hfcd6e152_e54ee94a,
        64'hed26f506_f1221028,
        64'h002c4605_e42a7171,
        64'hb769d575_250191cf,
        64'hf0ef85a2_7502bf61,
        64'h2501f20f_e0ef7502,
        64'he411f155_25019f5f,
        64'he0ef1008_faf518e3,
        64'h4791d94d_2501836f,
        64'hf0ef00a8_4581f161,
        64'h2501951f_e0efcaa2,
        64'h00a84589_96cfe0ef,
        64'h00a8100c_02800613,
        64'hfc878de3_01492783,
        64'hc89d88c1_cc0d0005,
        64'h041bad8f_e0ef0009,
        64'h45037902_80826149,
        64'h794674e6_640a60aa,
        64'h451dcb81_0014f793,
        64'h00b5c483_c59975e2,
        64'heb890207_f79300b7,
        64'hc7834519_6786e105,
        64'h2501e3bf_e0efe0be,
        64'h1008081c_65a2e905,
        64'h2501ca0f_e0eff8ca,
        64'hfca6e122_e5061008,
        64'h002c4605_e42a7175,
        64'hb7b100f4_0523fbf7,
        64'hf79300a4_4783f55d,
        64'h25016480_40ef0304,
        64'h05930017_c5034685,
        64'h4c50601c_dba50407,
        64'hf79300a4_4783fcf9,
        64'h6ae34d1c_6008fcf9,
        64'h00e34509_4785b769,
        64'h449db7e1_2501a1cf,
        64'hf0ef85ca_6008f979,
        64'h2501b37f_e0ef167d,
        64'h10000637_4c0cb7dd,
        64'h450502f9_146357fd,
        64'h0005091b_94dfe0ef,
        64'h4c0cbf7d_84aa00a4,
        64'h05a3c539_00042a23,
        64'h2501a58f_f0ef484c,
        64'hef016008_00f40523,
        64'hc8180207_e793fed7,
        64'h72e34814_4458cf39,
        64'h0027f713_00a44783,
        64'h80826105_64a26902,
        64'h85266442_60e20007,
        64'h849bcb91_00b44783,
        64'he4910005_049bbc4f,
        64'he0ef842a_e04aec06,
        64'he426e822_1101bfad,
        64'h8a2abfbd_4a09b749,
        64'h4a05b7c5_39f10911,
        64'h2485e111_65820155,
        64'h75332501_abcfe0ef,
        64'he02e854a_b745fc0c,
        64'h94e33cfd_39f90909,
        64'h2485e391_8fd90087,
        64'h979b0009_47030019,
        64'h4783038b_91632000,
        64'h09930344_091385ce,
        64'he9212501_d10fe0ef,
        64'h0015899b_85220009,
        64'h9e631afd_4c094481,
        64'h49814901_10000ab7,
        64'h504cb74d_009b2023,
        64'h00f402a3_0017e793,
        64'hc8040054_4783fef9,
        64'h63e32905_4c1c2485,
        64'he1110955_08630935,
        64'h08632501_a55fe0ef,
        64'h852285ca_4a8559fd,
        64'h44814909_02fb9f63,
        64'h47850004_4b838082,
        64'h61656ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h694664e6_85527406,
        64'h70a600fb_202302f7,
        64'h6263ffec_871b481c,
        64'h01842c83_6000000a,
        64'h1c630005_0a1be7cf,
        64'he0efec66_f062f45e,
        64'hfc56e4ce_e8caeca6,
        64'hf486e0d2_8522002c,
        64'h46018b2e_e42af85a,
        64'h8432f0a2_7159bfcd,
        64'h44198082_616564e6,
        64'h740670a6_8522c10f,
        64'he0ef1028_85a6c489,
        64'hcf816786_e8010005,
        64'h041b872f_f0efe4be,
        64'h1028083c_65a2e00d,
        64'h0005041b_edafe0ef,
        64'hf486f0a2_1028002c,
        64'h460184ae_e42aeca6,
        64'h7159bf65_84aad16d,
        64'hbf7d0004_2a2300f5,
        64'h16634791_2501f8bf,
        64'he0ef8522_4581c68f,
        64'he0ef8522_85ca0004,
        64'h2a2302f5_13634791,
        64'h2501b32f_f0ef8522,
        64'h45810224_30238082,
        64'h614564e2_69428526,
        64'h740270a2_0005049b,
        64'hc5ffe0ef_85224581,
        64'h00091f63_e8890005,
        64'h049bd98f_e0ef892e,
        64'h842af406_e84aec26,
        64'hf0227179_80820141,
        64'h640260a2_00043023,
        64'he1192501_dbafe0ef,
        64'h842ae406_e0221141,
        64'hb7c1fcf5_01e34791,
        64'hbfdd4525_80826121,
        64'h744270e2_f971fcf5,
        64'h0be34791_2501cbdf,
        64'he0ef00f4_14230067,
        64'hd7838522_458167e2,
        64'hc448e30f_e0ef0007,
        64'hc50367e2_a02d0004,
        64'h30234515_e7898bc1,
        64'h00b5c783_cd996c0c,
        64'he5292501_97cff0ef,
        64'hf01c101c_e01c8522,
        64'h65a267e2_e1152501,
        64'hfe6fe0ef_0828002c,
        64'h4601842a_c52de42e,
        64'hf822fc06_7139b7bd,
        64'hc45c0137_87bb4134,
        64'h84bbcc0c_445cfaf5,
        64'hfae34f9c_601cfaba,
        64'hfee3fd45_88e30005,
        64'h059bc4bf_e0efbf69,
        64'h84cee599_0005059b,
        64'hfddfe0ef_cb818b89,
        64'h600800a4_4783b765,
        64'hcc0cc84c_b5ed4905,
        64'h00f405a3_478500f5,
        64'h976357fd_bded4909,
        64'h00f405a3_478900f5,
        64'h97634785_0005059b,
        64'h814ff0ef_e595484c,
        64'hbfb19ca9_0094d49b,
        64'hcd112501_c87fe0ef,
        64'h6008d7b5_1ff4f793,
        64'hc45c9fa5_445c0499,
        64'hea634a85_5a7dd1c1,
        64'h9c9dc45c_27814c0c,
        64'h8ff94130_07bb02c6,
        64'hed630337_563b0336,
        64'hd6bbfff4_869b377d,
        64'hc7290097_999b0025,
        64'h47836008_bf59cc44,
        64'hed352501_219040ef,
        64'h85ce0017_c5038626,
        64'h4685601c_00f40523,
        64'hfbf7f793_00a44783,
        64'hed512501_26b040ef,
        64'h0017c503_85ce4685,
        64'h601cc385_0407f793,
        64'h03040993_00a44783,
        64'hfc960ee3_4c50d3e5,
        64'h1ff7f793_445c4481,
        64'hbf7d00f4_05230207,
        64'he79300a4_4783c81c,
        64'hfcf778e3_4818445c,
        64'he4bd0004_26234458,
        64'h84bae391_8b8900a4,
        64'h47830097_77634818,
        64'h80826121_6aa26a42,
        64'h69e27902_74a2854a,
        64'h744270e2_0007891b,
        64'hcf8900b4_47830009,
        64'h17630005_091bfb4f,
        64'he0ef84ae_842ae456,
        64'he852ec4e_fc06f04a,
        64'hf426f822_7139b709,
        64'hfe9465e3_fee78fa3,
        64'h24050785_00074703,
        64'h97369281_02041693,
        64'h67220789_bddd4545,
        64'hb7e900c6_8023377d,
        64'hfc964603_962a1088,
        64'h92010207_1613b7c1,
        64'h2785b731_9c3d0136,
        64'h8023fff7_c7930127,
        64'h1a6396b2_920166a2,
        64'h02069613_00e586bb,
        64'h40f405bb_fff7871b,
        64'h04e46263_0037871b,
        64'heb05fc97_47039736,
        64'h10949301_02079713,
        64'h4781f5cf_e0ef1828,
        64'h100cb759_4509f8e5,
        64'h16e367a2_4711dd61,
        64'h2501a9ef_f0ef1828,
        64'h45810145_0e632501,
        64'h8a7fe0ef_0007c503,
        64'h65c677e2_e1052501,
        64'he48ff0ef_18284581,
        64'hf9492501_f63fe0ef,
        64'h18284581_c2aa8cdf,
        64'he0ef0007_c50365c6,
        64'h77e2f555_2501e6ef,
        64'hf0ef1828_4581fd45,
        64'h2501f89f_e0ef1828,
        64'h45858082_61497a06,
        64'h79a67946_74e6640a,
        64'h60aa0007_8023078d,
        64'h00e78123_02f00713,
        64'h0e941863_00e780a3,
        64'h03a00713_00e78023,
        64'h0307071b_13474703,
        64'h00008717_e50567a2,
        64'h4501040a_12634a16,
        64'hc2be02f0_09934bdc,
        64'h597d8426_77e2ecbe,
        64'h081ce529_2501acdf,
        64'he0ef1828_002c4601,
        64'h84ae0005_0023f0d2,
        64'hf4cef8ca_e122e506,
        64'he42afca6_7175bfd9,
        64'h4415fcf4_1ee34791,
        64'hb7c5c8c8_97bfe0ef,
        64'h0004c503_74a2cb99,
        64'h8bc100b5_c7838082,
        64'h616564e6_740670a6,
        64'h8522cbd8_575277a2,
        64'he9916586_e41d0005,
        64'h041bcd2f_f0efe4be,
        64'h1028083c_65a2ec19,
        64'h0005041b_b3bfe0ef,
        64'heca6f486_f0a21028,
        64'h002c4601_e42a7159,
        64'hbfe5452d_80826105,
        64'h60e24501_1ea78623,
        64'h00008797_00054a63,
        64'h95bfe0ef_ec060028,
        64'he42a1101_80820141,
        64'h640260a2_00043023,
        64'he1192501_9cbfe0ef,
        64'h8522e901_2501efff,
        64'hf0ef842a_e406e022,
        64'h11418082_01416402,
        64'h60a24505_ebbfe06f,
        64'h014160a2_640200f5,
        64'h02234785_00f40523,
        64'hfdf7f793_600800a4,
        64'h47830007_89a30007,
        64'h892300e7_8ca300d7,
        64'h8da30460_07130086,
        64'hd69b00e7_8c230210,
        64'h07130106_d69b00e7,
        64'h8aa30087_571b0107,
        64'h571b0107_171b00e7,
        64'h8a232701_0107571b,
        64'h0107169b_00e78d23,
        64'h00078ba3_00078b23,
        64'h485800e7_8fa300d7,
        64'h8f230187_571b0107,
        64'h569b00d7_8ea300e7,
        64'h8e230086_d69b0106,
        64'hd69b0107_169b4818,
        64'h00e785a3_02076713,
        64'h00b7c703_741ce15d,
        64'h2501b77f_e0ef6008,
        64'h500c00f4_0523fbf7,
        64'hf79300a4_4783ed55,
        64'h25015e10_40ef0304,
        64'h05930017_c5034685,
        64'h4c50601c_c3950407,
        64'hf793cf69_0207f713,
        64'h00a44783_e1752501,
        64'hacffe0ef_842ae406,
        64'he0221141_bd2d499d,
        64'hb5f9c81c_bf4100f4,
        64'h05230407_e79300a4,
        64'h47839dbf_e0ef9522,
        64'h85d28626_03050513,
        64'h0007849b_0127f463,
        64'h40ab87bb_1ff57513,
        64'h0009049b_444801a4,
        64'h2e23fd09_25016230,
        64'h40ef85da_4685001d,
        64'hc50300e7_fa63445c,
        64'h481800c7_8e634c5c,
        64'hbdd100fa_a0239fa5,
        64'h000aa783_c45c9fa5,
        64'h4099093b_445c9a3e,
        64'h93810204_97930094,
        64'h949b00f4_0523fbf7,
        64'hf79300a4_4783a4ff,
        64'he0ef855a_95d22000,
        64'h06139181_15820097,
        64'h959b0297_f26341a5,
        64'h87bb4c4c_f1512501,
        64'h6bf040ef_85d286a6,
        64'h001dc503_419704bb,
        64'h00f77463_9fb5002d,
        64'hc703c4b5_8d320007,
        64'h849b00a6_863b0099,
        64'h579b000c_869bd159,
        64'h250197cf_f0ef856e,
        64'h4c0c0004_3d8300f4,
        64'h0523fbf7_f79300a4,
        64'h4783f969_250170d0,
        64'h40ef85da_0017c503,
        64'h46854c50_601cc38d,
        64'h0407f793_00a44783,
        64'hc85ce311_cc1c4858,
        64'hbf994985_00f405a3,
        64'h47850187_9763b795,
        64'h00f40523_0207e793,
        64'h00a44783_12f76a63,
        64'h4818445c_f3fd0005,
        64'h079bd86f_f0ef4c0c,
        64'hb7594989_00f405a3,
        64'h478902e7_98634705,
        64'hcb914581_485cef01,
        64'h040c9a63_0ffcfc93,
        64'h0197fcb3_37fd0025,
        64'h47830097_5c9b6008,
        64'h14079363_1ff77793,
        64'h04090463_44585c7d,
        64'h03040b13_20000b93,
        64'h04f76c63_0127873b,
        64'h445c1807_8f638b89,
        64'h00a44783_80826165,
        64'h6da26d42_6ce27c02,
        64'h7ba27b42_7ae26a06,
        64'h69a66946_64e6854e,
        64'h740670a6_0007899b,
        64'hc39d00b4_47830009,
        64'h97630005_099bcb5f,
        64'he0ef8ab6_89328a2e,
        64'h842a0006_a023e46e,
        64'he86aec66_f062f45e,
        64'hf85aeca6_f486fc56,
        64'he0d2e4ce_e8caf0a2,
        64'h7159b59d_499dbf9d,
        64'hbd1fe0ef_855295a2,
        64'h86260305_85930007,
        64'h849b0127_f46340bb,
        64'h87bb1ff5_f5930009,
        64'h049b444c_01a42e23,
        64'hf1152501_018050ef,
        64'h85da0017_c503863a,
        64'h4685601c_00f40523,
        64'hfbf7f793_672200a4,
        64'h4783f139_250106c0,
        64'h50efe43a_85da4685,
        64'h001dc503_c38d0407,
        64'hf79300a4_478304e6,
        64'h01634c50_b70500fa,
        64'ha0239fa5_000aa783,
        64'hc45c9fa5_4099093b,
        64'h445c9a3e_93810204,
        64'h97930094_949bc5ff,
        64'he0ef9552_85da2000,
        64'h06139101_15020097,
        64'h951b0097_fc6341a5,
        64'h07bb4c48_c3850407,
        64'hf79300a4_4783f94d,
        64'h25010a60_50ef85d2,
        64'h863a86a6_001dc503,
        64'h419684bb_00f6f463,
        64'h9fb1002d_c683c4b5,
        64'h8d3a0007_849b00a6,
        64'h073b0099_579b000c,
        64'h861bd579_2501b98f,
        64'hf0ef856e_4c0c0004,
        64'h3d83cc08_b7a54985,
        64'h00f405a3_47850185,
        64'h1763b7e5_2501bd6f,
        64'hf0ef4c0c_b7414989,
        64'h00f405a3_478900a7,
        64'hec634785_4848eb11,
        64'h020c9963_0ffcfc93,
        64'h0197fcb3_37fd0025,
        64'h47830097_5c9b6008,
        64'h12079063_1ff77793,
        64'h4458fa09_0ce35c7d,
        64'h03040b13_20000b93,
        64'h0006091b_00f67463,
        64'h893e40f9_07bb445c,
        64'h01042903_16078963,
        64'h8b8500a4_47838082,
        64'h61096de2_7d027ca2,
        64'h7c427be2_6b066aa6,
        64'h6a4669e6_790674a6,
        64'h854e7446_70e60007,
        64'h899bc39d_662200b4,
        64'h47830009_98630005,
        64'h099be91f_e0ef8ab6,
        64'he4328a2e_842a0006,
        64'ha023ec6e_f06af466,
        64'hf862fc5e_e0daf0ca,
        64'hf4a6fc86_e4d6e8d2,
        64'heccef8a2_7119b7d5,
        64'h491db7e5_49118082,
        64'h61496b46_6ae67a06,
        64'h79a67946_74e6854a,
        64'h640a60aa_00f49423,
        64'h0134b023_0004ae23,
        64'h0004a623_c8880069,
        64'hd783dbbf_e0ef01c4,
        64'h0513c8c8_f33fe0ef,
        64'h0009c503_000485a3,
        64'hd09c0144_8523f480,
        64'h0309a783_85a279a2,
        64'h020a6a13_c399008a,
        64'h7793e3ad_8b850009,
        64'h84630029_f993e72d,
        64'h0107f713_00b44783,
        64'hf565a085_4921f609,
        64'h81e30049_f993e3d9,
        64'h8bc500b4_4783a895,
        64'h892ac90d_250183af,
        64'hf0ef0135_262385da,
        64'h39fd7522_e9112501,
        64'he3fff0ef_030aab03,
        64'h855685ce_04098b63,
        64'h00fa8223_0005099b,
        64'h00040aa3_00040a23,
        64'h00040da3_00040d23,
        64'h4785fc9f_e0ef85a2,
        64'h000ac503_00040fa3,
        64'h00040f23_00040ea3,
        64'h00040e23_000405a3,
        64'h00e40c23_00040ba3,
        64'h00040b23_00e40823,
        64'h000407a3_00040723,
        64'h00f40ca3_00f408a3,
        64'h02100713_04600793,
        64'h7aa2cfcd_008a7793,
        64'h6406e949_008a6a13,
        64'h2501e75f_f0ef1028,
        64'h00f51663_4791c54d,
        64'hc3e101f9_fa1301c9,
        64'hf7934519_e011e119,
        64'h64062501_b6dff0ef,
        64'he4be1028_083c65a2,
        64'h14091063_0005091b,
        64'h9d6ff0ef_1028002c,
        64'h8a7984aa_89b20005,
        64'h30231405_0d634925,
        64'he42ee8da_ecd6f0d2,
        64'hf4cefca6_e122e506,
        64'hf8ca7175_bfe5452d,
        64'h80826121_70e22501,
        64'ha0eff0ef_0828080c,
        64'h460100f6_18634785,
        64'hcb114501_e39897aa,
        64'h00070023_c3196762,
        64'h00070023_c3196622,
        64'h631800a7_8733050e,
        64'h8c078793_00009797,
        64'h04054263_83eff0ef,
        64'hf42ee432_e82efc06,
        64'h1028ec2a_7139b759,
        64'h4505bf5d_0009049b,
        64'h00f402a3_0017e793,
        64'h00544783_c81c2785,
        64'h01378a63_481cf15d,
        64'h25018aff_f0ef8522,
        64'h85a64601_03390763,
        64'hfb490ce3_bf754501,
        64'h00091463_0005091b,
        64'hec8ff0ef_852285a6,
        64'h00f4fa63_4c1c59fd,
        64'h4a05fcf5_fde384ae,
        64'h842ae052_e44ee84a,
        64'hf406ec26_f0227179,
        64'h4d1c8082_61456a02,
        64'h69a26942_64e27402,
        64'h70a24509_80824509,
        64'h00b7ed63_47858082,
        64'h610564a2_85266442,
        64'h60e200e7_82234705,
        64'h601c82af_f0ef462d,
        64'h6c08700c_84cff0ef,
        64'h45810200_06136c08,
        64'he0850005_049ba42f,
        64'hf0ef6008_484ce49d,
        64'h0005049b_fa9ff0ef,
        64'h842aec06_e426e822,
        64'h11018082_610564a2,
        64'h644260e2_451d00f5,
        64'h13634791_dd792501,
        64'hbcdff0ef_85224585,
        64'hcb990097_8d630007,
        64'hc7836c1c_ed092501,
        64'ha8cff0ef_6008484c,
        64'h0e500493_e50d2501,
        64'h88fff0ef_842ae426,
        64'hec06e822_45811101,
        64'hbfe54511_b7cd0004,
        64'h2a23d945_2501c13f,
        64'hf0ef8522_45818082,
        64'h614569a2_694264e2,
        64'h740270a2_45010097,
        64'h9a630017_b79317e1,
        64'h8bfd0337_80630327,
        64'h026303f7_f79300b7,
        64'hc783c321_0007c703,
        64'h6c1ce129_2501afaf,
        64'hf0ef6008_a0b1c90d,
        64'he199484c_49bd0e50,
        64'h09134511_84aef406,
        64'h842ae44e_e84aec26,
        64'hf0227179_bdf90ff7,
        64'h77130017_e7933701,
        64'heea866e3_0ff57513,
        64'hf9f7051b_eea87ae3,
        64'h0ff57513_fbf7051b,
        64'hbd6d4519_f11710e3,
        64'h00088663_00054883,
        64'hcf050513_00008517,
        64'h00054c63_4185551b,
        64'h0187151b_02b6f263,
        64'hfd370ae3_f95704e3,
        64'hf94706e3_f4e374e3,
        64'h00074703_97229301,
        64'h17020017_061b8732,
        64'h45ad46a1_0ff7f793,
        64'h0027979b_05659a63,
        64'hbdb9c4c8_af2ff0ef,
        64'h0007c503_609cdbe5,
        64'h8bc100b5_c7836c8c,
        64'hfbf58b91_b73d4515,
        64'hfb0dbf15_4501e807,
        64'h03e30004_bc230004,
        64'ha623cb89_0207f793,
        64'h0047f713_f4e518e3,
        64'h4711c505_00b7c783,
        64'h709c4511_bf654701,
        64'hbdfd00e9_05a39432,
        64'h92011602_00876713,
        64'h00d79463_46918bb1,
        64'h01076713_00b69463,
        64'h45850037_f6930ff7,
        64'hf7930027_979b0165,
        64'h966300d9_00234695,
        64'h00d51563_0e500693,
        64'h00094503_c6ed4711,
        64'ha06d2685_00e50023,
        64'h954a9101_02069513,
        64'h0027e793_a8dd0505,
        64'ha0d14865_02000313,
        64'h478145a1_47014681,
        64'hb7ad0240_0793943a,
        64'h12f6e063_02000693,
        64'hf7578be3_bf954709,
        64'hbf1d0405_80826121,
        64'h6b026aa2_6a4269e2,
        64'h790274a2_744270e2,
        64'h0004bc23_2501a85f,
        64'hf0ef8526_4581b791,
        64'hc55c4bdc_611cbf75,
        64'hdfdff0ef_85264581,
        64'hfed608e3_fff7c683,
        64'hfff74603_07850705,
        64'h0cb78d63_00b78593,
        64'h709cef91_8ba100b7,
        64'h4783c7e5_00074783,
        64'h6c98e96d_2501cdaf,
        64'hf0ef6088_48cc1005,
        64'h10632501_adbff0ef,
        64'h85264581_00f905a3,
        64'h02000793_943a0947,
        64'h9763470d_1b378e63,
        64'h00244783_00f900a3,
        64'h02e00793_0b379063,
        64'h00144783_01390023,
        64'h0d379263_00044783,
        64'hb40ff0ef_854a0200,
        64'h0593462d_0204b903,
        64'h0d578063_0d478263,
        64'h00044783_4b2102e0,
        64'h099305c0_0a9302f0,
        64'h0a130ae7_fc6347fd,
        64'h00044703_0004a623,
        64'h04050ce7_906305c0,
        64'h071300e7_8663842e,
        64'h84aa02f0_07130005,
        64'hc783e05a_e456e852,
        64'hec4ef04a_fc06f426,
        64'hf8227139_b7e9db1c,
        64'h27855b1c_2a856018,
        64'hf1412501_d1cff0ef,
        64'h01450223_b7b9c848,
        64'ha83ff0ef_85a6c804,
        64'h6008d91c_415787bb,
        64'h591c00fa_ed630025,
        64'h47836008_4a0502aa,
        64'h2823aa5f_f0ef8552,
        64'h85a60004_3a03beef,
        64'hf0ef0345_05134581,
        64'h20000613_6008f579,
        64'h2501dd8f_f0ef6008,
        64'hfcf48de3_57fdfcf4,
        64'h8be34785_d4bd451d,
        64'h0005049b_e81ff0ef,
        64'h480cf60a_0ee306f4,
        64'he0634d1c_6008b761,
        64'h450500f4_946357fd,
        64'hbf494509_0097e463,
        64'h47850005_049bb27f,
        64'hf0effc0a_9fe30157,
        64'hfab337fd_00495a9b,
        64'h00254783_bf5d4501,
        64'hec1c97ce_03478793,
        64'h01241523_0996601c,
        64'hfcf775e3_0009071b,
        64'h00855783_e18dc85c,
        64'h61082785_480c0009,
        64'h9d63842a_8a2e00f9,
        64'h7993d7ed_495c8082,
        64'h61216aa2_6a4269e2,
        64'h790274a2_744270e2,
        64'h4511eb99_93c1e456,
        64'he852ec4e_f4260309,
        64'h17932905_f822fc06,
        64'h00a55903_f04a7139,
        64'hbfad4405_f6f50fe3,
        64'h4785dd61_2501dbbf,
        64'hf0ef8526_85ce8622,
        64'hbf4900f4_82a30017,
        64'he7930054_c783c89c,
        64'h37fdfae7_83e3577d,
        64'hc4c0489c_02099063,
        64'he9052501_de9ff0ef,
        64'h852685a2_167d1000,
        64'h0637b76d_fb2411e3,
        64'h05450863_fd5507e3,
        64'hc9012501_c05ff0ef,
        64'h852685a2_4409bf55,
        64'h4905b7d5_faf47ee3,
        64'h894e4c9c_80826121,
        64'h6aa26a42_69e27902,
        64'h74a27442_70e28522,
        64'h547d00f4_1d6357fd,
        64'h0887f863_47850005,
        64'h041bc43f_f0efa821,
        64'h4401052a_606304f4,
        64'h63632405_4c9c5afd,
        64'h4a05844a_04f97763,
        64'h4d1c0409_0a6300c5,
        64'h2903e19d_89ae84aa,
        64'he456e852_f04af822,
        64'hfc06ec4e_f4267139,
        64'hbf3d4989_b745012a,
        64'h81a300fa_81230189,
        64'h591b0109_579b00fa,
        64'h80a30087_d79b0324,
        64'h0a230107_d79b9426,
        64'h0109179b_01256933,
        64'h8d71f000_06372501,
        64'hda0ff0ef_85569aa6,
        64'h03440a93_1fc47413,
        64'h0024141b_f80996e3,
        64'h0005099b_fd8ff0ef,
        64'h9dbd0075_d59b515c,
        64'hbf790144_82230324,
        64'h0aa30089_591b0109,
        64'h591b0109_191b0324,
        64'h0a239426_1fe47413,
        64'h0014141b_fc0992e3,
        64'h0005099b_811ff0ef,
        64'h9dbd0085_d59b515c,
        64'hb7e90127_e9339bc1,
        64'h00f97913_0089591b,
        64'h0347c783_015487b3,
        64'h80826121_6aa26a42,
        64'h69e27902_74a2854e,
        64'h744270e2_00f48223,
        64'h4785032a_8a239aa6,
        64'h0ff97913_0049591b,
        64'hc40d1ffa_fa930009,
        64'h9f630005_099b86bf,
        64'hf0ef9dbd_8526009a,
        64'hd59b50dc_00f48223,
        64'h478502fa_0a239a26,
        64'h0ff7f793_8fd98ff5,
        64'h0049179b_00f7f713,
        64'h16c16685_0347c783,
        64'h014487b3_cc191ffa,
        64'h7a130ff9_7793001a,
        64'h0a9b8805_06099663,
        64'h0005099b_8b9ff0ef,
        64'h9dbd009a_559b00ba,
        64'h0a3b515c_0015da1b,
        64'h15479463_0ee78863,
        64'h470d0ae7_8f63842e,
        64'h89324709_00054783,
        64'h0af5f063_498984aa,
        64'h4d1c16ba_75634a05,
        64'he456ec4e_f04af426,
        64'hf822fc06_e8527139,
        64'h80826105_64a28526,
        64'h644260e2_00e78223,
        64'h4705601c_00e78023,
        64'h57156c1c_f3cff0ef,
        64'h45810200_06136c08,
        64'hec990005_049b933f,
        64'hf0ef6008_484ce495,
        64'h0005049b_f33ff0ef,
        64'h842aec06_e426e822,
        64'h110100a5_5583b78d,
        64'h4505bfc1_413484bb,
        64'hf6f476e3_4f9c0009,
        64'h3783f68a_fbe30144,
        64'h0c630005_041be6ff,
        64'hf0efbf75_2501e59f,
        64'hf0ef0134_f66385a2,
        64'h00093503_4a850992,
        64'h5a7d843a_0027c983,
        64'h8722b75d_45010099,
        64'h3c2300a9_2a2394be,
        64'h03478793_049688bd,
        64'h00093783_9d3d0044,
        64'hd79bd171_00892823,
        64'h5788fce4_f7e30087,
        64'hd703eb15_579800e6,
        64'h9463470d_0007c683,
        64'he02184ae_fee474e3,
        64'h4f98611c_80826121,
        64'h6aa26a42_69e27902,
        64'h74a27442_70e24509,
        64'h00f41c63_892a4785,
        64'h00b51523_e456e852,
        64'hec4ef426_fc06f04a,
        64'h4540f822_71398082,
        64'h853e4785_b76517fd,
        64'h25011000_07b7807f,
        64'hf0ef954a_03450513,
        64'h1fc57513_0024151b,
        64'hf9352501_a39ff0ef,
        64'h9dbd0075_d59b515c,
        64'hb7598fc9_0087979b,
        64'h03494503_03594783,
        64'h99221fe4_74130014,
        64'h141bfd59_2501a63f,
        64'hf0ef9dbd_0085d59b,
        64'h515cbf45_8fe9157d,
        64'h6505bf65_8391c019,
        64'h8fc50087_979b8805,
        64'h03494783_994e1ff9,
        64'hf993f579_2501a93f,
        64'hf0ef0344_c483854a,
        64'h9dbd94ca_1ff4f493,
        64'h0099d59b_0014899b,
        64'h02492783_80826145,
        64'h853e69a2_694264e2,
        64'h740270a2_57fdc911,
        64'h2501ac7f_f0ef9dbd,
        64'h0094d59b_9cad515c,
        64'h0015d49b_00f71e63,
        64'h08d70e63_468d06d7,
        64'h0c63842e_46890005,
        64'h470302e5_f963892a,
        64'he44eec26_f022f406,
        64'he84a7179_4d180eb7,
        64'hf7634785_80824501,
        64'h80829d2d_02d585bb,
        64'h55480025_458300f6,
        64'hf96337f9_ffe5869b,
        64'h4d1c8082_610564a2,
        64'h644260e2_00a03533,
        64'h250158d0_50ef4581,
        64'h46010014_45030004,
        64'h02a35990_50ef85a6,
        64'h4685d810_22f401a3,
        64'h22e40123_20d40ca3,
        64'h20d40c23_0187d79b,
        64'h0107d71b_260522e4,
        64'h00a322f4_00230720,
        64'h06930014_45030087,
        64'h571b0107_571b0107,
        64'h971b5010_20e40f23,
        64'h445c20f4_0fa30187,
        64'hd79b0107_d71b20e4,
        64'h0ea320f4_0e230087,
        64'h571b0107_571b0107,
        64'h971b20e4_0d2302e4,
        64'h0ba30410_0713481c,
        64'h20f40da3_02f40b23,
        64'h06100793_02f40aa3,
        64'h02f40a23_05200793,
        64'h22f409a3_faa00793,
        64'h22f40923_05500793,
        64'ha01ff0ef_85264581,
        64'h20000613_03440493,
        64'h0af71b63_47850054,
        64'h47030cf7_1063478d,
        64'h00044703_ed692501,
        64'hbffff0ef_842ae426,
        64'hec06e822_1101bdc5,
        64'h9cbd0017_d79b8885,
        64'h029787bb_478db701,
        64'h0014949b_00f91563,
        64'h4789d41c_9fb5e00a,
        64'h05e3b545_a25ff0ef,
        64'h05440513_b5b90005,
        64'h099ba33f_f0ef0584,
        64'h0513b351_47810004,
        64'h2a230124_002300f4,
        64'h13233cf7_16230000,
        64'h971793c1_17c22785,
        64'h3da7d783_00009797,
        64'hc448a63f_f0ef2204,
        64'h0513c808_a6dff0ef,
        64'h21c40513_00f51c63,
        64'h27278793_25016141,
        64'h77b7a83f_f0ef2184,
        64'h051302f5_17632527,
        64'h87932501_416157b7,
        64'ha99ff0ef_03440513,
        64'h04f71263_a5570713,
        64'h4107d79b_776d0107,
        64'h979b8fd9_0087979b,
        64'h000402a3_23244703,
        64'h23344783_e13d2501,
        64'hce5ff0ef_8522001a,
        64'h859b06f7_1b634705,
        64'h4107d79b_0107979b,
        64'h8fd90087_979b0644,
        64'h47030654_478308f9,
        64'h1963478d_00f402a3,
        64'hf8000793_c45cc81c,
        64'h57fdee99_e7e32481,
        64'h0094d49b_1ff4849b,
        64'h0024949b_d408b17f,
        64'hf0ef0604_0513f00a,
        64'h15e310e9_1263470d,
        64'hd05c0354_2023cc04,
        64'hd4580157_87bb2489,
        64'h00ea873b_490d00b6,
        64'h73630905_165500b9,
        64'h39336641_19556905,
        64'hdd8d84ae_0364d5bb,
        64'h40c504bb_f4c564e3,
        64'h873200d7_063b9f3d,
        64'h004a571b_27810339,
        64'h06bbdfb1_8fd90087,
        64'h979b2501_04244703,
        64'h04344783_14050e63,
        64'h8d450085_151b0474,
        64'h44830484_4503f3c1,
        64'h00fa7793_01441423,
        64'h00fa6a33_008a1a1b,
        64'h04544783_04644a03,
        64'hffc900fb_77b3fffb,
        64'h079bfa0b_03e30164,
        64'h01230414_4b03faf7,
        64'h69e30ff7_f7930124,
        64'h01a3fff9_079b4705,
        64'h01342e23_04444903,
        64'h29811a09_866300f9,
        64'he9b30089_999b04a4,
        64'h478304b4_4983fef7,
        64'h11e32000_07134107,
        64'hd79b0107_979b8fd9,
        64'h0087979b_03f44703,
        64'h04044783_bfb947b5,
        64'hc1194a81_f6e504e3,
        64'h4785470d_b7bd00e5,
        64'h19634785_470dfe99,
        64'h15e30491_c10de9df,
        64'hf0ef8522_85d6000a,
        64'h87634509_0004aa83,
        64'h01048913_ff2a14e3,
        64'h09910941_00a9a023,
        64'h2501c5bf_f0ef854a,
        64'hc7894501_ffc94783,
        64'h89a623a4_0a131fa4,
        64'h0913848a_04f51a63,
        64'h4785ee1f_f0ef8522,
        64'h4581f569_89110009,
        64'h0463fb71_478d0015,
        64'h77130500_60ef00a4,
        64'h00a30004_00230ff4,
        64'hf5138082_6161853e,
        64'h6b426ae2_7a0279a2,
        64'h794274e2_640660a6,
        64'h47a9c111_89110009,
        64'h0563e38d_00157793,
        64'h13e060ef_00144503,
        64'hcb850004_47830089,
        64'hb023c015_47b184aa,
        64'h638097ba_65478793,
        64'h00009797_00351713,
        64'h02054e63_47addd9f,
        64'hf0ef8932_852e89aa,
        64'h00053023_e85aec56,
        64'hf052fc26_e0a2e486,
        64'hf44ef84a_715dbfcd,
        64'h450d8082_61056902,
        64'h64a26442_60e200a0,
        64'h35338d05_01257533,
        64'h2501d33f_f0ef0864,
        64'h05130097_8c634501,
        64'h0127f7b3_14650493,
        64'h00544537_fff50913,
        64'h01000537_0005079b,
        64'hd59ff0ef_06a40513,
        64'h02f71f63_a5570713,
        64'h4107d79b_776d0107,
        64'h979b8fd9_0087979b,
        64'h45092324_47032334,
        64'h4783e52d_2501fa3f,
        64'hf0ef842a_d91c0005,
        64'h022357fd_e04ae426,
        64'hec06e822_11018082,
        64'h61056902_64a26442,
        64'h60e28522_0324a823,
        64'h597d4405_c1192501,
        64'h1f4060ef_03448593,
        64'h864a4685_0014c503,
        64'hec190005_041bfddf,
        64'hf0ef892e_84aa02b7,
        64'h87634401_e04ae426,
        64'hec06e822_1101591c,
        64'h80824501_f8dff06f,
        64'hc3990045_4783b7f9,
        64'h4505b7e5_397d26c0,
        64'h60ef85ce_86269cbd,
        64'h46850014_45034c5c,
        64'hff2a74e3_4a050034,
        64'h49038082_61456a02,
        64'h69a26942_64e27402,
        64'h70a24501_00e7eb63,
        64'h40f487bb_00040223,
        64'h4c58505c_e1312501,
        64'h2ae060ef_85ce8626,
        64'h46850015_4503842a,
        64'h03450993_e052e84a,
        64'hf4065904_e44eec26,
        64'hf0227179_8082853e,
        64'h27818fd9_0107979b,
        64'h8fd50087_979b0145,
        64'hc6830155_c78300d5,
        64'h1d630007_079b8f5d,
        64'h0087979b_468d01a5,
        64'hc70301b5_c7838082,
        64'h45258082_014160a2,
        64'h4525c391_45010015,
        64'h77933200_60ef0017,
        64'hc503e406_114102e6,
        64'h90630085_57030067,
        64'hd683c70d_0007c703,
        64'hcb85611c_c915bfd5,
        64'h85074703_0000a717,
        64'h8082853a_e11c0006,
        64'h871b0789_00b66663,
        64'h0ff6f593_fd06869b,
        64'h577d4605_0007c683,
        64'hb7dd0705_a00d577d,
        64'h00d70663_00178693,
        64'h00c69863_02d5fc63,
        64'h00074683_03a00613,
        64'h02000593_cf99873e,
        64'h611c8082_61056902,
        64'h64a26442_60e20004,
        64'h002300f4_93238fd9,
        64'h0087979b_01694703,
        64'h01794783_00f49223,
        64'h8fd90087_979b0189,
        64'h47030199_4783c088,
        64'hf59ff0ef_00f58423,
        64'h84ae01c9_051300b9,
        64'h4783fcc7_9ee30685,
        64'h040500e4_00230405,
        64'h00640023_01179563,
        64'h0e500713_01071463,
        64'h00a70e63_27850006,
        64'hc703462d_02e00313,
        64'h48a54815_86ca0200,
        64'h05134781_01853903,
        64'hcfa50095_8413e04a,
        64'he426ec06_e8221101,
        64'h495cbfcd_050500b5,
        64'h00238082_00f61363,
        64'h367d57fd_b7f5fee5,
        64'h0fa30585_05050005,
        64'hc7038082_00f61363,
        64'h367d57fd_80822501,
        64'h8d5d0562_8fd907c2,
        64'h00354503_00254783,
        64'h8f5d07a2_00054703,
        64'h00154783_80820141,
        64'h60a23020_00730ff0,
        64'h000f0000_100f7ac0,
        64'h30efbba5_05130000,
        64'h95173417_907307fe,
        64'h47853007_90738fd9,
        64'h88070713_67093000,
        64'h27f37d00_30efbbe5,
        64'h05130000_95177dc0,
        64'h30efba25_05130000,
        64'h95178307_b58382e7,
        64'hb823f007_07136705,
        64'h80e7b423_8f75e406,
        64'h16fd1141_ff8006b7,
        64'h8087b703_300017b7,
        64'hb7d914fd_b7e9c35f,
        64'hf0efbfc1_710a8493,
        64'h7bf050ef_4501dff1,
        64'h54fd000a_2783bfc5,
        64'hc4fff0ef_fc075de3,
        64'h03379713_83093783,
        64'h02074563_03379713,
        64'h83093783_5a0b0493,
        64'hf4bfe0ef_8522e78d,
        64'h0009a783_e4a99e07,
        64'haf230000_a797a007,
        64'ha5230000_a797a007,
        64'hab230000_a797a007,
        64'ha7230000_a797a007,
        64'h9d230000_a797a4f7,
        64'h01a30000_a7170054,
        64'h4783a4f7_07230000,
        64'ha7170044_4783a4f7,
        64'h0ca30000_a7170034,
        64'h4783a6f7_02230000,
        64'ha7170024_4783a6f7,
        64'h07a30000_a7173000,
        64'h19370014_4783a6f7,
        64'h0f230000_a7170026,
        64'h2b376a89_00044783,
        64'h0d7030ef_c6c50513,
        64'h00009517_a945c583,
        64'h0000a597_a9d64603,
        64'h0000a617_aa66c683,
        64'h0000a697_ab184803,
        64'h0000a817_ab87c783,
        64'h0000a797_abf74703,
        64'h0000a717_113030ef,
        64'h80e7b423_8f4d91c1,
        64'h15c2ac2a_0a130000,
        64'haa170080_07378087,
        64'hb5838007_b60382e7,
        64'hb4234721_cbc50513,
        64'h00009517_8087b703,
        64'h8007b703_80e7b423,
        64'h934180a7_b0231742,
        64'h91013000_17b71502,
        64'h8f558f71_0ff6f693,
        64'h82a10086_971bf006,
        64'h06130100_063746b2,
        64'hf4fff0ef_b1498993,
        64'h0000a997_44814522,
        64'h7d8050ef_006885a2,
        64'h46097e20_50efb4f7,
        64'h05a30000_a717b4e4,
        64'h04130000_a4170028,
        64'hb5a58593_0000a597,
        64'h07f00793_4611b6f7,
        64'h05230000_a717578d,
        64'hb6f709a3_0000a717,
        64'h4789b6f7_0e230000,
        64'ha71703e0_0793b8f7,
        64'h03a30000_a71747e1,
        64'hb8078823_0000a797,
        64'h1e7030ef_e85aec56,
        64'hf052f44e_f84afc26,
        64'he0a2e486_d6c50513,
        64'h00009517_715d8082,
        64'h25018d5d_8d7900ff,
        64'h07370085_151b8fd9,
        64'h8f750085_571bf006,
        64'h86938fd9_66c10185,
        64'h579b0185_171b8082,
        64'h91411542_8d5d0522,
        64'h0085579b_80826145,
        64'h64e27402_70a28522,
        64'h8aeff0ef_bfc50513,
        64'h0000a517_04500693,
        64'hbf475703_0000a717,
        64'hbf088893_0000a897,
        64'h85a68622_47b20007,
        64'ha803c0a7_87930000,
        64'ha7970cb0_50eff406,
        64'h0068c525_85930000,
        64'ha5974611_84ae8432,
        64'hec26f022_7179bfc1,
        64'h4785eb9f_f0ef8082,
        64'h610564a2_644260e2,
        64'hc3c00c20_07b72ad0,
        64'h30efe0a5_05130000,
        64'h9517e799_0206c163,
        64'h03371693_8304b703,
        64'h300014b7_47812401,
        64'hec06e426_43c0e822,
        64'h0c2007b7_1101b7e1,
        64'hff06bc23_06a12605,
        64'h00083803_00d78833,
        64'h80826101_01135f81,
        64'h34838526_60013403,
        64'h60813083_8287b823,
        64'h300017b7_0405aa1f,
        64'hf0ef8626_02e64463,
        64'h97c285b6_30000837,
        64'h8f95868a_83f502d7,
        64'h473b1782_270546a1,
        64'h00776713_9fad377d,
        64'h8005859b_658502d5,
        64'h1a638066_86936685,
        64'hc6918005_069b0001,
        64'h550300d1_00230086,
        64'hd69b0106_d69b0106,
        64'h969b00d1_00a38726,
        64'h46d496aa_068e9ebd,
        64'h8006869b_7007f793,
        64'h0084179b_ea254390,
        64'hd2878793_0000a797,
        64'hcfb52781_8ff1fff7,
        64'hc79300c5_963b1010,
        64'h05938a1d_08b86963,
        64'h35b95f20_0813ffc5,
        64'h849b2581_60113423,
        64'h5e913c23_630c8387,
        64'hb783972a_30000537,
        64'h9f2d8406_871b0387,
        64'h75936685_0034171b,
        64'h00f67413_26016081,
        64'h30239f01_01138307,
        64'hb6033000_17b7bba5,
        64'h46013e90_30eff2e5,
        64'h05130000_951785aa,
        64'hb36900f4_16236080,
        64'h079300f4_1f230024,
        64'hd78300f4_1e230004,
        64'hd78302f4_142301e4,
        64'h578302f4_132302a0,
        64'h061301c4_57832770,
        64'h50ef8522_85ca4619,
        64'h281050ef_00640513,
        64'hdf058593_0000a597,
        64'h46192930_50ef854e,
        64'he0058593_0000a597,
        64'h46192a30_50ef854a,
        64'h85ce4619_00f59a23,
        64'h01658993_02058913,
        64'h20000793_eaf719e3,
        64'he427d783_0000a797,
        64'h0285d703_ecf711e3,
        64'he5048493_0000a497,
        64'he587d783_0000a797,
        64'h0265d703_b1e1fa65,
        64'h05130000_9517b9c9,
        64'hf9850513_00009517,
        64'hb9f1f725_05130000,
        64'h9517b1dd_f5c50513,
        64'h00009517_b9c5f4e5,
        64'h05130000_9517b9ed,
        64'hf3050513_00009517,
        64'hb311f2a5_05130000,
        64'h9517b339_f1450513,
        64'h00009517_bb21f065,
        64'h05130000_9517b30d,
        64'hef050513_00009517,
        64'hb335eea5_05130000,
        64'h9517b799_355050ef,
        64'h0868eda5_85930000,
        64'ha5974611_f4f70de3,
        64'h02045703_f6f701e3,
        64'h17fd67c1_01e45703,
        64'hf6e787e3_5fe00713,
        64'hbf95ca0f_f0ef02a4,
        64'h051385ca_53b030ef,
        64'hf1050513_00009517,
        64'hcb6ff0ef_852285a6,
        64'h54f030ef_f1450513,
        64'h00009517_02e79863,
        64'h4d200713_b765d47f,
        64'he0ef02a4_0513f1e5,
        64'h85930000_a597f1a6,
        64'h06130000_a617f1e6,
        64'h86930000_a697f7e9,
        64'h439cf2a7_87930000,
        64'ha797c799_439cf3a7,
        64'h87930000_a797f2f7,
        64'h2b230000_a71747e2,
        64'h04e69463_04300713,
        64'h80826161_79a27942,
        64'h74e26406_60a65080,
        64'h60ef4501_02a40593,
        64'hff89061b_f4c78793,
        64'h0000a797_66a24762,
        64'h429050ef_e436f6f7,
        64'h2b230000_a717f765,
        64'h05130000_a517f6e5,
        64'h85930000_a5974619,
        64'h47e2f8d7_9b230000,
        64'ha79704e7_9b6301c1,
        64'h56830450_071300e1,
        64'h0e230234_470300e1,
        64'h0ea301c1_19030224,
        64'h470300e1_0e232781,
        64'h02744703_00e10ea3,
        64'h01c11783_00f10e23,
        64'h02544783_00f10ea3,
        64'h02644703_02444783,
        64'hbdb5ffa5_05130000,
        64'h9517b559_fec50513,
        64'h00009517_bd41fde5,
        64'h05130000_9517a06d,
        64'hda5fe0ef_450185a2,
        64'h02f41223_862601c1,
        64'h578300a1_0e238121,
        64'h00a10ea3_db9ff0ef,
        64'h00f41e23_0029d783,
        64'h00f41d23_0009d783,
        64'h02f41023_02240513,
        64'hfde4859b_01c45783,
        64'h00f41f23_02041223,
        64'h02040123_01a45783,
        64'h509050ef_854a0765,
        64'h85930000_a5974619,
        64'h519050ef_852285ca,
        64'h461910f7_1c630a87,
        64'hd7830000_a7970204,
        64'h570312f7_14630b69,
        64'h89930000_a9970be7,
        64'hd7830000_a79701e4,
        64'h5703b73d_1dc50513,
        64'h00009517_f0f59ce3,
        64'h08800793_26f58963,
        64'h0ff00793_26f58863,
        64'h08900793_b73df4f5,
        64'h8ae31d25_05130000,
        64'h951706c0_079326f5,
        64'h8b630670_079300b7,
        64'hef6328f5_86630840,
        64'h0793bf91_f6f58de3,
        64'h1c050513_00009517,
        64'h05e00793_28f58463,
        64'h05c00793_b7bdf8f5,
        64'h8ae31aa5_05130000,
        64'h95170320_079328f5,
        64'h876302f0_079300b7,
        64'hef632af5_82630330,
        64'h079304b7_e2632cf5,
        64'h82630620_0793b7c9,
        64'h1a850513_00009517,
        64'hfaf596e3_02900793,
        64'h2af58663_02100793,
        64'hbf6dfef5_80e318e5,
        64'h05130000_951747d9,
        64'h16f58a63_47c500b7,
        64'hed632cf5_826347f5,
        64'ha4317c90_30effef5,
        64'h91e31725_05130000,
        64'h951747a1_18f58263,
        64'h4799a41d_7e3030ef,
        64'h30850513_00009517,
        64'h02f58363_16c50513,
        64'h00009517_478910f5,
        64'h84634785_02b7e363,
        64'h1af58363_479104b7,
        64'he5631cf5_826347b1,
        64'h08b7e763_32f58963,
        64'h02e00793_01744583,
        64'h679050ef_1ac50513,
        64'h0000a517_461985ca,
        64'h00640913_68d050ef,
        64'h46110828_84b205e9,
        64'h44079a63_8005079b,
        64'h0af50e63_6dd78793,
        64'h67a13cf5_0563842e,
        64'h80678793_f44ef84a,
        64'hfc26e486_e0a26785,
        64'h715dbf55_943e00e1,
        64'h578300f1_072300d1,
        64'h478300f1_07a334f9,
        64'h090900c1_47836df0,
        64'h50ef0068_460985ca,
        64'h80826145_91416942,
        64'h64e21542_fff54513,
        64'h740270a2_95220104,
        64'h5513942a_90411442,
        64'h01045513_02904463,
        64'h440184ae_892af406,
        64'he84aec26_f0227179,
        64'h80821e25_05130000,
        64'h9517bf75_22c50513,
        64'h00009517_84078793,
        64'hfce608e3_22c50513,
        64'h00009517_83878713,
        64'hbfe921a5_05130000,
        64'h95178287_879300c7,
        64'h4963fee6_09e323e5,
        64'h05130000_95178307,
        64'h87138082_faf612e3,
        64'h22050513_00009517,
        64'h81878793_00e60a63,
        64'h22050513_00009517,
        64'h81078713_80820141,
        64'h2a850513_0000a517,
        64'h60a21240_40efe406,
        64'h2b850513_0000a517,
        64'h2c058593_00009597,
        64'h9e3d1141_7c07879b,
        64'h77fd04c7_c9632ce5,
        64'h05130000_951787f7,
        64'h87936785_c3ad24e5,
        64'h05130000_95178006,
        64'h079b04c7_496306e6,
        64'h0b632725_05130000,
        64'h95178087_871308a7,
        64'h4463862a_0ce50763,
        64'h82078713_67858082,
        64'h953e057e_450597aa,
        64'h20000537_e3089536,
        64'h00178693_00756513,
        64'h157d631c_35470713,
        64'h0000a717_80824000,
        64'h05378082_057e4505,
        64'h8082853e_4785bf99,
        64'h03840413_2a057ed0,
        64'h50ef856a_4581864e,
        64'h1f6040ef_856285ea,
        64'h9d3e864e_40f989b3,
        64'h01843d03_0337f163,
        64'h701c0284_39830660,
        64'h60ef856a_85ee864e,
        64'h21e040ef_856686ce,
        64'h85ea866e_80826165,
        64'h853e6da2_6d426ce2,
        64'h7c027ba2_7b427ae2,
        64'h6a0669a6_694664e6,
        64'h740670a6_478d24c0,
        64'h40ef2d25_05130000,
        64'h9517864a_02bafa63,
        64'h95ce00b4_8db30184,
        64'h3d03640c_04098d63,
        64'h02043983_272040ef,
        64'h855e85d2_cbc1741c,
        64'h09679b63_401ca835,
        64'h478100fa_64630384,
        64'hd783332c_8c930000,
        64'h9c97352c_0c130000,
        64'h9c17312b_8b930000,
        64'h9b974b05_4a01942a,
        64'h84aa892e_06eae663,
        64'h478d9722_020ada93,
        64'he46ee86a_ec66f062,
        64'hf45ef85a_e0d2e4ce,
        64'he8caeca6_f4860205,
        64'h9a93fc56_7100f0a2,
        64'h02f70733_71590380,
        64'h07930385_570310e6,
        64'h97634709_00454683,
        64'h10e69c63_478957f7,
        64'h0713464c_47370005,
        64'h668312b7_f4630400,
        64'h0793bfd5_8f8d2505,
        64'h8082e21c_00b7f463,
        64'h45019181_87aa1582,
        64'hbf390705_01070023,
        64'h0005d463_4185d59b,
        64'h0185959b_c5190975,
        64'h75130005_450300bc,
        64'h05330007_4583bfdd,
        64'h4701bf1d_3cfdfe97,
        64'h6ae32705_672204e0,
        64'h70efe43a_855eb75d,
        64'h00c58023_0ff67613,
        64'h00ea85b3_0006c603,
        64'hbf6500c5_90239241,
        64'h164295d6_00171593,
        64'h0006d603_006d1c63,
        64'hbfc1e190_95d60037,
        64'h15936290_011d1863,
        64'hbf856862_78820705,
        64'h96d27322_674266a2,
        64'h3ae040ef_e436e83a,
        64'hec42f046_f41a855a,
        64'h65829201_1602c190,
        64'h260195d6_00271593,
        64'h4290030d_1b63b795,
        64'h557dd135_022070ef,
        64'h99369281_168241b4,
        64'h043b66a2_3ea040ef,
        64'hfa060c23_e43645e5,
        64'h05130000_951785d6,
        64'h963e011c_0ac5ed63,
        64'h415705bb_0006861b,
        64'h02e00813_875603bd,
        64'h06bb0d9d_e66399ba,
        64'h03470733_9301020d,
        64'h971305b6_6c630007,
        64'h061b4309_48a14811,
        64'h470186ce_000c8d9b,
        64'h008cf463_00040d9b,
        64'h446040ef_4a450513,
        64'h00009517_85ca8082,
        64'h616d6daa_6d4a6cea,
        64'h7c0a7baa_7b4a7aea,
        64'h6a0e69ae_694e64ee,
        64'h740e70ae_4501e00d,
        64'h3d8c0c13_00008c17,
        64'h450b8b93_00009b97,
        64'h4e8b0b13_00009b17,
        64'h03810a93_020a5a13,
        64'h0017849b_e03e020d,
        64'h1a13001d_179b03ac,
        64'hdcbb4cc1_000c9563,
        64'h02ccdcbb_04000c93,
        64'h00e7f663_84368d32,
        64'h89ae892a_04000793,
        64'he56ef162_f55ef95a,
        64'hfd56e1d2_eda6f586,
        64'he96ae5ce_e9caf1a2,
        64'h02c7073b_8cbaed66,
        64'h71514e80_406f6105,
        64'h54050513_00009517,
        64'h64a26902_85a6864a,
        64'h60e26442_502040ef,
        64'h53850513_00009517,
        64'h85a2c801_512040ef,
        64'h89325425_05130000,
        64'h95170585_14590087,
        64'hf46300e4_5433942a,
        64'h47a500d4_14334405,
        64'h03b6869b_02f50533,
        64'h47a9c10d_44018d7d,
        64'hfff7c793_00e797b3,
        64'h57fdb7f5_59450513,
        64'h00009517_85aafb07,
        64'h9de32785_5620406f,
        64'h61055aa5_05130000,
        64'h951785aa_690264a2,
        64'h60e26442_e495e04a,
        64'he822ec06_0007c483,
        64'he42697c2_11015f68,
        64'h08130000_a8179381,
        64'h1782cd85_00e555b3,
        64'h03c6871b_02f886bb,
        64'h481958d9_4781862e,
        64'hb78d5ca5_05130000,
        64'h951785aa_5ba0406f,
        64'h61055fa5_05130000,
        64'h95176902_64a285ca,
        64'h862660e2_64425d40,
        64'h40ef60a5_05130000,
        64'h951785a2_c8015e40,
        64'h40ef84b2_61450513,
        64'h00009517_f86102f4,
        64'h5433bfc1_02e45433,
        64'ha039943e_00144413,
        64'h03243413_02e47433,
        64'h02f457b3_06400713,
        64'h02877463_06300713,
        64'hc70502f4_773347a9,
        64'h0287e663_47293e80,
        64'h0793c021_02f555b3,
        64'h02f57433_bf7d2407,
        64'h87934685_b7d9a007,
        64'h87934681_64a0406f,
        64'h610566a5_05130000,
        64'h951785aa_690264a2,
        64'h60e26442_02091663,
        64'he426e822_ec060007,
        64'h4903e04a_97361101,
        64'h6e870713_0000a717,
        64'h3e800793_46890ca7,
        64'hf7633e70_079304a7,
        64'h676323f7_8713000f,
        64'h47b704a7_6963862e,
        64'h9ff78713_3b9ad7b7,
        64'h8082612d_450160ee,
        64'h6ae040ef_6c450513,
        64'h00009517_002cfebf,
        64'hf0efed86_45050c80,
        64'h0613002c_7115f73f,
        64'hf06f4581_862e86b2,
        64'h80826145_69a26942,
        64'h64e2854a_740270a2,
        64'h27c060ef_6dc58593,
        64'h00009597_00890533,
        64'hffd4841b_00f44463,
        64'hffe4879b_9c296c40,
        64'h40ef954a_70c60613,
        64'h00009617_86ce40a4,
        64'h85bb0095_5d630009,
        64'h8f63842a_6e2040ef,
        64'h854a85a6_72460613,
        64'h00009617_bfc70713,
        64'h00009717_72c68693,
        64'h00009697_c509fce6,
        64'h86930000_a6978932,
        64'h89ae84b6_f022f406,
        64'he44ee84a_ec267179,
        64'hbfdd7600_40ef8562,
        64'hb7e90905_76a040ef,
        64'h856600fb_e7630ff7,
        64'hf793fe05_879b0007,
        64'hc583012a_07b3b781,
        64'h04852405_78a040ef,
        64'h2b850513_0000a517,
        64'h00f45b63_0009079b,
        64'hff047913_7a2040ef,
        64'h855aff2d_cce32d85,
        64'h7ae040ef_8556a029,
        64'h00f97913_4d81fffd,
        64'h4913028d_1d637c40,
        64'h40ef7b25_05130000,
        64'h95170104_c583dbe5,
        64'hb7c57d80_40ef8562,
        64'ha0317e00_40ef8556,
        64'h7e6040ef_31450513,
        64'h0000a517_ffb912e3,
        64'h09057f80_40ef8566,
        64'h02fbe263_0ff7f793,
        64'hfe05879b_0007c583,
        64'h012487b3_4dc14901,
        64'h017040ef_855ae7a9,
        64'hc42900f4_77938082,
        64'h61656da2_6d426ce2,
        64'h7c027ba2_7b427ae2,
        64'h6a0669a6_694664e6,
        64'h740670a6_03344163,
        64'hfff58d1b_824c8c93,
        64'h0000ac97_834c0c13,
        64'h0000ac17_06000b93,
        64'h828b0b13_0000ab17,
        64'h540a8a93_0000aa97,
        64'h4401ff05_049389ae,
        64'h8a2ae46e_e8caf486,
        64'he86aec66_f062f45e,
        64'hf85afc56_e0d2e4ce,
        64'heca6f0a2_7159b7cd,
        64'h097040ef_9e07ae23,
        64'h0000b797_85450513,
        64'h0000a517_80826151,
        64'h641260b2_85220b50,
        64'h40ef83a5_05130000,
        64'ha5178125_85930000,
        64'ha597860a_c10d842a,
        64'hdedff0ef_85220d50,
        64'h40ef8325_05130000,
        64'ha5178325_85930000,
        64'ha597842a_00054603,
        64'h00154683_00254703,
        64'h00354783_00454803,
        64'h00554883_e222e606,
        64'h716d8082_7f010113,
        64'h7c813983_7d013903,
        64'h7d813483_7e013403,
        64'h45017e81_30836165,
        64'h8cfff0ef_86c685a6,
        64'h18085632_6882fbaf,
        64'hf0ef03e1_0513863e,
        64'h86c285a2_67c26822,
        64'hf8aff0ef_d64e0521,
        64'h051385a2_864a86ba,
        64'h943e7fc4_04136762,
        64'h747d97ba_81078793,
        64'h10186785_7bc060ef,
        64'hd602e83e_ec3ae442,
        64'h893689b2_e04605a1,
        64'h051384aa_71597d31,
        64'h34237d21_38237c91,
        64'h3c237e81_30237e11,
        64'h34238101_011319d0,
        64'h406f8e25_05130000,
        64'ha51785aa_80826125,
        64'h7aa27a42_79e26906,
        64'h64a66446_450160e6,
        64'h911a6305_96bff0ef,
        64'h85ce86a6_10084652,
        64'h855ff0ef_460156fd,
        64'h02e10513_85a2821f,
        64'hf0ef0440_06130430,
        64'h06930421_051385a2,
        64'h943e1451_978a020a,
        64'h879312f1_1c233537,
        64'h87936799_12f11b23,
        64'h26378793_77e105f0,
        64'h60ef04f1_06230661,
        64'h05134641_479985ce,
        64'h04f11523_10100793,
        64'h027060ef_ca3e04a1,
        64'h05134581_0f000613,
        64'h0fc00793_08d060ef,
        64'h000107a3_15410223,
        64'h14f101a3_14510513,
        64'h460585ca_57fd0a70,
        64'h60ef13f1_05134611,
        64'h95beff04_0593978a,
        64'h020a8793_12f10f23,
        64'h479112f1_0ea30370,
        64'h07930cb0_60ef0141,
        64'h07a31a68_460585ca,
        64'h993e978a_020a8793,
        64'h12f11d23_13500793,
        64'hc83e4a05_fef40913,
        64'h439cb027_87930000,
        64'hb7970a90_60ef8526,
        64'h55fd4619_94beff84,
        64'h0493978a_020a8793,
        64'h747d2c10_40efca02,
        64'h6a859f25_05130000,
        64'ha517911a_89aaf456,
        64'hf852fc4e_e0cae4a6,
        64'he8a2ec86_711d737d,
        64'hb35d2e90_40ef9de5,
        64'h05130000_a517bf45,
        64'h9d850513_0000a517,
        64'h95be978a_d0040593,
        64'h35078793_678530d0,
        64'h40ef9d25_05130000,
        64'ha5173190_40ef9ce5,
        64'h05130000_a51700fa,
        64'h20234785_de0796e3,
        64'h000a2783_bbcd3350,
        64'h40ef9da5_05130000,
        64'ha517b501_343040ef,
        64'h9d050513_0000a517,
        64'h95be978a_f0040593,
        64'h35048793_35b040ef,
        64'h9d850513_0000a517,
        64'h95bee004_0593978a,
        64'h35048793_373040ef,
        64'h02f5d5bb_e107879b,
        64'h678502f6_763b02f5,
        64'hf6bb02f5_d63b03c0,
        64'h0793d4f7_1e230000,
        64'hb7170121_5783d6f7,
        64'h13230000_b7179fe5,
        64'h05130000_a51755c2,
        64'h01015783_3b3040ef,
        64'h9f050513_0000a517,
        64'h01014583_01114603,
        64'h01214683_01314703,
        64'h3cf040ef_9ec50513,
        64'h0000a517_01814583,
        64'h01914603_01a14683,
        64'h01b14703_3eb040ef,
        64'h00b14703_dcf71323,
        64'h0000b717_9ec50513,
        64'h0000a517_00814583,
        64'h35215783_dcf71e23,
        64'h0000b717_00914603,
        64'h00a14683_35015783,
        64'h41f040ef_9ec50513,
        64'h0000a517_35014583,
        64'h35114603_35214683,
        64'h35314703_28d060ef,
        64'h01490593_4611953e,
        64'hcb840513_978a3504,
        64'h87936485_2a5060ef,
        64'h0e880109_05934611,
        64'h45f040ef_a1c50513,
        64'h0000a517_00fa2023,
        64'h47851207_9a63000a,
        64'h2783b311_d00d0023,
        64'h2d1060ef_9d228562,
        64'h866ab759_cc048513,
        64'hbb29cef4_2023401c,
        64'h00f40023_ce344783,
        64'h00f400a3_ce244783,
        64'h00f40123_ce144783,
        64'h00f401a3_ce044783,
        64'h309060ef_4611953e,
        64'hce048513_978a3507,
        64'h87936785_bfdd855a,
        64'h4611bbb1_325060ef,
        64'h85564611_b39df00d,
        64'h00233330_60ef9d22,
        64'h953e866a_f0048513,
        64'h978a3507_87936785,
        64'ha00d953e_978a3507,
        64'h87936785_4611cd04,
        64'h85138082_3b010113,
        64'h35013d03_35813c83,
        64'h36013c03_36813b83,
        64'h37013b03_37813a83,
        64'h38013a03_38813983,
        64'h39013903_39813483,
        64'h3a013403_3a813083,
        64'h911a6305_cebff0ef,
        64'h0e8885de_86ca5672,
        64'hbd5ff0ef_35e10513,
        64'h85a24601_56fdba1f,
        64'hf0ef3721_051385a2,
        64'h04400613_04300693,
        64'h943ecec4_0413978a,
        64'h350a8793_46f11423,
        64'h35378793_679946f1,
        64'h13232637_879377e1,
        64'h3e1060ef_36f10e23,
        64'h39610513_85de4799,
        64'h464136f1_1d231010,
        64'h07933a90_60efde3e,
        64'h37a10513_45810f00,
        64'h06131020_079340f0,
        64'h60ef4731_0d230001,
        64'h03a346f1_0ca347b1,
        64'h051385a6_460557fd,
        64'h429060ef_47410a23,
        64'h47510513_461195be,
        64'hcf440593_978a350a,
        64'h879346f1_09a30360,
        64'h079344b0_60ef4741,
        64'h072346f1_05134611,
        64'h4a1195be_cf040593,
        64'h978a350a_879346f1,
        64'h06a30320_079346f0,
        64'h60efc0d2_46c10513,
        64'h85a64605_94becb74,
        64'h0493c2a6_978a350a,
        64'h879346f1_15231350,
        64'h079300f1_03a3478d,
        64'h447060ef_854a55fd,
        64'h4619993e_cf840913,
        64'h978a350a_879365d0,
        64'h40efde02_54e25a52,
        64'hc0850513_0000a517,
        64'h4c1060ef_953e4611,
        64'h01490593_ce840513,
        64'h978a350a_87934d70,
        64'h60ef013c_a023953e,
        64'h46110109_0593ce44,
        64'h05134985_978a350a,
        64'h87936a85_16079263,
        64'h000ca783_3ae79d63,
        64'h470938e7_81634719,
        64'h24e78163_0007859b,
        64'h747d4715_00614783,
        64'hf8e79ce3_0ff00713,
        64'h24e78563_03800713,
        64'haad94605_cb648513,
        64'hfae798e3_03500713,
        64'h22e78063_03300713,
        64'h00f76e63_22e78363,
        64'h03600713_b759e00d,
        64'h00235530_60ef9d22,
        64'h953e866a_e0048513,
        64'h978a3507_87936785,
        64'hfee794e3_473d22e7,
        64'h85634731_b77d7250,
        64'h40efe325_05130000,
        64'ha51785b6_22e78963,
        64'hcc848513_470d2ae7,
        64'h89634705_02f76263,
        64'h24e78163_471904f7,
        64'h6b6326e7_8d630007,
        64'h869b01a9_89bb0589,
        64'h02a00713_29890f07,
        64'hc7830015_cd030139,
        64'h07b395ca_0f098593,
        64'h9c3a9b3a_49818a36,
        64'h8cb28bae_d0048c13,
        64'hcb848b13_970a3507,
        64'h87139aba_cd848a93,
        64'h970a3507_871374fd,
        64'h678526f7_11634789,
        64'h00054703_a0017ad0,
        64'h40efd325_05130000,
        64'ha51785aa_00e7ea63,
        64'h892a5800_073797aa,
        64'hd0040023_f0040023,
        64'he0040023_ca040b23,
        64'hce042023_d00007b7,
        64'h943e747d_978a911a,
        64'h35078793_35a13823,
        64'h35913c23_37813023,
        64'h37713423_37613823,
        64'h37513c23_39413023,
        64'h39313423_38913c23,
        64'h3a113423_39213823,
        64'h3a813023_6785737d,
        64'hc5010113_fadff06f,
        64'h614564e2_00e4859b,
        64'h70a27402_852200f4,
        64'h162347a1_68d060ef,
        64'h85b64619_852266a2,
        64'h699060ef_e436f406,
        64'h46190519_84b2842a,
        64'hec26f022_71798082,
        64'h01416402_60a28522,
        64'hfa5ff0ef_e4064501,
        64'h85aa8622_0005841b,
        64'he0221141_bff105a1,
        64'h25050116_b02396ba,
        64'h010686bb_0035169b,
        64'h0005b883_808280c7,
        64'h3823973e_678500f5,
        64'h47636805_450102d7,
        64'hc7bb2785_0077e793,
        64'hfff6079b_8007bc23,
        64'h97ba46a1_67856398,
        64'h13878793_0000b797,
        64'h80826145_740270a2,
        64'h00f41523_fff7c793,
        64'h9fb94107_d71b9fb9,
        64'h93411742_4107579b,
        64'hfed79ce3_9f31ffe7,
        64'hd6030789_470187a2,
        64'h01440693_74d060ef,
        64'h01040513_002c4611,
        64'h759060ef_00c40513,
        64'h00041523_006c4611,
        64'h00f404a3_47c576f0,
        64'h60efec3e_00840513,
        64'h00041323_082c4621,
        64'h47c17830_60ef0044,
        64'h05130161_05934609,
        64'h791060ef_00f11b23,
        64'hc4360509_084c57fd,
        64'h460900f1_1a238fd9,
        64'h0087979b_0ff77713,
        64'h0087d713_c632842a,
        64'h419c00f5_10230457,
        64'h879b6785_c19c27d1,
        64'hf022f406_7179419c,
        64'h80820005_132300f5,
        64'h122300d5_112300c5,
        64'h10238fd9_0087979b,
        64'h0ff77713_c19c0087,
        64'hd7138ed9_06a20086,
        64'hd71b8e59_27a10622,
        64'h0086571b_419cc19c,
        64'h2785c319_0017f713,
        64'h419cbfcd_fda00513,
        64'h80826121_74a27442,
        64'h70e29782_85a66562,
        64'h701ce509_c39ff0ef,
        64'h842a0830_65a2c105,
        64'hc7dff0ef_84b2e42e,
        64'hf822fc06_f4267139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2655c,
        64'h862686ca_6562e519,
        64'hc75ff0ef_083065a2,
        64'hc115cb7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2615c,
        64'h862686ca_6562e519,
        64'hcb5ff0ef_083065a2,
        64'hc115cf7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hb7e16522_f569cdbf,
        64'hf0ef8526_85ce0030,
        64'hbfc90284_8493c501,
        64'h6a3060ef_854a608c,
        64'h296050ef_855285ca,
        64'h60908082_61216a42,
        64'h69e27902_74a27442,
        64'h70e24501_00849b63,
        64'h942602f4_043302ea,
        64'h0a130000_aa1789ae,
        64'h892afc06_e852ec4e,
        64'hf04a0280_079302f4,
        64'h043b840d_8c053a24,
        64'h84930000_b4973aa4,
        64'h04130000_b417f426,
        64'hf822639c_29c78793,
        64'h0000b797_7139bfdd,
        64'h45018082_61056442,
        64'h60e2fda0_05138302,
        64'h610560e2_65a26442,
        64'h85220003_0e630205,
        64'h3303c919_db9ff0ef,
        64'he42eec06_4108842a,
        64'he8221101_bfc56562,
        64'hf96dd97f_f0ef0830,
        64'h80826145_70a24501,
        64'he50965a2_de1ff0ef,
        64'hf406e42e_7179bfc1,
        64'h5479fcf7_1be30ff0,
        64'h079300c7_c70367a2,
        64'h04e080ef_6522f565,
        64'h842adcff_f0ef85a6,
        64'h00308522_80826145,
        64'h64e27402_70a28522,
        64'h543507a0_80ef0ee5,
        64'h05130000_a51700f4,
        64'hcf63445c_39a050ef,
        64'h0f050513_0000a517,
        64'h85a6842a_c11dfda0,
        64'h0413e47f_f0ef84ae,
        64'hf406ec26_f0227179,
        64'h80826145_694264e2,
        64'h740270a2_85220b40,
        64'h80ef6522_3d2050ef,
        64'h11850513_0000a517,
        64'h864a608c_ed01842a,
        64'he45ff0ef_84aa85ca,
        64'h0030c11d_fda00413,
        64'he8dff0ef_892eec26,
        64'hf406e84a_f0227179,
        64'hb7d92405_0f2080ef,
        64'h65224100_50ef854e,
        64'h85a20127_896300c7,
        64'hc78367a2_ed09e83f,
        64'hf0ef8526_85a20030,
        64'h80826121_69e27902,
        64'h74a27442_70e200f4,
        64'h496344dc_17498993,
        64'h0000a997_0ff00913,
        64'h440184aa_cd01eebf,
        64'hf0efec4e_f04af426,
        64'hf822fc06_7139bfd5,
        64'h54798082_61457402,
        64'h70a28522_158080ef,
        64'h00f70963_00c54703,
        64'h0ff00793_6562e911,
        64'h842aee7f_f0ef0830,
        64'h65a2c105_fda00413,
        64'hf2dff0ef_e42ef406,
        64'hf0227179_b7c1fda0,
        64'h0513bf65_24051920,
        64'h80ef4981_65224b40,
        64'h50ef8552_00099563,
        64'h2485cb99_0087c783,
        64'h67a2ed19_f29ff0ef,
        64'h854a85a2_00308082,
        64'h61216a42_69e27902,
        64'h74a27442_70e24501,
        64'hc0915535_00f44d63,
        64'h00c92783_01ca0a13,
        64'h0000ba17_44014481,
        64'h4985892a_cd31f9bf,
        64'hf0efe852_ec4ef04a,
        64'hf426f822_fc067139,
        64'hbfe54501_80820141,
        64'h60a26108_c509fbbf,
        64'hf0efe406_1141b7f5,
        64'h02870713_fea68de3,
        64'h47148082_853a4701,
        64'h00e79563_97ba02d7,
        64'h87b30280_069302d7,
        64'h87bb878d_8f9961a7,
        64'h87930000_b7976294,
        64'h62470713_0000b717,
        64'h51068693_0000b697,
        64'hb7edfda0_07138302,
        64'h853e85b2_00030563,
        64'h01853303_8082853a,
        64'he21c97b6_470102a7,
        64'h87b30a00_051300b7,
        64'hd963454c_0005cc63,
        64'h5735c285_87ae6914,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h000a2e2e_2e746e65,
        64'h6d6f6d20_61207469,
        64'h61772065_7361656c,
        64'h50202165_6e616972,
        64'h41206d6f_7266206f,
        64'h6c6c6548_ffdff06f,
        64'h10500073_34102373,
        64'h342022f3_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_4ce090ef,
        64'hfec5c6e3_02058593,
        64'h0005bc23_0005b823,
        64'h0005b423_0005b023,
        64'hd9060613_0000c617,
        64'h83058593_0000c597,
        64'h30579073_09078793,
        64'h00000797_00078067,
        64'h40b787b3_00d787b3,
        64'h01478793_00000797,
        64'hfcc5cce3_02068693,
        64'h02058593_00e6bc23,
        64'h0185b703_00e6b823,
        64'h0105b703_00e6b423,
        64'h0085b703_00e6b023,
        64'h0005b703_0006b703,
        64'hff810113_01b11113,
        64'h0110011b_fe0e9ae3,
        64'h0085b703_fffe8e93,
        64'h0005b703_240e8e9b,
        64'h000f4eb7_01169693,
        64'hfff6869b_000066b7,
        64'h81c60613_0000c617,
        64'hfc058593_00000597,
        64'h000280e7_13050513,
        64'h00000517_09428293,
        64'h00008297_000280e7,
        64'h06e28293_00008297,
        64'h01111113_fff1011b,
        64'h00006137_11249463,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
