/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module etherboot (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 6034;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h87fe705c_00000000,
        64'h87fe709a_00000000,
        64'h00000000_ffffffff,
        64'h00000006_00000000,
        64'h87feb5b0_cc33aa55,
        64'h00000000_2f7c5c2d,
        64'h00000000_87feb3f8,
        64'h00000000_ffffffff,
        64'h00006772_615f6473,
        64'h0000646d_635f6473,
        64'h00000000_0c000000,
        64'h00000000_ffffffff,
        64'h00000000_00000000,
        64'h00000000_43000000,
        64'h00000000_004b4d47,
        64'h00004b4d_47545045,
        64'h00000003_0f060301,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'haaaaaaaa_aaaaaaaa,
        64'h55555555_55555555,
        64'h5851f42d_4c957f2d,
        64'h10000000_20000000,
        64'h10325476_98badcfe,
        64'hefcdab89_67452301,
        64'h00000002_464c457f,
        64'hcccccccc_cccccccd,
        64'h00000a0d_70617274,
        64'h00000000_000a7473,
        64'h65742065_68636143,
        64'h00000000_00000a74,
        64'h6f6f6220_50544654,
        64'h00000000_00000a74,
        64'h73657420_4d415244,
        64'h00000000_00000a74,
        64'h6f6f6220_49505351,
        64'h00000000_00000000,
        64'h0a746f6f_62204453,
        64'h00000000_0000000a,
        64'h5825203d_20646565,
        64'h73206d6f_646e6152,
        64'h000a5825_2c582520,
        64'h3d20676e_69747465,
        64'h73206863_74697753,
        64'h0000000a_5825203d,
        64'h205d6425_5b707773,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h0a646c25_2e646c25,
        64'h203d2049_5043202c,
        64'h73656c63_79632064,
        64'h6c25202c_736e6f69,
        64'h74637572_74736e69,
        64'h20646c25_202c424b,
        64'h6425203d_20746573,
        64'h5f676e69_6b726f77,
        64'h00000000_00000000,
        64'h0a2e2979_6c6e6f28,
        64'h2032206e_6f697372,
        64'h65762065_736e6563,
        64'h694c2063_696c6275,
        64'h50206c61_72656e65,
        64'h4720554e_47206568,
        64'h74207265_646e7520,
        64'h6465736e_6563694c,
        64'h00000000_0000000a,
        64'h2e6e6f62_617a6143,
        64'h2073656c_72616843,
        64'h20323130_322d3130,
        64'h30322029_43282074,
        64'h68676972_79706f43,
        64'h00000000_0000000a,
        64'h29746962_2d642528,
        64'h20302e33_2e34206e,
        64'h6f697372_65762072,
        64'h65747365_746d656d,
        64'h00000a74_73657420,
        64'h4d415244_206c6174,
        64'h656d2065_7261420a,
        64'h00000a2e_656e6f44,
        64'h00000000_000a6b6f,
        64'h0000203a_73252020,
        64'h00000073_73657264,
        64'h6441206b_63757453,
        64'h00000000_00000a3a,
        64'h00000000_0075252f,
        64'h00752520_706f6f4c,
        64'h00000000_000a7025,
        64'h7830206f_74207025,
        64'h78302073_69206567,
        64'h6e617220_74736574,
        64'h00000000_00082008,
        64'h00000000_00000008,
        64'h08080808_08080808,
        64'h08082020_20202020,
        64'h20202020_20080808,
        64'h08080808_08080808,
        64'h00000000_0000000a,
        64'h2e2e2e74_73657420,
        64'h7478656e_206f7420,
        64'h676e6970_70696b53,
        64'h00000000_000a2e78,
        64'h25783020_74657366,
        64'h666f2074_6120656e,
        64'h696c2073_73657264,
        64'h64612064_61622065,
        64'h6c626973_736f7020,
        64'h3a455255_4c494146,
        64'h00000000_00007525,
        64'h20676e69_74736574,
        64'h00000000_00007525,
        64'h20676e69_74746573,
        64'h00000000_00080808,
        64'h08080808_08080808,
        64'h00000000_00202020,
        64'h20202020_20202020,
        64'h00000000_0000000a,
        64'h7025203d_20327020,
        64'h2c702520_3d203170,
        64'h00000a2e_78257830,
        64'h20746573_66666f20,
        64'h74612078_25783020,
        64'h3d212078_25783020,
        64'h3a455255_4c494146,
        64'h00000000_000a7325,
        64'h206e6f69_74636e75,
        64'h66202c64_2520656e,
        64'h696c202c_73252065,
        64'h6c696620_2c64656c,
        64'h69616620_7325206e,
        64'h6f697472_65737361,
        64'h00000a72_6564616f,
        64'h6c20746f_6f622065,
        64'h67617473_20747372,
        64'h69662064_65736162,
        64'h20746f6f_622d750a,
        64'h00000000_216b7369,
        64'h6420746e_756f6d75,
        64'h206f7420_6c696166,
        64'h00000000_0021656c,
        64'h69662065_736f6c63,
        64'h206f7420_6c696166,
        64'h0000000a_21746f6f,
        64'h62206e65_706f206f,
        64'h74206465_6c696146,
        64'h00000000_00000000,
        64'h6e69622e_746f6f62,
        64'h00000000_00000a79,
        64'h726f6d65_6d206f74,
        64'h6e69206e_69622e74,
        64'h6f6f6220_64616f4c,
        64'h00000000_0000000a,
        64'h21726576_69726420,
        64'h44532074_6e756f6d,
        64'h206f7420_6c696146,
        64'h00000000_0000000a,
        64'h2e2e2e70_25207373,
        64'h65726464_61207461,
        64'h206d6172_676f7270,
        64'h20646564_616f6c20,
        64'h65687420_746f6f42,
        64'h00000000_5c2d2f7c,
        64'h000a7825_203d206c,
        64'h61757463_61202c58,
        64'h25203d20_64657269,
        64'h75716572_206e656c,
        64'h00000000_00000000,
        64'h0a2e6e6f_69746172,
        64'h65706f20_50544654,
        64'h206c6167_656c6c49,
        64'h00000000_000a2e64,
        64'h656c6c61_63207172,
        64'h775f656c_646e6168,
        64'h00000000_00000a2e,
        64'h646e6520_656c6966,
        64'h20657669_65636552,
        64'h00000000_00000000,
        64'h0a64253d_657a6973,
        64'h6b636f6c_62202c22,
        64'h73252220_3a717277,
        64'h00000000_0000002f,
        64'h00000000_000a646c,
        64'h25202e67_6e6f6c20,
        64'h6f6f7420_68746170,
        64'h20747365_75716552,
        64'h00000064_6c252065,
        64'h646f6320_68746977,
        64'h2064656c_69616620,
        64'h64616572_20666c65,
        64'h000a7972_6f6d656d,
        64'h20524444_206f7420,
        64'h666c6520_64616f6c,
        64'h00000000_00000000,
        64'h0a732520_3d202964,
        64'h252c7025_2835646d,
        64'h00000000_0000000a,
        64'h6425203d_20687467,
        64'h6e656c20_656c6946,
        64'h00000000_00636d6d,
        64'h00000029_73252820,
        64'h00006425_203a7325,
        64'h00000000_00004453,
        64'h00000000_434d4d65,
        64'h00000000_00000000,
        64'h0a646e75_6f662074,
        64'h6f6e2064_25206563,
        64'h69766544_20434d4d,
        64'h0000297a_484d3030,
        64'h32282030_30325348,
        64'h00000000_00297a48,
        64'h4d383032_28203430,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282030,
        64'h35524444_20534855,
        64'h00000000_0000297a,
        64'h484d3030_31282030,
        64'h35524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282035,
        64'h32524453_20534855,
        64'h00000000_00000029,
        64'h7a484d35_32282032,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d32_35282032,
        64'h35524444_20434d4d,
        64'h0000297a_484d3235,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000029_7a484d30,
        64'h35282064_65657053,
        64'h20686769_48204453,
        64'h0000297a_484d3632,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000000_00000079,
        64'h63616765_4c204453,
        64'h00000000_00007963,
        64'h6167656c_20434d4d,
        64'h00000064_252e6425,
        64'h00000000_63256325,
        64'h63256325_63256325,
        64'h00000078_34302578,
        64'h34302520_726e5320,
        64'h78363025_206e614d,
        64'h00000000_00000a21,
        64'h646e756f_66206473,
        64'h635f7478_65206f4e,
        64'h00000000_00000000,
        64'h0a65646f_6d206120,
        64'h7463656c_6573206f,
        64'h7420656c_62616e75,
        64'h00000000_00000000,
        64'h0a217463_656c6573,
        64'h20656761_746c6f76,
        64'h206f7420_646e6f70,
        64'h73657220_746f6e20,
        64'h64696420_64726143,
        64'h0000000a_746e6573,
        64'h65727020_64726163,
        64'h206f6e20_3a434d4d,
        64'h00000000_0000000a,
        64'h64656e6f_69746974,
        64'h72617020_79646165,
        64'h726c6120_64726143,
        64'h00000000_000a7367,
        64'h6e697474_65732079,
        64'h74696c69_6261696c,
        64'h65722065_74697277,
        64'h206e6f69_74697472,
        64'h61702064_656c6c6f,
        64'h72746e6f_63207473,
        64'h6f682074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000a29_7525203e,
        64'h20752528_206d756d,
        64'h6978616d_20736465,
        64'h65637865_20657a69,
        64'h73206465_636e6168,
        64'h6e65206c_61746f54,
        64'h00000000_0000000a,
        64'h65747562_69727474,
        64'h61206465_636e6168,
        64'h6e652074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0a64656e,
        64'h67696c61_20657a69,
        64'h73207075_6f726720,
        64'h50572043_4820746f,
        64'h6e206e6f_69746974,
        64'h72617020_69255047,
        64'h0000000a_64656e67,
        64'h696c6120_657a6973,
        64'h2070756f_72672050,
        64'h57204348_20746f6e,
        64'h20616572_61206465,
        64'h636e6168_6e652061,
        64'h74616420_72657355,
        64'h00000a65_7a697320,
        64'h70756f72_67205057,
        64'h20434820_656e6966,
        64'h65642074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_000a676e,
        64'h696e6f69_74697472,
        64'h61702074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0000000a,
        64'h61657261_20617461,
        64'h64207265_73752064,
        64'h65636e61_686e6520,
        64'h726f6620_64657269,
        64'h75716572_20342e34,
        64'h203d3e20_434d4d65,
        64'h00000000_000a2978,
        64'h6c257830_2878616d,
        64'h20736465_65637865,
        64'h20786c25_78302072,
        64'h65626d75_6e206b63,
        64'h6f6c6220_3a434d4d,
        64'h00000000_00000a64,
        64'h6d632070_6f747320,
        64'h646e6573_206f7420,
        64'h6c696166_20636d6d,
        64'h00000000_000a7964,
        64'h61657220_64726163,
        64'h20676e69_74696177,
        64'h2074756f_656d6954,
        64'h0000000a_58383025,
        64'h7830203a_726f7272,
        64'h45207375_74617453,
        64'h00000000_65646f6d,
        64'h206e776f_6e6b6e55,
        64'h00000000_00006473,
        64'h5f637369_72776f6c,
        64'h00000078_25782520,
        64'h00000020_3a78250a,
        64'h00000000_0a732574,
        64'h69622d64_25203a68,
        64'h74646957_20737542,
        64'h00000000_0000203a,
        64'h79746963_61706143,
        64'h00000000_00000a73,
        64'h25203a79_74696361,
        64'h70614320_68676948,
        64'h00000a64_25203a64,
        64'h65657053_20737542,
        64'h00000000_00000a20,
        64'h63256325_63256325,
        64'h6325203a_656d614e,
        64'h00000000_00000000,
        64'h0a782520_3a4d454f,
        64'h00000000_0a782520,
        64'h3a444920_72657275,
        64'h74636166_756e614d,
        64'h00000000_000a7325,
        64'h203a6563_69766544,
        64'h00202020_3a434d4d,
        64'h00000000_52444420,
        64'h00000000_00006f4e,
        64'h00000000_00736559,
        64'h0000000a_7825203d,
        64'h2074736f_68202c78,
        64'h25207461_20646574,
        64'h61657263_20636d6d,
        64'h00000000_00000a64,
        64'h25206f74_20646567,
        64'h6e616863_206b7361,
        64'h6d202c64_65747265,
        64'h736e6920_64726143,
        64'h00000000_0000000a,
        64'h6425206f_74206465,
        64'h676e6168_63206b73,
        64'h616d202c_6465766f,
        64'h6d657220_64726143,
        64'h000a7475_6f656d69,
        64'h74207325_203a6473,
        64'h5f637369_72776f6c,
        64'h00726464_615f6573,
        64'h61625f64_73203d3d,
        64'h20657361_625f6473,
        64'h00000000_00000063,
        64'h2e636d6d_5f637369,
        64'h72776f6c_2f637273,
        64'h00000000_00000000,
        64'h66656463_62613938,
        64'h37363534_33323130,
        64'h007f7c5d_5b3f3e3d,
        64'h3c3b3a2e_2c2b2a22,
        64'h00007f7c_5d5b3f3e,
        64'h3d3c3b3a_2c2b2a22,
        64'h0000000a_2e783230,
        64'h253a7832_30253a78,
        64'h3230253a_78323025,
        64'h3a783230_253a7832,
        64'h3025203d_20737365,
        64'h72646461_2043414d,
        64'h00000a78_6c253a78,
        64'h6c25203d_2043414d,
        64'h00000000_00000a78,
        64'h25203d20_5d64255b,
        64'h4d454f20_49505351,
        64'h000a7264_64612043,
        64'h414d2070_75746553,
        64'h0000000a_21747075,
        64'h72726574_6e692064,
        64'h656c646e_61686e75,
        64'h00000000_00000a78,
        64'h25783020_3d206570,
        64'h79745f6f_746f7270,
        64'h00000000_0a297825,
        64'h28206465_74726f70,
        64'h7075736e_75203d20,
        64'h6f746f72_70205049,
        64'h000a5741_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a534c50_4d203d20,
        64'h6f746f72_50205049,
        64'h00000000_000a4554,
        64'h494c5044_55203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505443_53203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a504d4f_43203d20,
        64'h6f746f72_50205049,
        64'h00000000_0000004d,
        64'h00000000_0000000a,
        64'h5041434e_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000a48,
        64'h50544545_42203d20,
        64'h6f746f72_50205049,
        64'h000a5054_4d203d20,
        64'h6f746f72_50205049,
        64'h00000a48_41203d20,
        64'h6f746f72_50205049,
        64'h000a5053_45203d20,
        64'h6f746f72_50205049,
        64'h000a4552_47203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505653_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000036,
        64'h00000000_00000000,
        64'h0a504343_44203d20,
        64'h6f746f72_50205049,
        64'h00000a50_54203d20,
        64'h6f746f72_50205049,
        64'h000a5044_49203d20,
        64'h6f746f72_50205049,
        64'h000a3a73_746e6574,
        64'h6e6f6320_74736574,
        64'h0000000a_3a726564,
        64'h61656820_74736574,
        64'h000a5055_50203d20,
        64'h6f746f72_50205049,
        64'h000a5047_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000054,
        64'h00000000_00000000,
        64'h0a504950_49203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000047,
        64'h00006425_2b544553,
        64'h46464f5f_524c5052,
        64'h00000000_3f3f3f3f,
        64'h00000000_00544553,
        64'h46464f5f_524c5052,
        64'h00000000_00544553,
        64'h46464f5f_44414252,
        64'h00000000_00005445,
        64'h5346464f_5f525352,
        64'h00000000_00544553,
        64'h46464f5f_53434652,
        64'h00544553_46464f5f,
        64'h4c525443_4f49444d,
        64'h00000000_00544553,
        64'h46464f5f_53434654,
        64'h00000000_00544553,
        64'h46464f5f_524c5054,
        64'h00000000_54455346,
        64'h464f5f49_4843414d,
        64'h00000000_54455346,
        64'h464f5f4f_4c43414d,
        64'h00000000_000a3b29,
        64'h78257830_2c302c78,
        64'h25287465_736d656d,
        64'h00000000_0a3b2978,
        64'h2578302c_78257830,
        64'h2c782528_6e666c65,
        64'h00000a70_2520726f,
        64'h72726520_7974696e,
        64'h61732072_64646170,
        64'h00000020_3a5d6425,
        64'h5b6e6f69_74636553,
        64'h000a7325_20202020,
        64'h00786c6c_2a302520,
        64'h00003a78_6c383025,
        64'h00732542_69632520,
        64'h00000000_00732573,
        64'h65747942_20756c25,
        64'h0073257a_48632520,
        64'h00000000_646c252e,
        64'h00000000_00756c25,
        64'h00000000_00000000,
        64'h73257a48_20756c25,
        64'h00000000_00007325,
        64'h00000000_00732520,
        64'h3a646c69_7542202c,
        64'h00000000_73257325,
        64'h00000000_00000a0a,
        64'h00000058_32302520,
        64'h00000000_0000002e,
        64'h00000000_00006325,
        64'h00000000_00000020,
        64'h20202020_20202020,
        64'h000a5245_46464f5f,
        64'h50434844_20726f66,
        64'h20676e69_74696157,
        64'h00000a73_25203a73,
        64'h25206563_69766564,
        64'h206e6f20_59524556,
        64'h4f435349_44205043,
        64'h48442064_6e657320,
        64'h74276e64_6c756f43,
        64'h000a5832_30253a58,
        64'h3230253a_58323025,
        64'h3a583230_253a5832,
        64'h30253a58_32302520,
        64'h3a204341_4d207325,
        64'h00000000_30687465,
        64'h00000000_000a2973,
        64'h2528726f_72726570,
        64'h000a5952_45564f43,
        64'h5349445f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_0000000a,
        64'h64252065_646f6370,
        64'h6f205043_48442064,
        64'h656c646e_61686e55,
        64'h00000000_0a642520,
        64'h6e6f6974_706f2064,
        64'h656c646e_61686e75,
        64'h00000000_0000000a,
        64'h73252072_6f727245,
        64'h00000000_00000a64,
        64'h65737566_65722073,
        64'h73657264_64612064,
        64'h65747365_75716552,
        64'h00000000_0000000a,
        64'h4b414e20_50434844,
        64'h00000000_0a444550,
        64'h50494b53_204b4341,
        64'h000a2273_2522203d,
        64'h20656d61_6e74736f,
        64'h4820746e_65696c43,
        64'h00000a22_73252220,
        64'h3d206e69_616d6f44,
        64'h00000000_0000000a,
        64'h7364253a_6d64253a,
        64'h68642520_3d20656d,
        64'h69742065_7361654c,
        64'h000a6425_2e64252e,
        64'h64252e64_2520203a,
        64'h73736572_64646120,
        64'h6b73616d_2074654e,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h61207265_74756f52,
        64'h00000000_00000000,
        64'h0a64252e_64252e64,
        64'h252e6425_20203a73,
        64'h73657264_64412050,
        64'h49207265_76726553,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h41205049_20746e65,
        64'h696c4320_50434844,
        64'h00000000_0000000a,
        64'h4b434120_50434844,
        64'h0000000a_54534555,
        64'h5145525f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_00000000,
        64'h0a702520_2c726f72,
        64'h7265206c_616e7265,
        64'h746e6920_70636864,
        64'h00000a29_73252c73,
        64'h25287075_6b6f6f6c,
        64'h000a6563_69766564,
        64'h206e776f_6e6b6e75,
        64'h00000000_203a6425,
        64'h20656369_7665440a,
        64'h00203a64_25206563,
        64'h69766564_2073250a,
        64'h00000000_00203a64,
        64'h25206563_69766544,
        64'h00000000_00000000,
        64'h73736572_6464612d,
        64'h63616d2d_6c61636f,
        64'h6c006874_6469772d,
        64'h6f692d67_65720074,
        64'h66696873_2d676572,
        64'h00737470_75727265,
        64'h746e6900_746e6572,
        64'h61702d74_70757272,
        64'h65746e69_00646565,
        64'h70732d74_6e657272,
        64'h75630076_65646e2c,
        64'h76637369_72007974,
        64'h69726f69_72702d78,
        64'h616d2c76_63736972,
        64'h0073656d_616e2d67,
        64'h65720064_65646e65,
        64'h7478652d_73747075,
        64'h72726574_6e690073,
        64'h65676e61_7200656c,
        64'h646e6168_702c7875,
        64'h6e696c00_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h00100000_00000000,
        64'h00000044_00000000,
        64'h67000000_10000000,
        64'h03000000_00000064,
        64'h6e727768_2d637369,
        64'h72776f6c_1b000000,
        64'h0e000000_03000000,
        64'h00003030_30303030,
        64'h34344064_6e727768,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h00800000_00000000,
        64'h00000043_00000000,
        64'h67000000_10000000,
        64'h03000000_00007fe3,
        64'h023e1800_47010000,
        64'h06000000_03000000,
        64'h03000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303334,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_00636d6d,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_02000000,
        64'h25010000_04000000,
        64'h03000000_02000000,
        64'h14010000_04000000,
        64'h03000000_00000100,
        64'h00000000_00000042,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00000000_30303030,
        64'h30303234_40636d6d,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h04000000_3a010000,
        64'h04000000_03000000,
        64'h02000000_30010000,
        64'h04000000_03000000,
        64'h01000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h00c20100_06010000,
        64'h04000000_03000000,
        64'h80f0fa02_4b000000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000041_00000000,
        64'h67000000_10000000,
        64'h03000000_00303537,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00000030_30303030,
        64'h30313440_74726175,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000000,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'hffff0000_01000000,
        64'hca000000_08000000,
        64'h03000000_00333130,
        64'h2d677562_65642c76,
        64'h63736972_1b000000,
        64'h10000000_03000000,
        64'h00003040_72656c6c,
        64'h6f72746e_6f632d67,
        64'h75626564_01000000,
        64'h02000000_02000000,
        64'hbb000000_04000000,
        64'h03000000_02000000,
        64'hb5000000_04000000,
        64'h03000000_03000000,
        64'hfb000000_04000000,
        64'h03000000_07000000,
        64'he8000000_04000000,
        64'h03000000_00000004,
        64'h00000000_0000000c,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h09000000_01000000,
        64'h0b000000_01000000,
        64'hca000000_10000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00000c00,
        64'h00000000_00000002,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_01000000,
        64'h03000000_01000000,
        64'hca000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6e696c63,
        64'h01000000_c3000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000008_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h01000000_bb000000,
        64'h04000000_03000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00007663_73697200,
        64'h656e6169_7261202c,
        64'h7a687465_1b000000,
        64'h13000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h31344074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha8060000_59010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'he0060000_38000000,
        64'h39080000_edfe0dd0,
        64'h00000000_fffff994,
        64'hfffff95a_fffff982,
        64'hfffff95a_fffff970,
        64'hfffff95c_fffff948,
        64'h00000000_64726143,
        64'h2d445320_726f6620,
        64'h746f6f62_2d752064,
        64'h6573696d_696e696d,
        64'h20435349_52776f4c,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00020000_00010000,
        64'h0000c000_00008000,
        64'h00006000_00004000,
        64'h00002000_00001000,
        64'h00000800_00000400,
        64'h00000200_00000100,
        64'h00000080_00000040,
        64'h00000020_00000000,
        64'h0bebc200_0c65d400,
        64'h02faf080_05f5e100,
        64'h02faf080_017d7840,
        64'h03197500_03197500,
        64'h02faf080_018cba80,
        64'h017d7840_017d7840,
        64'h00989680_000f4240,
        64'h000186a0_00002710,
        64'h50463c37_322d2823,
        64'h1e19140f_0d0c0a00,
        64'h00000000_00000000,
        64'h00000000_10000000,
        64'h00000001_00000000,
        64'h20000000_00000002,
        64'h00000000_40000000,
        64'h00000005_00000001,
        64'h20000000_00000006,
        64'h00000001_40000000,
        64'h70000000_00000000,
        64'h70000000_00000002,
        64'h70000000_00000004,
        64'h60000000_00000005,
        64'h30000000_00000001,
        64'h30000000_00000003,
        64'h00000000_40050100,
        64'h40050000_40040500,
        64'h40040401_40040400,
        64'h40040300_40040200,
        64'h40040100_40040000,
        64'h00000000_87feb560,
        64'h00000000_87feb548,
        64'h00000000_87feb530,
        64'h00000000_87feb518,
        64'h00000000_87feb500,
        64'h00000000_87feb4e8,
        64'h00000000_87feb4d0,
        64'h00000000_87feb4b8,
        64'h00000000_87feb4a0,
        64'h00000000_87feb488,
        64'h00000000_87feb478,
        64'h00000000_87feb468,
        64'hffffb988_ffffb988,
        64'hffffb988_ffffb988,
        64'hffffb984_ffffb980,
        64'hffffb980_ffffb95a,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_87fe4d0e,
        64'h00000000_87fe4ab0,
        64'h00000000_87fe4ea2,
        64'h00646374_65675f63,
        64'h6d6d5f64_72616f62,
        64'h00000002_0000ffff,
        64'h004c4b40_004c4b40,
        64'h00300000_20000000,
        64'h00000000_87fe9e88,
        64'h00000000_87feb150,
        64'h00717269_5f646e65,
        64'h5f617461_645f6473,
        64'h5f637369_72776f6c,
        64'h00000000_00007172,
        64'h695f646d_635f6473,
        64'h5f637369_72776f6c,
        64'h00007172_695f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0067616c,
        64'h665f7470_75727265,
        64'h746e695f_74696177,
        64'h5f637369_72776f6c,
        64'h00000000_646d635f,
        64'h74726174_735f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0000006e,
        64'h655f7172_695f6473,
        64'h00000000_00007475,
        64'h6f656d69_745f6473,
        64'h00000000_0000657a,
        64'h69736b6c_625f6473,
        64'h00000000_00000074,
        64'h6e636b6c_625f6473,
        64'h00000000_00000000,
        64'h74657365_725f6473,
        64'h00000000_74726174,
        64'h735f646d_635f6473,
        64'h00000000_0000676e,
        64'h69747465_735f6473,
        64'h00000000_00007669,
        64'h645f6b6c_635f6473,
        64'h00000000_00000000,
        64'h6e67696c_615f6473,
        64'h00000000_00006465,
        64'h6c5f7465_735f6473,
        64'h5f637369_72776f6c,
        64'h09020b04_0d060f08,
        64'h010a030c_050e0700,
        64'h020f0c09_0603000d,
        64'h0a070401_0e0b0805,
        64'h0c07020d_08030e09,
        64'h040f0a05_000b0601,
        64'heb86d391_2ad7d2bb,
        64'hbd3af235_f7537e82,
        64'h4e0811a1_a3014314,
        64'hfe2ce6e0_6fa87e4f,
        64'h85845dd1_ffeff47d,
        64'h8f0ccc92_655b59c3,
        64'hfc93a039_ab9423a7,
        64'h432aff97_f4292244,
        64'hc4ac5665_1fa27cf8,
        64'he6db99e5_d9d4d039,
        64'h04881d05_d4ef3085,
        64'heaa127fa_289b7ec6,
        64'hbebfbc70_f6bb4b60,
        64'h4bdecfa9_a4beea44,
        64'hfde5380c_6d9d6122,
        64'h8771f681_fffa3942,
        64'h8d2a4c8a_676f02d9,
        64'hfcefa3f8_a9e3e905,
        64'h455a14ed_f4d50d87,
        64'hc33707d6_21e1cde6,
        64'he7d3fbc8_d8a1e681,
        64'h02441453_d62f105d,
        64'he9b6c7aa_265e5a51,
        64'hc040b340_f61e2562,
        64'h49b40821_a679438e,
        64'hfd987193_6b901122,
        64'h895cd7be_ffff5bb1,
        64'h8b44f7af_698098d8,
        64'hfd469501_a8304613,
        64'h4787c62a_f57c0faf,
        64'hc1bdceee_242070db,
        64'he8c7b756_d76aa478,
        64'h02020202_02020202,
        64'h10020202_02020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02010101_01010101,
        64'h10010101_01010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h08101010_10020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02424242_42424210,
        64'h10101010_10010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h01414141_41414110,
        64'h10101010_10100404,
        64'h04040404_04040404,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h08080808_08080808,
        64'h08080808_08080808,
        64'h08082828_28282808,
        64'h08080808_08080808,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h0000bf5d_b8fff0ef,
        64'hd73fb0ef_0f450513,
        64'h00002517_b7e1c94f,
        64'h80efd85f_b0ef0f65,
        64'h05130000_2517bfe9,
        64'hab7ff0ef_d97fb0ef,
        64'h0f850513_00002517,
        64'hb7f5edbf_f0ef8522,
        64'hdabfb0ef_0fc50513,
        64'h00002517_a001929f,
        64'he0ef8522_dbffb0ef,
        64'h10050513_00002517,
        64'h878297ba_439c97ba,
        64'h078a6ca7_07130000,
        64'h071702f7_64634719,
        64'h0054579b_0ff47413,
        64'hfd391be3_deffb0ef,
        64'h25818552_688c0004,
        64'hb823dfdf_b0ef8622,
        64'h24012581_6080608c,
        64'he09c0905_85560007,
        64'hc7830169_07b34991,
        64'h140a0a13_00002a17,
        64'h130a8a93_00002a97,
        64'h440004b7_2f4b0b13,
        64'h00002b17_4901c16f,
        64'h80effe94_16e3e41f,
        64'hb0ef0405_854a0004,
        64'h059b6390_078e0134,
        64'h07b34495_15490913,
        64'h00002917_088009b7,
        64'h4401fb4f_e0ef1565,
        64'h05130000_2517f8ef,
        64'he0efe05a_e456e852,
        64'hec4ef04a_f426f822,
        64'hfc067139_fd6fe06f,
        64'h21850513_00002517,
        64'h9cffe06f_014160a2,
        64'he9bfb06f_0141d065,
        64'h05130000_251740a0,
        64'h05b360a2_00055c63,
        64'hbabf70ef_f3050513,
        64'h00000517_ebffb0ef,
        64'he406d125_05130000,
        64'h25171141_bf612441,
        64'hed3fb0ef_855aff54,
        64'h92e3eddf_b0ef8552,
        64'hd9fff0ef_24854589,
        64'h0007c503_97ce9381,
        64'h17820094_07bb4481,
        64'hefbfb0ef_8552dbdf,
        64'hf0ef8522_45a1b745,
        64'h00fb3023_04a19381,
        64'h178200c4_579b2421,
        64'he0bff0ef_85a68082,
        64'h61616b42_6ae27a02,
        64'h79a27942_74e26406,
        64'h60a60324_6863ec6b,
        64'h0b130000_2b174ac1,
        64'h338a0a13_00001a17,
        64'h4401d9ff_d0ef8526,
        64'h002c9201_16024089,
        64'h063be4df_f0ef002c,
        64'h05446363_0154053b,
        64'h44000b37_ff860a1b,
        64'h440184aa_89328aae,
        64'h89aae486_e85aec56,
        64'hf052f44e_f84afc26,
        64'he0a2715d_80826125,
        64'h7aa27a42_79e26906,
        64'h64a66446_60e6fa1f,
        64'hb0eff325_05130000,
        64'h2517ff24_91e3fb1f,
        64'hb0ef854e_e73ff0ef,
        64'h24854589_ff87c503,
        64'h97ba9381_10181782,
        64'h009407bb_49213c69,
        64'h89930000_19974481,
        64'hfdbfb0ef_3d450513,
        64'h00001517_ea3ff0ef,
        64'h45a1854a_feffb0ef,
        64'hf8050513_00002517,
        64'hff4992e3_ffffb0ef,
        64'h8556ec1f_f0ef2985,
        64'h45890007_c50397a6,
        64'h93811782_013407bb,
        64'h4a21412a_8a930000,
        64'h1a974981_826fc0ef,
        64'h42050513_00001517,
        64'heefff0ef_854a45a1,
        64'h83afc0ef_fcc50513,
        64'h00002517_ff4991e3,
        64'h84afc0ef_8556f0df,
        64'hf0ef2985_4589ff07,
        64'hc50397ba_93811018,
        64'h17820134_07bb4a21,
        64'h460a8a93_00001a97,
        64'h4981874f_c0ef46e5,
        64'h05130000_1517f3df,
        64'hf0ef854a_45a1feb7,
        64'h90e30705_06850605,
        64'h37e10107_002300f5,
        64'h58330106_802300f9,
        64'hd8330106_002300fa,
        64'h583355e1_03800793,
        64'h083886a6_0810f31f,
        64'hf0ef454d_89aa4589,
        64'h46010034_f3fff0ef,
        64'h454d8a2a_45894601,
        64'h0034f4df_f0eff456,
        64'hf852fc4e_ec86c63e,
        64'hc43a454d_842a4589,
        64'h460184ae_0034e4a6,
        64'he8a20587_e7938f55,
        64'h0089179b_0189571b,
        64'h30068693_00a7893b,
        64'h6685e0ca_004007b7,
        64'h711da1ff_e06f0141,
        64'h60a26402_00044503,
        64'h943e3fa7_87930000,
        64'h2797883d_febff0ef,
        64'h250135fd_0045551b,
        64'h00b7d863_842a4785,
        64'he406e022_1141bfe1,
        64'hf7100691_27850006,
        64'he6038082_73884400,
        64'h07b7ffe5_37fdc319,
        64'h8b097a98_440006b7,
        64'h3e800793_00b7ef63,
        64'h44000737_47812581,
        64'hf7888d51_440007b7,
        64'h0106161b_8d5d0085,
        64'h979b8082_25017b88,
        64'h440007b7_80822501,
        64'h6b880007_b8234400,
        64'h07b78082_25016388,
        64'h440007b7_8082e388,
        64'h440007b7_91011502,
        64'hbff1f5df_f0ef4541,
        64'hf63ff0ef_4521f69f,
        64'hf0ef4511_f6fff0ef,
        64'h4509f75f_f0ef4505,
        64'hf7bff0ef_4501e406,
        64'h1141bf51_c00028f3,
        64'hc02026f3_fac710e3,
        64'h9f2fc06f_48450513,
        64'h00002517_02a74733,
        64'h02a767b3_02b345bb,
        64'h02c74733_40000593,
        64'h02a68733_411686b3,
        64'h3e800513_c00026f3,
        64'h8e15c020_267302b7,
        64'h1d632705_fe0813e3,
        64'h97aa387d_00078023,
        64'h97aa0007_802397aa,
        64'h00078023_97aa0007,
        64'h80234000_081387f2,
        64'h45a901f6_1e134681,
        64'h48814701_00c5131b,
        64'h46058082_80826145,
        64'h69a26942_64e27402,
        64'h70a2ff24_17e3e6df,
        64'hf0ef2405_01358533,
        64'h46054685_008495b3,
        64'h497901f4_99934441,
        64'ha92fc0ef_44852265,
        64'h05130000_2517aa0f,
        64'hc0ef4ea5_05130000,
        64'h2517aacf_c0ef4c65,
        64'h05130000_2517ab8f,
        64'hc0ef4aa5_05130000,
        64'h25170400_0593c19f,
        64'he0efe44e_e84aec26,
        64'hf022f406_4ac50513,
        64'h00002517_7179bfa1,
        64'h0485ae4f_c0ef2765,
        64'h05130000_2517b7e9,
        64'h4a89af4f_c0ef4be5,
        64'h05130000_25179782,
        64'h852285ce_6642008a,
        64'h3783b0cf_c0ef4ce5,
        64'h05130000_2517c58d,
        64'h000a3583_02f74963,
        64'h6762010a_2783b28f,
        64'hc0ef856e_ed15920f,
        64'hf0ef8522_65a2b38f,
        64'hc0ef856a_85e6b40f,
        64'hc0ef8562_b46fc0ef,
        64'h855e85ca_00090663,
        64'hb52fc0ef_855a85a6,
        64'h80826149_7da27d42,
        64'h7ce26c06_6ba66b46,
        64'h6ae67a06_79a67946,
        64'h74e68556_640a60aa,
        64'hb7afc0ef_54c50513,
        64'h00002517_02997863,
        64'h068a0a13_00003a17,
        64'h558d8d93_00002d97,
        64'h558d0d13_00002d17,
        64'h550c8c93_00002c97,
        64'h550c0c13_00002c17,
        64'h550b8b93_00002b97,
        64'h550b0b13_00002b17,
        64'h44854a81_e43e99a2,
        64'h0034d793_e83e0014,
        64'hd9930044_d793bd8f,
        64'hc0efec36_e506f46e,
        64'hf86afc66_e0e2e4de,
        64'he8daecd6_f0d2f4ce,
        64'h56850513_00002517,
        64'h85aa962a_84ae842a,
        64'hfca6e122_fff58613,
        64'h8932f8ca_71758082,
        64'h6505b789_547dbf29,
        64'h0d85e73f_e0ef0007,
        64'hc50397ea_8b8d0007,
        64'h8b1b001b_079be87f,
        64'he0ef4521_ef91034d,
        64'hf7b300f6_932393c1,
        64'h17c20064_d78300f6,
        64'h922393c1_17c20044,
        64'hd78300f6_912393c1,
        64'h17c20024_d78300f6,
        64'h902393c1_17c20004,
        64'hd783e388_66c267e2,
        64'h16a7b823_00003797,
        64'h8d419101_14021502,
        64'h8c518d59_0106161b,
        64'h0105151b_67026622,
        64'hfdbfd0ef_e02afe1f,
        64'hd0efe42a_fe7fd0ef,
        64'h842afedf_d0efe836,
        64'hec3eb775_8c4a8bce,
        64'h4a858082_61497da2,
        64'h7d427ce2_6c066ba6,
        64'h6b466ae6_7a0679a6,
        64'h794674e6_640a60aa,
        64'h8522cd4f_c0ef6465,
        64'h05130000_2517020a,
        64'h8863e579_842aa82f,
        64'hf0ef854a_85ce866e,
        64'h059d9563_97de00fc,
        64'h06b3003d_97934d81,
        64'h8c4e8bca_9c4d0d13,
        64'h00003d17_9c4a0a13,
        64'h21048493_00003497,
        64'h4a81f73f_e0ef4b01,
        64'h8cb2f46e_e122e506,
        64'hf86afc66_e0e2e4de,
        64'he8daecd6_fca66a05,
        64'h02000513_89ae892a,
        64'hf0d2f4ce_f8ca7175,
        64'hbfa1547d_bf0d0d85,
        64'hfa9fe0ef_0007c503,
        64'h97e68b8d_00078a9b,
        64'h001a879b_fbdfe0ef,
        64'h4521ef91_0ba1033d,
        64'hf7b3ffa7_95e300d6,
        64'h00230ff6_f6930785,
        64'h00fb8633_0006c683,
        64'h018786b3_4781e288,
        64'h28a7b423_00003797,
        64'h8d4166e2_91011402,
        64'h15028c51_0106161b,
        64'h8d5d0105_151b6642,
        64'h67a28fcf_e0efe42a,
        64'h902fe0ef_e82a908f,
        64'he0ef842a_90efe0ef,
        64'hec36b775_8ba68b4a,
        64'h4a058082_61497da2,
        64'h7d427ce2_6c066ba6,
        64'h6b466ae6_7a0679a6,
        64'h794674e6_640a60aa,
        64'h8522df4f_c0ef7665,
        64'h05130000_2517020a,
        64'h0863ed45_842aba2f,
        64'hf0ef8526_85ca866e,
        64'h04fd9563_96da003d,
        64'h96936782_4d214d81,
        64'h8bca8b26_ae4c8c93,
        64'h00003c97_9c498993,
        64'h328c0c13_00003c17,
        64'h4a01892f_f0ef4a81,
        64'he032f46e_f86ae122,
        64'he506fc66_e0e2e4de,
        64'he8daecd6_f0d26985,
        64'h02000513_892e84aa,
        64'hf4cef8ca_fca67175,
        64'hb7e95b7d_b7490605,
        64'h00b83023_e30c85d6,
        64'he11185e2_00167513,
        64'h80826109_6de27d02,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e67906,
        64'h74a6855a_744670e6,
        64'hea2fc0ef_7ec50513,
        64'h00002517_fafb90e3,
        64'h04000793_2b85fbb4,
        64'h1be38c56_2405e931,
        64'h8b2ac5ef_f0ef854a,
        64'h85ce6622_ecefc0ef,
        64'h856a85da_ed6fc0ef,
        64'he4328552_06f61063,
        64'h974e00e9_08330036,
        64'h17136782_4601fffc,
        64'h4a93ef4f_c0ef8566,
        64'h85da0084_8b3bf00f,
        64'hc0ef8552_4401003b,
        64'h949b0177_9c334785,
        64'h4da17f2d_0d130000,
        64'h2d177eac_8c930000,
        64'h2c977e2a_0a130000,
        64'h2a17f2cf_c0ef4b81,
        64'he03289ae_f862e0da,
        64'he4d6f4a6_f8a2fc86,
        64'hec6ef06a_f466fc5e,
        64'he8d2ecce_7fc50513,
        64'h00002517_892af0ca,
        64'h7119bf75_5dfdbfc5,
        64'h85bafe08_1be385c6,
        64'hb7610605_e10ce28c,
        64'h85be0008_1363859a,
        64'h008bea63_00167813,
        64'h80826109_6de27d02,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e67906,
        64'h74a6856e_744670e6,
        64'hfa2fc0ef_8ec50513,
        64'h00003517_f8f41be3,
        64'h08000793_2405ed29,
        64'h8daad56f_f0ef8526,
        64'h85ca6622_fc6fc0ef,
        64'h856685a2_fcefc0ef,
        64'he432854e_05461c63,
        64'h96ca00d4_85330036,
        64'h16934601_fff7c313,
        64'hfff74893_8fd5008d,
        64'h16b300fd_17b30024,
        64'h079b8f5d_00ed1733,
        64'h00fd17b3_408b07bb,
        64'h408a873b_80ffc0ef,
        64'h856285a2_817fc0ef,
        64'h854e8fac_8c930000,
        64'h3c9703f0_0b930810,
        64'h0b134d05_07f00a93,
        64'h900c0c13_00003c17,
        64'h8f898993_00003997,
        64'h843fc0ef_44018a32,
        64'h892eec6e_fc86f06a,
        64'hf466f862_fc5ee0da,
        64'he4d6e8d2_eccef0ca,
        64'hf8a29125_05130000,
        64'h351784aa_f4a67119,
        64'hb7f15dfd_bfe5e19c,
        64'he31cbf61_0605e194,
        64'he314008c_66638082,
        64'h61096de2_7d027ca2,
        64'h7c427be2_6b066aa6,
        64'h6a4669e6_790674a6,
        64'h856e7446_70e68a9f,
        64'hc0ef9f25_05130000,
        64'h3517fb54_17e32405,
        64'he1398daa_e58ff0ef,
        64'h852685ca_66228c9f,
        64'hc0ef856a_85a28d1f,
        64'hc0efe432_85520566,
        64'h1a63974a_00e485b3,
        64'h00361713_4601fff6,
        64'hc693fff7_c7930089,
        64'h96b300f9_97b3408b,
        64'h87bb8fdf_c0ef8566,
        64'h85a2905f_c0ef8552,
        64'h08000a93_9ecd0d13,
        64'h00003d17_03f00c13,
        64'h498507f0_0b939eec,
        64'h8c930000_3c979e6a,
        64'h0a130000_3a17931f,
        64'hc0ef4401_8b32892e,
        64'hec6efc86_f06af466,
        64'hf862fc5e_e0dae4d6,
        64'he8d2ecce_f0caf8a2,
        64'ha0050513_00003517,
        64'h84aaf4a6_7119b7f1,
        64'h5dfdbfe5_e298e398,
        64'hbf610605_e28ce38c,
        64'h008c6663_80826109,
        64'h6de27d02_7ca27c42,
        64'h7be26b06_6aa66a46,
        64'h69e67906_74a6856e,
        64'h744670e6_997fc0ef,
        64'hae050513_00003517,
        64'hfb541be3_2405e139,
        64'h8daaf46f_f0ef8526,
        64'h85ca6622_9b7fc0ef,
        64'h856a85a2_9bffc0ef,
        64'he4328552_05661a63,
        64'h97ca00f4_86b30036,
        64'h17934601_008995b3,
        64'h00e99733_408b873b,
        64'h9e3fc0ef_856685a2,
        64'h9ebfc0ef_85520800,
        64'h0a93ad2d_0d130000,
        64'h3d1703f0_0c134985,
        64'h07f00b93_ad4c8c93,
        64'h00003c97_acca0a13,
        64'h00003a17_a17fc0ef,
        64'h44018b32_892eec6e,
        64'hfc86f06a_f466f862,
        64'hfc5ee0da_e4d6e8d2,
        64'heccef0ca_f8a2ae65,
        64'h05130000_351784aa,
        64'hf4a67119_bff159fd,
        64'hb74d0605_e29ce31c,
        64'h80826125_6c426be2,
        64'h7b027aa2_7a4279e2,
        64'h690664a6_854e6446,
        64'h60e6a6df_c0efbb65,
        64'h05130000_3517f94c,
        64'h19e30c05_e91d89aa,
        64'h81dff0ef_852285a6,
        64'h6622a8df_c0ef855e,
        64'h85cea95f_c0efe432,
        64'h854a0556_17639726,
        64'h00e406b3_00361713,
        64'h46018fd9_038c1713,
        64'h8fd9030c_17138fd9,
        64'h028c1713_8fd9020c,
        64'h17138fd9_018c1713,
        64'h0187e7b3_8fd9010c,
        64'h1793008c_1713ad9f,
        64'hc0ef855a_85ce000c,
        64'h099bae5f_c0ef854a,
        64'h10000a13_bccb8b93,
        64'h00003b97_bc4b0b13,
        64'h00003b17_bbc90913,
        64'h00003917_b07fc0ef,
        64'h4c018ab2_84aefc4e,
        64'hec86e862_ec5ef05a,
        64'hf456f852_e0cae4a6,
        64'hbd050513_00003517,
        64'h842ae8a2_711db7e1,
        64'h5d7db779_0605e198,
        64'he398872a_c291876a,
        64'h00167693_bf49000b,
        64'h3d038082_61656d42,
        64'h6ce27c02_7ba27b42,
        64'h7ae26a06_69a66946,
        64'h64e6856a_740670a6,
        64'hb6bfc0ef_cb450513,
        64'h00003517_fb441ae3,
        64'h2405e529_8d2a91bf,
        64'hf0ef8526_85ca6622,
        64'hb8bfc0ef_856685a2,
        64'hb93fc0ef_e432854e,
        64'h05561c63_97ca00f4,
        64'h85b30036_1793fffd,
        64'h45134601_baffc0ef,
        64'h856285a2_000bbd03,
        64'hcba50014_7793bc1f,
        64'hc0ef854e_04000a13,
        64'hca8c8c93_00003c97,
        64'hca0c0c13_00003c17,
        64'hfa8b8b93_00003b97,
        64'hfa8b0b13_00003b17,
        64'hca898993_00003997,
        64'hbf3fc0ef_44018ab2,
        64'h892ee86a_f486ec66,
        64'hf062f45e_f85afc56,
        64'he0d2e4ce_e8caf0a2,
        64'hcc050513_00003517,
        64'h84aaeca6_7159bfc1,
        64'h54fdbf59_0605e198,
        64'he3988726_c2918766,
        64'h00167693_80826165,
        64'h6ce27c02_7ba27b42,
        64'h7ae26a06_69a664e6,
        64'h69468526_740670a6,
        64'hc53fc0ef_d9c50513,
        64'h00003517_fb541be3,
        64'h2405e129_84aaa03f,
        64'hf0ef854a_85ce6622,
        64'hc73fc0ef_856285a2,
        64'hc7bfc0ef_e4328552,
        64'h05661863_97ce00f9,
        64'h05b30036_179314fd,
        64'h46014090_0cb3c99f,
        64'hc0ef8885_855e85a2,
        64'hfff44493_ca7fc0ef,
        64'h85520400_0a93d8ec,
        64'h0c130000_3c17d86b,
        64'h8b930000_3b97d7ea,
        64'h0a130000_3a17cc9f,
        64'hc0ef4401_8b3289ae,
        64'hec66eca6_f486f062,
        64'hf45ef85a_fc56e0d2,
        64'he4cef0a2_d9450513,
        64'h00003517_892ae8ca,
        64'h7159bfc9_070500a8,
        64'h3023e288_00f70533,
        64'ha9dff06f_6121863a,
        64'h69e2854e_790274a2,
        64'h70e27442_00c71c63,
        64'h96ae00d9_88330037,
        64'h16934701_8fc59081,
        64'h178265a2_66021482,
        64'h8fc18cc9_0109179b,
        64'h0105151b_887fe0ef,
        64'h84aa88df_e0ef892a,
        64'h893fe0ef_842a899f,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7f100e8,
        64'h30238f69_00083703,
        64'he3148ee9_07856314,
        64'hb15ff06f_6121863e,
        64'h69e2854e_790274a2,
        64'h70e27442_00c79c63,
        64'h974e00e5_88330037,
        64'h97134781_8d5d9101,
        64'h178265a2_66021502,
        64'h8fc18d45_0109179b,
        64'h0105151b_8fffe0ef,
        64'h84aa905f_e0ef892a,
        64'h90bfe0ef_842a911f,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7f100e8,
        64'h30238f49_00083703,
        64'he3148ec9_07856314,
        64'hb8dff06f_6121863e,
        64'h69e2854e_790274a2,
        64'h70e27442_00c79c63,
        64'h974e00e5_88330037,
        64'h97134781_8d5d9101,
        64'h178265a2_66021502,
        64'h8fc18d45_0109179b,
        64'h0105151b_977fe0ef,
        64'h84aa97df_e0ef892a,
        64'h983fe0ef_842a989f,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7d100e8,
        64'h302302a7_57330008,
        64'h3703e314_02a6d6b3,
        64'h07856314_4505e111,
        64'hc0dff06f_6121863e,
        64'h69e2854e_790274a2,
        64'h70e27442_00c79c63,
        64'h974e00e5_88330037,
        64'h97134781_8d5d9101,
        64'h178265a2_66021502,
        64'h8fc18d45_0109179b,
        64'h0105151b_9f7fe0ef,
        64'h84aa9fdf_e0ef892a,
        64'ha03fe0ef_842aa09f,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7e100e8,
        64'h302302a7_07330008,
        64'h3703e314_02a686b3,
        64'h07856314_c89ff06f,
        64'h6121863e_69e2854e,
        64'h790274a2_70e27442,
        64'h00c79c63_974e00e5,
        64'h88330037_97134781,
        64'h8d5d9101_178265a2,
        64'h66021502_8fc18d45,
        64'h0109179b_0105151b,
        64'ha73fe0ef_84aaa79f,
        64'he0ef892a_a7ffe0ef,
        64'h842aa85f_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7f100e8_30238f09,
        64'h00083703_e3148e89,
        64'h07856314_d01ff06f,
        64'h6121863e_69e2854e,
        64'h790274a2_70e27442,
        64'h00c79c63_974e00e5,
        64'h88330037_97134781,
        64'h8d5d9101_178265a2,
        64'h66021502_8fc18d45,
        64'h0109179b_0105151b,
        64'haebfe0ef_84aaaf1f,
        64'he0ef892a_af7fe0ef,
        64'h842aafdf_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7f100e8_30238f29,
        64'h00083703_e3148ea9,
        64'h07856314_d79ff06f,
        64'h6121863e_69e2854e,
        64'h790274a2_70e27442,
        64'h00c79c63_974e00e5,
        64'h88330037_97134781,
        64'h8d5d9101_178265a2,
        64'h66021502_8fc18d45,
        64'h0109179b_0105151b,
        64'hb63fe0ef_84aab69f,
        64'he0ef892a_b6ffe0ef,
        64'h842ab75f_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7ad0485_a9dff0ef,
        64'h0007c503_97e20039,
        64'hf7930985_aadff0ef,
        64'h4521ef81_00adb023,
        64'h00acb023_8d419101,
        64'h14021502_01a46433,
        64'h00a96533_010d1d1b,
        64'h0105151b_0344f7b3,
        64'hbcbfe0ef_892abd1f,
        64'he0ef8d2a_bd7fe0ef,
        64'h842abddf_e0efe33f,
        64'hf06f6165_7ae28556,
        64'h7b4264e6_85da8626,
        64'h6da26d42_6ce27c02,
        64'h7ba26a06_69a66946,
        64'h70a67406_8befd0ef,
        64'h23050513_00003517,
        64'h03749b63_00fb0cb3,
        64'h00fa8db3_00349793,
        64'h598c0c13_00003c17,
        64'h9c4a0a13_4981b3ff,
        64'hf0ef4481_8bb28b2e,
        64'he46ee86a_ec66e8ca,
        64'hf0a2f486_f062f45e,
        64'hf85ae4ce_eca60200,
        64'h05138aaa_6a05fc56,
        64'he0d27159_bfa507a1,
        64'h05858082_61256ca2,
        64'h6c426be2_7b027aa2,
        64'h7a4279e2_690664a6,
        64'h644660e6_557d938f,
        64'hd0ef2625_05130000,
        64'h3517944f_d0ef2365,
        64'h05130000_3517058e,
        64'h02e60d63_40e98733,
        64'h00359713_c689873e,
        64'h8a856390_008586b3,
        64'hbf5d07a1_04856398,
        64'he39840e9_87330034,
        64'h9713c689_873e8a85,
        64'h008486b3_a8894501,
        64'h98afd0ef_2d450513,
        64'h00003517_fd5417e3,
        64'h040502b4_9b634581,
        64'h87ca9a4f_d0ef8562,
        64'h85e69acf_d0ef8552,
        64'h03649863_448187ca,
        64'h9bafd0ef_855e85e6,
        64'h00040c9b_9c6fd0ef,
        64'h85524ac1_2acc0c13,
        64'h00003c17_fff94993,
        64'h2a8b8b93_00003b97,
        64'h2a0a0a13_00003a17,
        64'h9eafd0ef_44018b2e,
        64'he466e4a6_ec86e862,
        64'hec5ef05a_f456f852,
        64'hfc4ee8a2_2b450513,
        64'h00003517_892ae0ca,
        64'h711dbf5d_0785a001,
        64'ha1afd0ef_2b450513,
        64'h00003517_85a28626,
        64'ha2afd0ef_29c50513,
        64'h00003517_6090600c,
        64'h02e80363_60980004,
        64'h38038082_61054501,
        64'h64a26442_60e200c7,
        64'h986300d5_043300d5,
        64'h84b30037_96934781,
        64'he426e822_ec061101,
        64'hbbbff06f_80824501,
        64'h80824501_80828082,
        64'h80828082_45098082,
        64'h45098082_4509bff9,
        64'h26052004_04136622,
        64'he37fc0ef_e4328522,
        64'h85b28082_61454501,
        64'h64e27402_70a20096,
        64'h186300c6_84bb842e,
        64'hf406ec26_f0227179,
        64'h80824505_80824505,
        64'h80824505_80820141,
        64'h8d7d6402_60a29522,
        64'h408007b3_f57ff0ef,
        64'he406952e_842ae022,
        64'h1141a001_cbbff0ef,
        64'h4505aecf_d0efe406,
        64'h32850513_00003517,
        64'h85aa862e_86b28736,
        64'h11418082_02f55533,
        64'h47a9b000_25738082,
        64'h45018082_45018082,
        64'h01414501_60a2ee5f,
        64'hc0ef4200_0537b28f,
        64'hd0efe406_33c50513,
        64'h00003517_11418082,
        64'h80826105_644260e2,
        64'h8522944f_f0ef4581,
        64'h6622c509_842afd1f,
        64'hf0efe432_8532ec06,
        64'he8221101_02b50633,
        64'h8082953e_055e10d0,
        64'h0513e308_95360017,
        64'h86930075_6513157d,
        64'h631ce127_07130000,
        64'h47178082_45018082,
        64'h24050513_000f4537,
        64'ha001d69f_f0efe406,
        64'h25011141_90020000,
        64'h0023ee1f_f0ef8522,
        64'hb7813a25_05130000,
        64'h3517c511_2501cb9f,
        64'ha0ef4501_01c58593,
        64'h00003597_4605bfb9,
        64'h3a850513_00003517,
        64'hc5112501_b9afb0ef,
        64'hc4050513_00004517,
        64'hbe2fd06f_014124e5,
        64'h05130000_351760a2,
        64'h64024080_05b3cf81,
        64'h439ce9e7_87930000,
        64'h47970005_4863842a,
        64'h902f90ef_ea07a623,
        64'h00004797_ea07ac23,
        64'h00004797_e9850513,
        64'h00000517_c26fd0ef,
        64'h27850513_00003517,
        64'hb7e13fa5_05130000,
        64'h3517c511_2501d9bf,
        64'ha0efcaa5_05130000,
        64'h45174025_85930000,
        64'h35974605_c56fd0ef,
        64'h3f050513_00003517,
        64'hc62fd06f_014160a2,
        64'h64023e25_05130000,
        64'h3517c911_2501d79f,
        64'ha0efe022_e406f265,
        64'h05130000_45170e65,
        64'h85930000_35974605,
        64'h11418302_0141dae5,
        64'h85930000_259760a2,
        64'h64028322_f1402573,
        64'h0ff0000f_0000100f,
        64'hcb2fd0ef_e4063fe5,
        64'h05130000_3517842a,
        64'h85aae022_1141bf95,
        64'hf687a423_00004797,
        64'h9c25bf5d_320010ef,
        64'h854ede7f_f0ef0009,
        64'h4503993e_00397913,
        64'h42878793_00003797,
        64'h0009099b_00c4591b,
        64'he05ff0ef_4521b775,
        64'hfaf72223_00004717,
        64'h4785d0cf_d0ef42e5,
        64'h05130000_351785a6,
        64'h04967563_4632fca7,
        64'ha1230000_4797c50d,
        64'h2501814f_b0efd965,
        64'h05130000_451785ca,
        64'h86260074_fcf72e23,
        64'h00004717_57fd8082,
        64'h612169e2_790274a2,
        64'h744270e2_fea7ac23,
        64'h00004797_c10d2501,
        64'hf3afb0ef_dcc50513,
        64'h00004517_02b78563,
        64'h84b2842e_892aec4e,
        64'hfc06f04a_f426f822,
        64'h7139439c_02478793,
        64'h00004797_80826105,
        64'h60e2e9ff_f0ef0091,
        64'h4503ea7f_f0ef0081,
        64'h4503f13f_f0efec06,
        64'h002c1101_80826145,
        64'h694264e2_740270a2,
        64'hfe9410e3_ec9ff0ef,
        64'h00914503_ed1ff0ef,
        64'h34610081_4503f3ff,
        64'hf0ef0ff5_7513002c,
        64'h00895533_54e10380,
        64'h0413892a_f406e84a,
        64'hec26f022_71798082,
        64'h61456942_64e27402,
        64'h70a2fe94_10e3f0bf,
        64'hf0ef0091_4503f13f,
        64'hf0ef3461_00814503,
        64'hf81ff0ef_0ff57513,
        64'h002c0089_553b54e1,
        64'h4461892a_f406e84a,
        64'hec26f022_71798082,
        64'h61056442_60e2f43f,
        64'hf0ef0091_4503f4bf,
        64'hf0ef0081_4503fb7f,
        64'hf0ef0ff4_7513002c,
        64'hf5dff0ef_00914503,
        64'hf65ff0ef_00814503,
        64'hfd1ff0ef_ec068121,
        64'h842a002c_e8221101,
        64'h808200f5_802300e5,
        64'h80a30007_c7830007,
        64'h470397aa_973e8111,
        64'h00f57713_f4c78793,
        64'h00002797_b7f50405,
        64'hfa5ff0ef_80820141,
        64'h640260a2_e5090004,
        64'h4503842a_e406e022,
        64'h11418082_00e78823,
        64'h02000713_00e78423,
        64'hfc700713_00e78623,
        64'h470d0007_822300e7,
        64'h8023476d_00e78623,
        64'hf8000713_00078223,
        64'h410007b7_808200a7,
        64'h0023dfe5_0207f793,
        64'h01474783_41000737,
        64'h80820205_75130147,
        64'hc5034100_07b78082,
        64'h00054503_808200b5,
        64'h00238082_61056902,
        64'h64a26442_60e2f47d,
        64'hfa1ff0ef_41240433,
        64'h854a8926_0084f363,
        64'h89226804_8493842a,
        64'he04aec06_e8220098,
        64'h94b7e426_11018082,
        64'h61056902_64a26442,
        64'h60e2fe85_6ee3f45f,
        64'hf0ef0405_944a0285,
        64'h54332404_0413000f,
        64'h443702a4_85333e20,
        64'h00ef892a_f63ff0ef,
        64'h84aae04a_e426e822,
        64'hec061101_808202a7,
        64'hd5330141_91011502,
        64'h640260a2_02f407b3,
        64'h24078793_000f47b7,
        64'h414000ef_842af95f,
        64'hf0efe022_e4061141,
        64'h80826105_64a28d05,
        64'h02a7d533_644260e2,
        64'h91011502_02f407b3,
        64'h3e800793_440000ef,
        64'h842afc1f_f0ef84aa,
        64'he426e822_ec061101,
        64'h80824501_80820141,
        64'h8d5d9101_17821502,
        64'h60a21007_e78310a7,
        64'ha22310e1_a0232705,
        64'h1001a703_00e57763,
        64'h878e1041_e7035040,
        64'h00efe406_11418082,
        64'hcf3ff06f_e6458593,
        64'h00004597_4611cb81,
        64'h07c7d783_00004797,
        64'h80822401_01132201,
        64'h39032281_34832301,
        64'h34032381_3083f63f,
        64'hf0ef8522_002cea2f,
        64'hf0efe802_c44a0828,
        64'h20400613_85a6e60f,
        64'hf0ef2211_3c230028,
        64'h21800613_45818932,
        64'h84ae842a_23213023,
        64'h22913423_22813823,
        64'hdc010113_ebfff06f,
        64'h614505c1_70a24190,
        64'h7402d8bf_f06f6145,
        64'h70a265a2_74028522,
        64'h8a3fd0ef_e42e78e5,
        64'h05130000_3517842a,
        64'h8b3fd06f_61457b65,
        64'h05130000_351770a2,
        64'h740202e7_8a63470d,
        64'h00e78e63_01e15783,
        64'h00f10f23_0115c783,
        64'h00f10fa3_47090105,
        64'hc783f022_f4067179,
        64'h80826105_690264a2,
        64'h644260e2_d49ff06f,
        64'h61056902_64a260e2,
        64'h6442905f_d0ef7d65,
        64'h05130000_35170087,
        64'hcf63278d_439c1667,
        64'h87930000_479716f7,
        64'h19230000_47172785,
        64'h0007d783_18078793,
        64'h00004797_240000ef,
        64'h02000513_d1bff0ef,
        64'h45151965_d5830000,
        64'h45972560_00ef4535,
        64'he2bff0ef_854af9e5,
        64'h85930000_4597faa7,
        64'h94230000_47974611,
        64'hcf1ff0ef_1c055503,
        64'h00004517_faa79e23,
        64'h00004797_d05ff0ef,
        64'h4511dabf_f0ef0044,
        64'h8513ffc4_059b06a7,
        64'h9a632501_0024d783,
        64'hd21ff0ef_1f055503,
        64'h00004517_08a79563,
        64'h25010004_d783d37f,
        64'hf0ef84ae_450d892a,
        64'h08c7df63_8432478d,
        64'he04ae426_ec06e822,
        64'h1101b791_22f71023,
        64'h00004717_4785eb1f,
        64'hf0ef854e_02458593,
        64'h00004597_461102a7,
        64'h98230000_4797d77f,
        64'hf0ef4501_02a79e23,
        64'h00004797_d85ff0ef,
        64'h26f73023_00004717,
        64'h26f73023_00004717,
        64'h451107e2_08100793,
        64'ha1bfd0ef_8cc50513,
        64'h00004517_858a4390,
        64'h27878793_00004797,
        64'hdf2ff0ef_850a85a2,
        64'hdfaff0ef_850a8e65,
        64'h85930000_459700f7,
        64'h096302f0_07930129,
        64'h4703deaf_f0ef850a,
        64'h6b858593_00003597,
        64'h863ff0ef_850a4581,
        64'h10000613_b7552af7,
        64'h2f230000_47172000,
        64'h07938082_615569b2,
        64'h695264f2_741270b2,
        64'ha8bfd0ef_91450513,
        64'h00004517_00a405b3,
        64'hf24ff0ef_6fc50513,
        64'h00003517_842af32f,
        64'hf0ef8522_04a7f263,
        64'h0ff00793_9526f42f,
        64'hf0ef71a5_05130000,
        64'h351784aa_f50ff0ef,
        64'h852230a7_ad230000,
        64'h479704e7_ee631ff0,
        64'h0793fff5_071be93f,
        64'hf0ef9526_0505f72f,
        64'hf0ef8526_00a404b3,
        64'h0505f7ef_f0ef892e,
        64'hea4aee26_f6068522,
        64'h89aae64e_01258413,
        64'hf2227169_80824501,
        64'h80820141_640260a2,
        64'h557d0085_036386ef,
        64'ha0ef8432_e406e022,
        64'h11416680_006f6105,
        64'h64a260e2_6442b39f,
        64'hd06f6105_9a450513,
        64'h00004517_40a005b3,
        64'h64a260e2_64420005,
        64'h5e6384df_90efef65,
        64'h05130000_0517b61f,
        64'hd0ef9b25_05130000,
        64'h4517b6df_d0ef9a65,
        64'h05130000_45178622,
        64'h86aa608c_e63fc0ef,
        64'h85a26088_b87fd0ef,
        64'h85a29c11_ec069ae5,
        64'h05130000_45176380,
        64'he8226090_3f448493,
        64'h00004497_e4264067,
        64'h87930000_47971101,
        64'h80826105_64a26442,
        64'he00c95a6_60e2600c,
        64'ha15ff0ef_ec066008,
        64'h85aa84ae_862ee426,
        64'h43040413_00004417,
        64'he8221101_808242f7,
        64'h3f230000_471742f7,
        64'h3f230000_471707e2,
        64'h08100793_5000006f,
        64'h03050513_014160a2,
        64'h640202a4_753b4529,
        64'hfe7ff0ef_357d02b4,
        64'h55bb45a9_00b7f863,
        64'h47a500a0_4563842e,
        64'he406e022_1141bff9,
        64'h0505fd07_879b9fb9,
        64'h02f587bb_00d66763,
        64'h0ff6f693_fd07069b,
        64'h8082853e_e3190005,
        64'h470345a9_46254781,
        64'haa5ff06f_95be9201,
        64'h16029181_1582639c,
        64'h4b878793_00004797,
        64'h80820141_00e15503,
        64'h00a10723_812100a1,
        64'h07a31141_fa5ff06f,
        64'h4581d7df_f06f0141,
        64'h05054581_462960a2,
        64'h6402f77d_8b110007,
        64'h4703973e_00054703,
        64'hfea47ae3_157d8082,
        64'h0141557d_640260a2,
        64'he7198b11_00074703,
        64'h973efff5_85130267,
        64'h87930000_2797fff5,
        64'hc70300a4_05b395bf,
        64'hf0efe589_842ae406,
        64'he0221141_bfd50789,
        64'hbff1052a_052ab7e9,
        64'he01c078d_00e69863,
        64'h04200713_0027c683,
        64'hfce69fe3_052a0690,
        64'h07130017_c683fed7,
        64'h16e306b0_069302d7,
        64'h076304d0_06938082,
        64'h01416402_60a202d7,
        64'h0e630470_069300e6,
        64'hea6302d7_04630007,
        64'hc70304b0_0693601c,
        64'hf87ff0ef_842ee406,
        64'he0221141_b7e1e008,
        64'hb7cdfc97_879b0ff7,
        64'hf793fe07_079bc609,
        64'h8a09b7d1_96be0505,
        64'h02d586b3_feb7f4e3,
        64'hfd07879b_00088b63,
        64'h00467893_80826105,
        64'h85366442_60e2ec05,
        64'h00089863_04467893,
        64'h00064603_00f80633,
        64'h0007079b_00054703,
        64'h10080813_00002817,
        64'h468100c1_6583e0ff,
        64'hf0efc632_ec06006c,
        64'h842ee822_1101bfd5,
        64'h0789bff1_052a052a,
        64'hb7e9e01c_078d00e6,
        64'h98630420_07130027,
        64'hc683fce6_9fe3052a,
        64'h06900713_0017c683,
        64'hfed716e3_06b00693,
        64'h02d70763_04d00693,
        64'h80820141_640260a2,
        64'h02d70e63_04700693,
        64'h00e6ea63_02d70463,
        64'h0007c703_04b00693,
        64'h601cf0df_f0ef842e,
        64'he406e022_11418082,
        64'h014140a0_053360a2,
        64'hf23ff0ef_e4060505,
        64'h1141f2df_f06f00e6,
        64'h846302d0_07130005,
        64'h4683b7e9_4501e088,
        64'hfcf718e3_47a9fd27,
        64'h9be30785_8f81cb01,
        64'h0007c703_fe8782e3,
        64'h67e2f5df_f0ef8522,
        64'h082c892a_862e8082,
        64'h61217902_74a27442,
        64'h70e25529_e90165a2,
        64'hb0dff0ef_84b2842a,
        64'he42e0006_3023f04a,
        64'hfc06f426_f8227139,
        64'hb7e1e008_b7cdfc97,
        64'h879b0ff7_f793fe07,
        64'h079bc609_8a09b7d1,
        64'h96be0505_02d586b3,
        64'hfeb7f4e3_fd07879b,
        64'h00088b63_00467893,
        64'h80826105_85366442,
        64'h60e2ec05_00089863,
        64'h04467893_00064603,
        64'h00f80633_0007079b,
        64'h00054703_25480813,
        64'h00002817_468100c1,
        64'h6583f63f_f0efc632,
        64'hec06006c_842ee822,
        64'h1101bf6d_47a9bf7d,
        64'h47a18082_050900e7,
        64'h93630780_07130ff7,
        64'hf7930207_879bc709,
        64'h8b050007_4703973e,
        64'h29870713_00002717,
        64'h00154783_02f71663,
        64'h03000793_00054703,
        64'h02f71c63_47c14198,
        64'hc19c47c1_c3b10447,
        64'hf7930007_c78397ba,
        64'h00254703_04d71b63,
        64'h07800693_0ff77713,
        64'h0207071b_c6898a85,
        64'h0006c683_00e786b3,
        64'h2e878793_00002797,
        64'h00154703_08f71163,
        64'h03000793_00054703,
        64'he7a9419c_b7f1377d,
        64'h87aabfa5_fef51be3,
        64'h0785f8b7_12e30007,
        64'hc70300d8_0a630087,
        64'h85130007_b803bfcd,
        64'h367d0785_f8b71fe3,
        64'h0007c703_d24d8a1d,
        64'heb1187aa_27018edd,
        64'h00365713_02079693,
        64'h8fd90107_179300b7,
        64'he7330085_97938e1d,
        64'h953e9381_02071793,
        64'hfaf50785_36fdfcb8,
        64'h1ce30007_c80387aa,
        64'h0007069b_40e7873b,
        64'h47a1c31d_00757713,
        64'hb7f5367d_0785feb7,
        64'h1ce30007_c7038082,
        64'h853e4781_e60187aa,
        64'h260100c7_ef630ff5,
        64'hf59347c1_b7ed853e,
        64'hfeb70be3_00150793,
        64'h00054703_80824501,
        64'h00c51463_0ff5f593,
        64'h962abfe9_0405d175,
        64'hf8bff0ef_397d8522,
        64'h85ce8626_80826145,
        64'h69a26942_64e27402,
        64'h70a28522_44010099,
        64'h5b630005_091bd13f,
        64'hf0ef8522_c8890005,
        64'h049bd1ff_f0ef89ae,
        64'he84af406_e44eec26,
        64'h852e842a_f0227179,
        64'hbfc50505_feb78de3,
        64'h00054783_808200c5,
        64'h1363962a_b7dd0585,
        64'h0505fbed_9f990005,
        64'hc7030005_47838082,
        64'h853e4781_00c51563,
        64'h962ab7fd_00f68023,
        64'h16fd0005_c78315fd,
        64'hd7e500e5_87b340b6,
        64'h073300c5_06b395b2,
        64'h80820141_640260a2,
        64'h8522f57f_f0ef00a5,
        64'he963842a_e406e022,
        64'h11418082_614564e2,
        64'h69428526_740270a2,
        64'h00040023_f79ff0ef,
        64'h944a864a_8522fff6,
        64'h091300c5_64636582,
        64'h892ace11_84aa6622,
        64'hdcdff0ef_e02ee84a,
        64'hf406e432_ec26852e,
        64'h842af022_7179bf65,
        64'hfee78fa3_0785fff5,
        64'hc7030585_bfe1469d,
        64'h00c508b3_87aa872e,
        64'hbfc100e5_07b3963e,
        64'h95ba070e_02f707b3,
        64'h57e10036_5713ff06,
        64'he8e340f8_8833ff07,
        64'hbc2307a1_ff873803,
        64'h07218082_02c79e63,
        64'h963e87aa_cb9d8b9d,
        64'h00a5e7b3_00b50a63,
        64'hbf6dfeb7_8fa30785,
        64'hbfe1fef7_3c230721,
        64'hbfd10ff5_f6934725,
        64'hbfc1963a_97aa078e,
        64'h02e78733_57610036,
        64'h57930106_ef6340e8,
        64'h8833469d_00c508b3,
        64'h872aff6d_377d8fd5,
        64'h07a28082_04c79063,
        64'h963e87aa_cb9d0075,
        64'h77938082_4501b7e5,
        64'h078900d7_80a300e7,
        64'h80238082_e3110017,
        64'hc703ce81_0007c683,
        64'h87aacf99_00054783,
        64'hc11d8082_610564a2,
        64'h85266442_60e2e008,
        64'h05050005_0023c501,
        64'hf73ff0ef_8526842a,
        64'hc891e822_ec066104,
        64'he4261101_bfd988a7,
        64'hbb230000_57970505,
        64'h00050023_c7810005,
        64'h4783c519_f9fff0ef,
        64'h852285a6_80826105,
        64'h64a26442_60e28522,
        64'h44018c07_b1230000,
        64'h5797ef81_00044783,
        64'h942af9df_f0ef85a6,
        64'h8522cc11_63808de7,
        64'h87930000_5797e519,
        64'h842a84ae_ec06e426,
        64'he8221101_bfd587ae,
        64'hb7e50505_fafd0007,
        64'hc6830785_fee68fe3,
        64'h80824501_eb190005,
        64'h4703bff9_0785bfd5,
        64'h872e8082_fe081be3,
        64'h00074803_070500c8,
        64'h0a638082_ea1140d7,
        64'h85330007_c60387aa,
        64'h86aabfcd_872eb7d5,
        64'h0785fe08_1be30007,
        64'h48030705_fed80fe3,
        64'h8082ea99_40c78533,
        64'h0007c683_87aa862a,
        64'hb7fd0785_808240a7,
        64'h8533e701_0007c703,
        64'h00b78563_87aa95aa,
        64'h80826105_644260e2,
        64'h4501fe85_7be3157d,
        64'h00b78663_00054783,
        64'h0ff5f593_952265a2,
        64'hfe5ff0ef_ec06842a,
        64'he42ee822_1101bfcd,
        64'h07858082_40a78533,
        64'he7010007_c70387aa,
        64'hbfcd0505_dffd8082,
        64'h00b79363_00054783,
        64'h0ff5f593_80824501,
        64'hbfcd0505_c3998082,
        64'h00b79363_00054783,
        64'h0ff5f593_8082853e,
        64'hff790505_e3994187,
        64'hd79b0187_979b40f7,
        64'h07bbfff5_c7830005,
        64'h47030585_a8394781,
        64'h00c59463_962e8082,
        64'h853ef37d_0505e399,
        64'h4187d79b_0187979b,
        64'h40f707bb_fff5c783,
        64'h00054703_0585b7cd,
        64'h87ba8082_000780a3,
        64'h00c71563_8082e291,
        64'hfed70fa3_00178713,
        64'hfff5c683_0585963e,
        64'hfb7d0017_86930007,
        64'hc70387b6_8082e219,
        64'h87aab7d5_87b68082,
        64'hfb75fee7_8fa30785,
        64'hfff5c703_0585eb09,
        64'h00178693_0007c703,
        64'h87aa8082_fb65fee7,
        64'h8fa30785_fff5c703,
        64'h058500c7_896387aa,
        64'h962a8082_fb75fee7,
        64'h8fa30785_fff5c703,
        64'h058587aa_80820141,
        64'h640260a2_8d411502,
        64'h9001fd1f_f0ef1402,
        64'h0005041b_fdbff0ef,
        64'he022e406_11418082,
        64'h01412501_640260a2,
        64'h8d410105_151bfe9f,
        64'hf0ef842a_fefff0ef,
        64'he022e406_1141fc3f,
        64'hf06fae25_05130000,
        64'h55178082_25018d5d,
        64'h00f717bb_40f007b3,
        64'h00f7553b_93ed836d,
        64'h8f3d0127_d713e118,
        64'h97360017_671302d7,
        64'h86b36518_6294611c,
        64'h8a868693_00005697,
        64'h1bc0106f_80826105,
        64'h690264a2_644260e2,
        64'h8522e99f_f0ef10f4,
        64'h00230247_c7838522,
        64'h0ea42e23_681c18f4,
        64'h34232ae7_87930000,
        64'h179718f4_30232be7,
        64'h87930000_179716f4,
        64'h3c2391c7_8793ffff,
        64'hf797e65f_f0ef0405,
        64'h28230325_3023e904,
        64'h10f502a3_47850ef5,
        64'h2c234799_c57c57fd,
        64'hcd21842a_200010ef,
        64'h45051c00_059384aa,
        64'h892ec7ad_639cc7bd,
        64'h651ccbad_511ccbbd,
        64'h4d5ccfad_44014d1c,
        64'hc1414401_e04ae426,
        64'hec06e822_1101b771,
        64'h600032a0_10ef98e5,
        64'h05130000_451701a9,
        64'h8863da4f_e0ef8566,
        64'h85e20097_8e63601c,
        64'hdb2fe0ef_855e85ca,
        64'h00090663_dbefe0ef,
        64'h638c855a_0fc42603,
        64'h681c8956_0007c363,
        64'h89524c1c_c7914901,
        64'h541cddcf_e06f6125,
        64'h57050513_00004517,
        64'h6d026ca2_6c426be2,
        64'h7b027aa2_7a4279e2,
        64'h690664a6_60e66446,
        64'h02941563_4d29a06c,
        64'h8c930000_4c970005,
        64'h0c1b422b_8b930000,
        64'h4b97422b_0b130000,
        64'h4b1741aa_8a930000,
        64'h4a9742aa_0a130000,
        64'h4a1789aa_e0caec86,
        64'he06ae466_e862ec5e,
        64'hf05af456_f852fc4e,
        64'h6080e8a2_c6c48493,
        64'h00005497_e4a6711d,
        64'h8082e308_e518e11c,
        64'he7886798_c8478793,
        64'h00005797_e5088082,
        64'hb207a023_00005797,
        64'he79ce39c_c9c78793,
        64'h00005797_b7d56000,
        64'ha9cff0ef_8522c781,
        64'h19a44783_80826105,
        64'h64a26442_60e20094,
        64'h176384be_ec06e426,
        64'h6380e822_ccc78793,
        64'h00005797_11018082,
        64'h4388b6a7_87930000,
        64'h57978082_0f850513,
        64'h8082c398_0015071b,
        64'h4388b827_87930000,
        64'h5797bfd5_55358082,
        64'h610564a2_644260e2,
        64'he0800f84_0413e501,
        64'hcf0ff0ef_842acd09,
        64'hf7dff0ef_84aee822,
        64'hec06e426_1101bfcd,
        64'hf8400513_bfe54501,
        64'h80826105_60e25535,
        64'heb3fe06f_610560e2,
        64'h00f70c63_0ff00793,
        64'h08154703_02b70063,
        64'h65a21035_4703c105,
        64'hfbdff0ef_e42eec06,
        64'h11014148_8082853e,
        64'hbfd187b6_00a60463,
        64'h0fc7a603_80820141,
        64'h853e4781_60a2f60f,
        64'he0efe406_53c50513,
        64'h00004517_85aa1141,
        64'h02e79063_6394631c,
        64'hd9870713_00005717,
        64'h80824501_80820141,
        64'h45016402_60a20dc0,
        64'h00ef13e0_00ef02c0,
        64'h0513fc5f_f0ef8522,
        64'h00055563_aeefe0ef,
        64'h852212a0_00efdcf7,
        64'h25230000_5717842a,
        64'he406e022_47851141,
        64'hef9d439c_de078793,
        64'h00005797_808218b5,
        64'h0d238082_557d8082,
        64'h557d8082_4501c56c,
        64'he54ff06f_fa100413,
        64'hf0eff06f_2006061b,
        64'h40010637_f0a60963,
        64'h4505f0c5_43638ca6,
        64'h02e34509_8a3d01a6,
        64'hd61bf2c5_1a634000,
        64'h063706bb_a42306eb,
        64'ha22306fb_a02304db,
        64'hae23018b_a50345e6,
        64'h475647c6_46b6ea05,
        64'h1163842a_93bfe0ef,
        64'hc4be855e_0107979b,
        64'h008c4601_07cbd783,
        64'hc2be479d_04f11023,
        64'h47a506fb_9e2304e1,
        64'h57830007_d663018b,
        64'ha783ec05_1b63842a,
        64'h96ffe0ef_c2be47d5,
        64'h855ec4be_0107979b,
        64'h008c4601_07cbd783,
        64'h04f11023_478d6da0,
        64'h00ef06cb_851300ec,
        64'h4641bf6d_11872583,
        64'h974e8379_02079713,
        64'hfcfc65e3_4581b7c9,
        64'hf521d31f_e0ef855e,
        64'h45850b70_06130ff6,
        64'hf693bb91_fd319fdf,
        64'he0ef855e_cb0ff0ef,
        64'h855e4601_18fbae23,
        64'h08bba223_0017b793,
        64'h17ed088b_a583ef8d,
        64'h1afba823_409ce79d,
        64'h0046f793_00892683,
        64'hf941808f_f0ef855e,
        64'h408c933f_e0ef855e,
        64'h02ebaa23_0017b713,
        64'h41b787b3_01a78663,
        64'h471100d7_89634721,
        64'h400006b7_00092783,
        64'hbb6d925f_e0ef58e5,
        64'h05130000_4517f764,
        64'h9fe304a1_fb9911e3,
        64'h0931973f_e0ef855e,
        64'h035baa23_08fba223,
        64'h180bae23_1a0ba823,
        64'h088ba783_ddbfe0ef,
        64'h855e4585_0b700613,
        64'h4681c131_debfe0ef,
        64'h855e0fb6_f6934585,
        64'h0b700613_00894683,
        64'hc3a18ff9_00fa77b3,
        64'h00092703_40dc04f7,
        64'h18630017_b79317ed,
        64'h00494703_409c1000,
        64'h0db72000_0d3718e9,
        64'h09130000_3917cbb5,
        64'h278100fa_77b300fa,
        64'h97bb409c_1e0c8c93,
        64'h00003c97_4c2d1aeb,
        64'h0b130000_3b174a85,
        64'hdb4ff0ef_19c48493,
        64'h00003497_00fa7a33,
        64'h855e4601_088ba583,
        64'h044ba783_040baa03,
        64'h04fba023_00c7e793,
        64'h040ba783_c7998b85,
        64'h04eba023_01076713,
        64'h040ba703_04eba023,
        64'h0217071b_c68900c7,
        64'hf693ce91_0027f693,
        64'h1adba423_03f7f693,
        64'h0c46c783_04fba023,
        64'h0017079b_70000737,
        64'hbb956ba5_05130000,
        64'h4517e691_ecf76ce3,
        64'h1a0bb683_400407b7,
        64'h04fba023_27851000,
        64'h07b7b8d1_02fba423,
        64'h47857e40_10ef8526,
        64'ha3ffe0ef_8a3d8abd,
        64'h0146561b_0106569b,
        64'h06248513_73c58593,
        64'h00004597_074ba603,
        64'ha5ffe0ef_04d48513,
        64'h74058593_00004597,
        64'h26810ff7_77130ff8,
        64'h78130ff7_f7930188,
        64'h569b0108_571b0088,
        64'h579b06cb_c603077b,
        64'hc883070b_a803a95f,
        64'he0effef5_36230245,
        64'h05137625_85930000,
        64'h459784aa_06fbc603,
        64'h074bd683_07abd703,
        64'h02c7d7b3_ed109201,
        64'h0a8bb783_d11c9fb9,
        64'h071200e0_37338f75,
        64'h02071613_76c19fb5,
        64'h068e00d0_36b38ef9,
        64'hf0068693_ff0106b7,
        64'h9fb5068a_00d036b3,
        64'h8ef90f06_8693f0f0,
        64'hf6b79fb5_00f037b3,
        64'h068600d0_36b32781,
        64'h8ef98ff9_ccc68693,
        64'haaa78793_ccccd6b7,
        64'haaaab7b7_08cba703,
        64'h00050623_00051523,
        64'h484000ef_855e08fb,
        64'ha82308fb_a6232000,
        64'h0793c799_19cba783,
        64'h1afbaa23_1b0ba783,
        64'h0adba223_0afba023,
        64'h02d606bb_02f757bb,
        64'h8a8d0106_d69b02e6,
        64'h073b3e80_0613c305,
        64'hc38d03f7_77132781,
        64'h0126d71b_8fd10186,
        64'hd61b8ff9_17fd67c1,
        64'h00cca683_08fbae23,
        64'h0087171b_1487a783,
        64'h97b6078a_2ec68693,
        64'h00003697_04d61c63,
        64'h800306b7_018ba603,
        64'h00f6f863_8bbd00c7,
        64'h579b46a5_008ca703,
        64'hfdb59ee3_fefdae23,
        64'h8fd98ff5_8f510087,
        64'hd79b8e69_0087961b,
        64'h8f510187_971b0187,
        64'hd61b0d91_000da783,
        64'hf0068693_00ff0537,
        64'h040d8593_66c1b545,
        64'h11872583_974e8379,
        64'h02079713_eaf768e3,
        64'h4581472d_b35d04fb,
        64'ha0230087_6793da06,
        64'hd9e3040b_a70302e7,
        64'h96938fd1_8ff50087,
        64'hd79b0087_961bf006,
        64'h869366c1_44dcfbe1,
        64'h8b8583a5_4cdcd005,
        64'h1ce3d61f_e0efdc3e,
        64'hf84af426_c556855e,
        64'h010c0400_07931030,
        64'hc33e47d5_08f11023,
        64'h4799020a_08633a7d,
        64'h09053ac5_4a159881,
        64'h19020100_0ab70ff1,
        64'h04934905_bbc58003,
        64'h0737de07_5ee30307,
        64'h971300eb_ac238002,
        64'h0737b519_a007071b,
        64'h80011737_b61ddf40,
        64'h0413cbdf_e0ef9265,
        64'h05130000_5517e6f4,
        64'h9fe349a7_87930000,
        64'h379704a1_eafa94e3,
        64'h47a10a91_8c9ff0ef,
        64'h855e8405_85934601,
        64'h180bae23_096ba223,
        64'h1afba823_017d85b7,
        64'h4785f3ed_37fd6702,
        64'h67a20e05_0c63e0df,
        64'he0efe03a_c93ae552,
        64'he16ee43e_855e110c,
        64'h01100400_07134791,
        64'hd502d33a_0af11023,
        64'h47b56702_e915e35f,
        64'he0efd53e_e03ad33a,
        64'h8cee855e_110c0107,
        64'h979b4601_475507cb,
        64'hd7830af1_10230370,
        64'h0793fe07_fd930ff1,
        64'h0793947f_f0ef855e,
        64'h460118fb_ae2308bb,
        64'ha2230017_b79317ed,
        64'h088ba583_14079a63,
        64'h1afba823_409c09b7,
        64'h94638bbd_010c4783,
        64'he941e91f_e0efc93e,
        64'he552e162_855e110c,
        64'h04000793_0110d53e,
        64'h00fde7b3_17c12d81,
        64'h810007b7_d33e47d5,
        64'h0af11023_47994d85,
        64'h0ce79163_470d01a7,
        64'h8663409c_dfdfe0ef,
        64'h855e02fb_aa23001c,
        64'hb79340fc_8cb31000,
        64'h07b700ec_88634791,
        64'h20000737_00ec8d63,
        64'h47a14000_07370e05,
        64'h1c638daa_971ff0ef,
        64'h855e0015_b59340bc,
        64'h85b31000_05b700fc,
        64'h88634591_200007b7,
        64'h00fc8d63_45a14000,
        64'h07b71407_81630197,
        64'hf7b300f9_77b340dc,
        64'h0007ac83_97d6109c,
        64'h840b0b1b_4a81017d,
        64'h8b371607_85632781,
        64'h00f977b3_00e797bb,
        64'h47854098_0a05fe07,
        64'hfc1383f9_79130ff1,
        64'h079300f9_793361e4,
        64'h84930000_3497020d,
        64'h1a13044b_a783f0be,
        64'h4d05040b_a903639c,
        64'h23078793_00005797,
        64'h1ef71863_800107b7,
        64'h018ba703_04fba023,
        64'h8fd92000_0737040b,
        64'ha7830007_596302d7,
        64'h971300eb_ac238001,
        64'h073720d7_02634689,
        64'h21270063_8b3d0187,
        64'hd71b04eb_ac238f55,
        64'h8f718ecd_0087571b,
        64'h8de90087_159b8ecd,
        64'h0187169b_0187559b,
        64'h40d804fb_aa232781,
        64'h8fd58ef1_f0070613,
        64'h8fd16741_0087569b,
        64'h8e698fd5_0087161b,
        64'h0187179b_0187569b,
        64'h00ff0537_4098b555,
        64'h8b1d9381_00f7571b,
        64'h17828fd5_01e7569b,
        64'h8ff50027_979b16f1,
        64'h6685b54d_08bba823,
        64'h00b515bb_89bd0165,
        64'hd59bbd99_40030637,
        64'ha7a94002_0637bb45,
        64'h842afe0a_16e33a7d,
        64'hc131850f_f0efd05a,
        64'hec56e826_855e108c,
        64'h08104b21_0a854a11,
        64'hd48206f1_10239881,
        64'h02091a93_03300793,
        64'h0bf10493_4905d2ca,
        64'hed05880f_f0efd4be,
        64'hd2ca855e_0107979b,
        64'h108c4601_07cbd783,
        64'h06f11023_03700793,
        64'h04fba023_27891000,
        64'h07b75407_5a63018b,
        64'ha703e005_1fe3842a,
        64'hffbfe0ef_855e00b5,
        64'h45830f70_00ef855e,
        64'he2051ae3_842ac9af,
        64'hf0ef855e_08fb80a3,
        64'h57fd08fb_aa234785,
        64'he40516e3_842a8e4f,
        64'hf0efc4be_c2ca855e,
        64'h008c0107_979b4601,
        64'h495507cb_d78304f1,
        64'h1023479d_902ff0ef,
        64'hc282c4be_04e11023,
        64'h855e008c_46010107,
        64'h979b4711_00e78e63,
        64'h577d04cb_a783c215,
        64'h08fba823_00e7f463,
        64'h20000793_090ba703,
        64'h08fba623_0107d463,
        64'h20000793_0afbb823,
        64'h0e0bb023_0c0bbc23,
        64'h0c0bb823_0c0bb423,
        64'h0c0bb023_0a0bbc23,
        64'h030787b3_00e797b3,
        64'h07090785_47219381,
        64'h17828fd9_8ff50107,
        64'h571b003f_06b70107,
        64'h979b1406_8e6302cb,
        64'ha683090b_a8231408,
        64'hdc63090b_a62300d5,
        64'h183b8abd_0107d69b,
        64'h08dba223_08dba423,
        64'h04cba823_180bae23,
        64'h1a0ba823_8a0500c7,
        64'hd61b02d6_06bb018b,
        64'ha8834505_1086a683,
        64'h0f864603_96ce964e,
        64'h068a8a3d_80498993,
        64'h00004997_8a9d0036,
        64'hd61b00cb_ac234006,
        64'h061b4001_0637a029,
        64'h40040637_0ea61ee3,
        64'h45111aa6_0f63450d,
        64'hbf0506fb_9e234785,
        64'h02fba623_8b8541e7,
        64'hd79b048b_a78300fb,
        64'hac234000_07b7bfe9,
        64'h1d7010ef_06400513,
        64'h12a96ee3_149010ef,
        64'h85260007_cc63048b,
        64'ha783f155_842ab36f,
        64'hf0ef855e_45853e80,
        64'h09139081_02051493,
        64'h16d010ef_4501b16f,
        64'hf0ef855e_0407c163,
        64'h180b8c23_048ba783,
        64'h8082615d_6db66d56,
        64'h6cf67c16_7bb67b56,
        64'h7af66a1a_69ba695a,
        64'h64fa741a_70ba8522,
        64'hd55d842a_d99ff0ef,
        64'h855ea031_020ba423,
        64'hf4fd34fd_100503e3,
        64'h842aaa0f_f0ef855e,
        64'h008c4601_4495cf81,
        64'h8b851b8b_a7831205,
        64'h00e3842a_abaff0ef,
        64'hc482c2be_855e008c,
        64'h479d4601_04f11023,
        64'h4789e7b5_180b8ca3,
        64'h198bc783_c7b1199b,
        64'hc7831ff0_10ef4501,
        64'h8baae3b5_4401e6ee,
        64'heaeaeee6_f2e2f6de,
        64'hfadafed6_e352e74e,
        64'heb4aef26_f706f322,
        64'h7161551c_b58584aa,
        64'hb595fa10_0493a10f,
        64'hf0efe4a5_05130000,
        64'h5517d965_c1cff0ef,
        64'h85224585_bfd118f4,
        64'h0c234785_0007d663,
        64'h443ced09_c34ff0ef,
        64'h85224581_c04ff0ef,
        64'h852202f5_1f63f920,
        64'h0793b55d_18f40ca3,
        64'h47850604_1e23d45c,
        64'h8b8541e7_d79bc43c,
        64'hcc188001_073700e6,
        64'h85638002_07374c14,
        64'hbf453310_10ef3e80,
        64'h05130609_0863397d,
        64'h0007ca63_47b2ed1d,
        64'hb8eff0ef_8522858a,
        64'h4601c43e_0197e7b3,
        64'h01871563_c43e0177,
        64'hf7b3c25a_4bdc0151,
        64'h10234c18_681ce13d,
        64'hbb6ff0ef_c402c252,
        64'h01311023_8522858a,
        64'h46014000_0cb78002,
        64'h0c3700ff_8bb74b05,
        64'h02900a93_4a550370,
        64'h09933e90_0913cc1c,
        64'h800207b7_00f71563,
        64'h0aa00793_00c14703,
        64'he911bf8f_f0efc23e,
        64'hc43a8522_858a4601,
        64'h47d50aa0_0713e399,
        64'h1aa00713_8ff94bdc,
        64'h00ff8737_681c00f1,
        64'h102347a1_000505a3,
        64'h45d000ef_8522f149,
        64'h84aacf2f_f0ef8522,
        64'hf1dff0ef_85224581,
        64'h4601b72f_f0ef8522,
        64'hd85c4785_08f42223,
        64'h1a042823_18042e23,
        64'h08842783_f94584aa,
        64'h97826b9c_679c8522,
        64'h681c4210_10ef7d00,
        64'h0513ba2f_f0ef8522,
        64'h02042c23_02f40823,
        64'h47851af4_2c23478d,
        64'hf93ff0ef_f3e54481,
        64'h541c8082_61097ca2,
        64'h7c427be2_6b066aa6,
        64'h6a4669e6_74a67906,
        64'h85267446_70e6f850,
        64'h0493bacf_f0effce5,
        64'h05130000_55170204,
        64'h2423eb8d_6b9c679c,
        64'h681cc509_f11ff0ef,
        64'h842ac17c_8fd9f466,
        64'hf862fc5e_e0dae4d6,
        64'he8d2ecce_f0caf4a6,
        64'hfc86f8a2_070d4b9c,
        64'h71191000_0737691c,
        64'h80828082_c2cff06f,
        64'h02c50823_dd0c0007,
        64'h059b00e7_f46385be,
        64'h27814f18_87ae00f5,
        64'hf3634f5c_6918ee09,
        64'hb7cdc402_fef414e3,
        64'h47858082_61217902,
        64'h74a27442_70e2d34f,
        64'hf0ef8526_858a4601,
        64'hc43e4789_00f41f63,
        64'h4791c24a_00f11023,
        64'h4799ed19_d52ff0ef,
        64'hc43ec24a_8526858a,
        64'h46010107_979b4955,
        64'h842e07c4_d78300f1,
        64'h10230370_079304f5,
        64'h92635529_478500f5,
        64'h866384aa_4791f04a,
        64'hf822fc06_f4267139,
        64'h80820141_640260a2,
        64'h45058302_014160a2,
        64'h64028522_00030763,
        64'h0187b303_679c681c,
        64'h00055e63_810ff0ef,
        64'h842ae406_e0221141,
        64'hb32ddd79_842a945f,
        64'hf0ef854a_45850a70,
        64'h061386ce_bb3d842a,
        64'h957ff0ef_854a4585,
        64'h09b00613_46850137,
        64'h9b630a7a_4783d4fb,
        64'h0de34785_ed19975f,
        64'hf0ef854a_458509c0,
        64'h061386de_fdb498e3,
        64'h0c110ff4_f493248d,
        64'hffac90e3_0ffafa93,
        64'h2ca12a85_e13999df,
        64'hf0ef854a_0ff6f693,
        64'h0196d6bb_45858656,
        64'h000c2683_4c818aa6,
        64'h09b00d93_4d61ffa4,
        64'h92e32ca1_0ff4f493,
        64'h2485e935_9cbff0ef,
        64'h854a4585_86260ff6,
        64'hf693019a_d6bb08f0,
        64'h0d134c81_ffb492e3,
        64'h2d210ff4_f4932485,
        64'hed499f1f_f0ef854a,
        64'h45858626_0ff6f693,
        64'h01acd6bb_08c00d93,
        64'h4d010880_049308f9,
        64'h2a2300a7_979b0e0a,
        64'h47830afa_07a34785,
        64'he569a21f_f0ef854a,
        64'h45850af0_06134685,
        64'he3958b85_0afa4783,
        64'he20b02e3_b51d547d,
        64'hdbaff0ef_1bc50513,
        64'h00005517_cb898b85,
        64'h09ba4783_bfd100f9,
        64'hf9b3fff7_c793b591,
        64'h370020ef_18c50513,
        64'h00005517_ef898b85,
        64'h0a6a4783_02d98263,
        64'hfcc592e3_872e0ff9,
        64'hf99300f9_e9b3c70d,
        64'h4189d99b_4187d79b,
        64'h8b050189_999b0187,
        64'h979b0027_571b00b5,
        64'h17bb0208_04630018,
        64'h78130017_581b4b18,
        64'h9726070e_0017059b,
        64'h46114505_47010016,
        64'he993c399_0fe6f993,
        64'h8b89c719_89b60017,
        64'hf7130a7a_46830084,
        64'hc783b5c1_e56ff0ef,
        64'h1d850513_00005517,
        64'h85ce0136_7a63963e,
        64'h09da4783_9e3d0087,
        64'h979b0106_161b09ea,
        64'h478309fa_4603ee05,
        64'h19e3842a_f94ff0ef,
        64'h854a85d2_fe0a7a13,
        64'h02f10a13_f00600e3,
        64'h1e850513_00005517,
        64'h8a09000b_8963fbc5,
        64'h96e387ae_05110821,
        64'h013309bb_0ffbfb93,
        64'h00dbebb3_00be96bb,
        64'hcb898b85_0107c783,
        64'h97a6078e_02088063,
        64'h00652023_02e8d33b,
        64'hb7f14b81_4a814c81,
        64'hb7c1ee4f_f0ef2065,
        64'h05130000_55170003,
        64'h0d6302e8_f33b0017,
        64'h859b0008_28834e11,
        64'h4e854781_89d68562,
        64'h00c48813_8c0a009c,
        64'h9c9be399_4b8502ea,
        64'hdabb02c9_2783bf41,
        64'h5429f24f_f0ef20e5,
        64'h05130000_5517cb89,
        64'h02ecf7bb_0005ac83,
        64'he79102ea_f7bb060a,
        64'h81630045_aa83db45,
        64'h20850513_00005517,
        64'h09892703_80822a01,
        64'h01132381_3d832401,
        64'h3d032481_3c832501,
        64'h3c032581_3b832601,
        64'h3b032681_3a832701,
        64'h3a032781_39832801,
        64'h39032881_34832901,
        64'h34032981_30838522,
        64'hf8400413_f96ff0ef,
        64'h23050513_00005517,
        64'he7b90016_779307e9,
        64'h460300e7_eb6320e5,
        64'h05130000_551784ae,
        64'h8b32892a_bfe78793,
        64'h3ffc07b7_9f3dbff7,
        64'h879bbffc_07b74d18,
        64'h0ac7e963_478923b1,
        64'h3c2325a1_30232591,
        64'h34232581_38232571,
        64'h3c232761_30232751,
        64'h34232741_38232731,
        64'h3c232921_30232891,
        64'h34232881_38232811,
        64'h3c23d601_01138082,
        64'h614569a2_694264e2,
        64'h740270a2_85220135,
        64'h05a315e0_10ef8526,
        64'h842a875f_f0ef8526,
        64'h85ca0009_1c6300f5,
        64'h1e63842a_57b5c519,
        64'hcc7ff0ef_84aa4585,
        64'h0b300613_8edd892e,
        64'h9be10079_f6930ff5,
        64'hf9930815_4783f022,
        64'hf406e44e_e84aec26,
        64'h7179b74d_84aab75d,
        64'hdf400493_f7d50b94,
        64'h4783e519_98dff0ef,
        64'h854a85a2_980101f1,
        64'h0413f1e9_258199f5,
        64'hffe4059b_f57184aa,
        64'hd1fff0ef_892a4585,
        64'h0b900613_842e4685,
        64'hfef760e3_4705ffc5,
        64'h879b8082_24010113,
        64'h22813483_22013903,
        64'h85262301_34032381,
        64'h308354a9_c5854681,
        64'h02b7e163_02f58863,
        64'h47892321_30232291,
        64'h34232281_38232211,
        64'h3c23dc01_0113bf45,
        64'h5929bf55_5951bf65,
        64'h1a04b023_5c8020ef,
        64'hd1691a04_b503892a,
        64'hbf4d08f4_aa2302f7,
        64'h07bb2785_27058bfd,
        64'h8b7d0057_d79b00a7,
        64'hd71b50fc_80822501,
        64'h01132281_39832301,
        64'h39032381_3483854a,
        64'h24013403_24813083,
        64'h08f48023_0a744783,
        64'h08d4ac23_02f686bb,
        64'h00a6969b_0dd44783,
        64'hf8dc07a6_0d442783,
        64'h00098663_c79954dc,
        64'h08f4aa23_00a6979b,
        64'hc7b98b85_0e044683,
        64'h0af44783_0af407a3,
        64'h4785ed35_e0bff0ef,
        64'h85264585_0af00613,
        64'h4685ce81_e3918bfd,
        64'h09c44783_c7898b85,
        64'h0a044783_f4fc07a6,
        64'hc319f4fc_54d89fb9,
        64'h08844703_9fb90087,
        64'h171b0894_47039fb9,
        64'h0107171b_0187979b,
        64'h08a44703_08b44783,
        64'hf8fc07ce_02e787b3,
        64'h0dd44783_02f70733,
        64'h0e044703_97ba08c4,
        64'h47039fb9_0087171b,
        64'h0107979b_468508d4,
        64'h470308e4_47830409,
        64'h8f63fca7_14e30621,
        64'h070de21c_07ce02b7,
        64'h87b30dd4_478302f5,
        64'h85b30e04_45830009,
        64'h8c634685_c39197ae,
        64'hffe74583_9fad0105,
        64'h959b0087_979b0007,
        64'h4583fff7_4783e0fc,
        64'h07c64681_09d40513,
        64'h0a844783_fcdc07c6,
        64'h0c848613_09140713,
        64'h0e244783_06f48fa3,
        64'h09c44783_c7898b89,
        64'h0a044783_00098a63,
        64'h08f480a3_0b344783,
        64'hc7890e24_4783e781,
        64'h0019f993_8b8506f4,
        64'h8f2309b4_49830a04,
        64'h4783f8dc_00d77363,
        64'h0147d693_07a68007,
        64'h07136705_0d442783,
        64'h00e7fd63_cc981ff7,
        64'h87934004_07b753b8,
        64'h97ba078a_1f470713,
        64'h00004717_1cf76b63,
        64'h47210c04_47831230,
        64'h10ef85a2_20000613,
        64'h1e050363_1a04b503,
        64'h1aa4b023_766020ef,
        64'h20000513_e7991a04,
        64'hb7831e05_1863892a,
        64'hc09ff0ef_84aa85a2,
        64'h980101f1_04131ce7,
        64'hf5634901_3ffc0737,
        64'h23313423_22913c23,
        64'h24813023_24113423,
        64'h9fb92321_3823bffc,
        64'h07b7db01_01134d18,
        64'hbfcdfc79_347d8082,
        64'h612174a2_744270e2,
        64'hd91ff0ef_85263e80,
        64'h0593e919_c53ff0ef,
        64'h8526858a_4601440d,
        64'hc43684aa_fc06f426,
        64'hf8228ed1_0106161b,
        64'h8edd0300_07b70086,
        64'h969bc23e_47f500f1,
        64'h10234799_71398082,
        64'h61216aa2_6a4269e2,
        64'h74a27902_85267442,
        64'h70e2fc09_99e39aa2,
        64'h02878433_9a224089,
        64'h89b308c9_6783fc85,
        64'h1ae3f01f_f0ef854a,
        64'h85d68652_86a2844e,
        64'h0089f363_0207e403,
        64'h01093783_89a6f96d,
        64'hecdff0ef_854a08c9,
        64'h2583a089_4481bd9f,
        64'hf0ef60a5_05130000,
        64'h551700b6_7a630144,
        64'h85b36810_00054d63,
        64'h8c9fa0ef_852200b4,
        64'h4583c11d_892a4820,
        64'h10ef8ab6_84b28a2e,
        64'h4148842a_ce05e456,
        64'he852ec4e_f04af426,
        64'hf822fc06_7139b7c5,
        64'h4401b7d5_0004841b,
        64'hb74d02f6_063bbf61,
        64'h47c58082_61256906,
        64'h64a66446_60e68522,
        64'hc43ff0ef_65450513,
        64'h00005517_c11dd55f,
        64'hf0efd23e_d402854a,
        64'h100c47f5_460102f1,
        64'h102347b1_0497f063,
        64'h4785e529_842ad75f,
        64'hf0efc83e_ca26d23a,
        64'h854a100c_47850030,
        64'hcc3ee42e_4755d432,
        64'hcf3108c9_27832601,
        64'h02f11023_02c92703,
        64'h47c906d7_f66384b6,
        64'h892a4785_e8a2ec86,
        64'he0cae4a6_711d8082,
        64'h4501bfd5_45018082,
        64'h612174a2_744270e2,
        64'hf8ed34fd_c901dcdf,
        64'hf0ef8522_858a4601,
        64'h4495cb91_8b891b84,
        64'h2783c11d_de3ff0ef,
        64'hc23e842a_f426fc06,
        64'hf822858a_460147d5,
        64'hc42e00f1_102347c1,
        64'h7139e7a9_19c52783,
        64'hbf7df920_0513d09f,
        64'hf0ef6fa5_05130000,
        64'h5517fc80_49e34501,
        64'hb7555d80_20ef3e80,
        64'h051300f0_57630014,
        64'h079b347d_fe04c6e3,
        64'h34fd8082_61257aa2,
        64'h7a4279e2_690664a6,
        64'h644660e6_fba00513,
        64'hd4bff0ef_72450513,
        64'h00005517_c78d0125,
        64'hf7b30547_93630135,
        64'hf7b3c789_1005f793,
        64'h45b2ed0d_e73ff0ef,
        64'h8556858a_4601e00a,
        64'h0a13e009_89930809,
        64'h09134495_c43e842e,
        64'h8aaaec86_f456e4a6,
        64'he8a26a05_6989fdf9,
        64'h49370107_979bf852,
        64'hfc4ee0ca_07c55783,
        64'hc23e47d5_00f11023,
        64'h47b5711d_80826145,
        64'h740270a2_c43c47b2,
        64'he119ec9f_f0ef8522,
        64'h858a4601_c43e8fd9,
        64'h8f554000_06b78f75,
        64'h600006b7_8ff58ff9,
        64'hf8078793_4ad40080,
        64'h07b74538_6914c195,
        64'h842ac402_c23ef406,
        64'hf0224785_00f11023,
        64'h47857179_80826145,
        64'h740270a2_85226cc0,
        64'h20ef7d00_0513e509,
        64'h842af21f_f0efc202,
        64'hc4020001_1023858a,
        64'h46018522_6ea020ef,
        64'hf4063e80_0513842a,
        64'hf0227179_b761fb60,
        64'h0513d551_56f010ef,
        64'h0d448513_0d440593,
        64'h461100f7_1a630e04,
        64'h47830e04_c70302f7,
        64'h10630c04_47830c04,
        64'hc70302f7_16630dd4,
        64'h47830dd4_c70302f7,
        64'h1c630a04_47830a04,
        64'hc703f579_f95ff0ef,
        64'h1a053483_22113c23,
        64'h22913423_85a29801,
        64'h01f10413_22813823,
        64'hdc010113_80822401,
        64'h01132281_34832301,
        64'h34032381_30834501,
        64'h80824501_00e6fe63,
        64'h40040737_4d148082,
        64'h616160a6_fd3ff0ef,
        64'hcc3ed402_e486100c,
        64'h20000793_0030e83e,
        64'he42e0785_17824785,
        64'hd23e47d5_02f11023,
        64'h47a1715d_83020007,
        64'hb303679c_691c8082,
        64'h8c850513_00006517,
        64'h80826108_953e8175,
        64'h64878793_00004797,
        64'h150200a7_eb6347ad,
        64'h8082557d_80820141,
        64'h640260a2_45018302,
        64'h014160a2_64028522,
        64'h00030763_0207b303,
        64'h679c681c_00055e63,
        64'hff5ff0ef_842ae406,
        64'he0221141_8082557d,
        64'h8082557d_b7e9659c,
        64'h95aa058e_05e135f1,
        64'hbfd9617c_bfe97d5c,
        64'h80826105_4501e91c,
        64'h64a26442_60e202f4,
        64'h57b39381_02049793,
        64'h0c5010ef_7540f55c,
        64'h08c52483_795c8782,
        64'h97bae426_e822ec06,
        64'h1101439c_97ba83f9,
        64'h6c070713_00004717,
        64'h02059793_04b7ee63,
        64'h479d8082_45018302,
        64'h00030363_0087b303,
        64'h679c691c_80826135,
        64'h645260f2_85221290,
        64'h20ef0808_842ae3ff,
        64'hf0efe436_eec6eac2,
        64'he6bee2ba_ea22ee06,
        64'h08081000_05931234,
        64'h862afe36_fa32f62e,
        64'h710d8082_616160e2,
        64'he69ff0ef_e436e4c6,
        64'he0c2fc3e_f83aec06,
        64'h10000593_1014862e,
        64'hf436f032_715d8082,
        64'h616160e2_e8dff0ef,
        64'he436e4c6_e0c2fc3e,
        64'hf83aec06_1034f436,
        64'h715db7f1_85220201,
        64'h03930005_059b4db0,
        64'h10ef8522_01247433,
        64'h60000084_0b13b5fd,
        64'h845ad93f_f0ef0084,
        64'h0b130201_03930004,
        64'h4503a809_ddbff0ef,
        64'h00280201_03930005,
        64'h059be37f_f0ef4008,
        64'h45a94601_0016b693,
        64'h00380084_0b13f8b5,
        64'h0693a811_45c10016,
        64'h36134685_00380084,
        64'h0b13fa85_0613f6e5,
        64'h10e30780_071302e5,
        64'h00630750_0713a00d,
        64'h46014685_00380084,
        64'h0b13f6e5_1ee30700,
        64'h071300a7_6c6306e5,
        64'h0e630730_0713b74d,
        64'h048d0024_c5038082,
        64'h61090007_051b6b06,
        64'h6aa66a46_69e67906,
        64'h74a67446_70e6f55d,
        64'h08f50963_06300793,
        64'h04d50f63_05800693,
        64'h02a6eb63_06d50f63,
        64'h06400693_04890014,
        64'hc5034781_00f6f363,
        64'h46a50ff7_f793fd07,
        64'h879bcb9d_0004c783,
        64'h03551063_47810489,
        64'h05450f63_0014c503,
        64'hbfe1e7bf_f0ef0201,
        64'h03930485_01350863,
        64'h04d7ff63_93811782,
        64'h76820017_079bc52d,
        64'h8f1d0004_c50377a2,
        64'h77420209_59130300,
        64'h0a9306c0_0a130250,
        64'h0993f82a_f02ef42a,
        64'hfc3e8436_84b2e0da,
        64'hfc86e4d6_e8d2ecce,
        64'hf4a6f8a2_597d011c,
        64'hf0ca7119_b7f10685,
        64'h01178023_00668023,
        64'h26050006_c8830007,
        64'hc30397ba_93811782,
        64'h40c807bb_b7d92585,
        64'hfea68fa3_0685bf5d,
        64'h00a8053b_808200b6,
        64'h1b63fff5_081b86ba,
        64'h25810006_80230015,
        64'h559b40e6_853b0685,
        64'h00f68023_02d00793,
        64'h00088763_02f5e963,
        64'h03000513_40e685bb,
        64'hfe718532_fea68fa3,
        64'h06850ff5_751302b6,
        64'h563b0305_051b046e,
        64'h67630ff3_751302b6,
        64'h733b0005_061b3859,
        64'h86ba4e25_0ff6f813,
        64'h04100693_c2190610,
        64'h06934885_40a0053b,
        64'he6810005_56634881,
        64'hbfe900d7_00230785,
        64'h0007c683_00d3b823,
        64'h00170693_8082852e,
        64'h00070023_00b6e663,
        64'h0103b703_40a786bb,
        64'h87aa9d9d_fff7059b,
        64'h00c6f563_8e9dfff7,
        64'h06930003_b7038f99,
        64'h92010205_96130103,
        64'hb7830083_b7038082,
        64'h45018082_00078023,
        64'h45050103_b78300a7,
        64'h002300f3_b8230017,
        64'h079300d7_fe639381,
        64'h17822785_40f707b3,
        64'h0003b683_0083b783,
        64'h0103b703_80826145,
        64'h45016a02_69a26942,
        64'h64e27402_70a22e80,
        64'h00ef27a5_05130000,
        64'h6517fd24_9fe30405,
        64'h2fa000ef_819100f5,
        64'hf6132485_854e0004,
        64'h458330c0_00ef8552,
        64'h85a6e789_01f4f793,
        64'h20000913_ccc98993,
        64'h00006997_ccca0a13,
        64'h00006a17_4481ed5f,
        64'hf0ef8426_45818526,
        64'h33a000ef_ccc50513,
        64'h00006517_fa460613,
        64'h00006617_e789c466,
        64'h06130000_6617584c,
        64'h19c42783_db9fb0ef,
        64'h2f058593_00006597,
        64'h74481020_30efcee5,
        64'h05130000_65173780,
        64'h00efce25_05130000,
        64'h6517c6a5_85930000,
        64'h6597c789_c7c58593,
        64'h00006597_545c3980,
        64'h00efcf25_05130000,
        64'h65175c0c_3a6000ef,
        64'h26010ff6_f6930ff7,
        64'hf7930ff7_77130187,
        64'hd61b0107_d69b0087,
        64'hd71bd025_05130000,
        64'h651706c4_4583583c,
        64'h3d2000ef_91c115c2,
        64'h0085d59b_d0c50513,
        64'h00006517_546c3e80,
        64'h00efd025_05130000,
        64'h651706f4_45833f80,
        64'h00ef638c_d0450513,
        64'h00006517_681c2060,
        64'h10ef842a_491010ef,
        64'h450144b0_10ef0001,
        64'hb5031b20_30efd1e5,
        64'h05130000_651784aa,
        64'h0aa030ef_e052e44e,
        64'he84aec26_f022f406,
        64'h20000513_71797940,
        64'h006f6105_468560e2,
        64'h66226442_85a24d30,
        64'h10efe42e_ec064501,
        64'h842ae822_11018082,
        64'h01416402_60a2557d,
        64'he3914505_703c1700,
        64'h30efcba5_05130000,
        64'h6517caa5_85930000,
        64'h659734c0_0613b666,
        64'h86930000_569702f4,
        64'h02634200_07b7e406,
        64'h6380e022_1141711c,
        64'h80822501_6108953e,
        64'h050e4200_07b7f73f,
        64'hf06f4200_05374581,
        64'h46098082_bff9557d,
        64'h18c030ef_8522b7e5,
        64'hc45c4785_d4fd4501,
        64'h88858082_614569a2,
        64'h694264e2_740270a2,
        64'h4501c45c_4789cb99,
        64'h0024f793_f4040124,
        64'h2423e01c_420007b7,
        64'h02098b63_4fe000ef,
        64'hdc850513_00006517,
        64'h862285aa_89aa7850,
        64'h10efbca5_05130000,
        64'h551785a2_cc1d5551,
        64'h842a1a40_30ef892e,
        64'h84b2e44e_f406e84a,
        64'hec26f022_04800513,
        64'h717908b0_41635535,
        64'hb7dd87ca_0ca139a0,
        64'h20efe43e_002c4621,
        64'h8566639c_00878913,
        64'hfa978de3_94be0009,
        64'h3c830109_648397a6,
        64'h67a1bf41_b1dff0ef,
        64'h8522b771_00f92623,
        64'h000cb783_dbd98b85,
        64'hbd956410_20ef4505,
        64'hd80c8ee3_c47ff0ef,
        64'h8522484c_c85c9bf5,
        64'h4c85485c_b4dff0ef,
        64'h8522ef8d_8b850089,
        64'h27830009_09630404,
        64'h30232b40_30ef8556,
        64'h85d20ca0_0613c5e6,
        64'h86930000_56970174,
        64'h8c630404_39036004,
        64'hcc9d4c85_8889c85c,
        64'h9bf9485c_c85c0027,
        64'he793485c_cbb5603c,
        64'hfeb690e3_0791872a,
        64'h2685c398_8f518361,
        64'hff873703_01068763,
        64'hc3900086_161bff87,
        64'h05136310_4591480d,
        64'h468100c9_0793018c,
        64'h871308e6_9f630037,
        64'hf693470d_02043c23,
        64'h00492783_cba97c1c,
        64'h332030ef_855685d2,
        64'h09c00613_cc468693,
        64'h00005697_017c8c63,
        64'h03843903_00043c83,
        64'hcfb50014_f7936580,
        64'h00efefa5_05130000,
        64'h651785ca_d1fff0ef,
        64'h85ca0049_6913ff39,
        64'h79138522_01442903,
        64'hc3950084_f7936800,
        64'h00efefa5_05130000,
        64'h651785ca_d47ff0ef,
        64'h85ca0089_6913ff39,
        64'h79138522_01442903,
        64'hc3950044_f793b27f,
        64'hf0ef8522_4581b6ff,
        64'hf0ef8522_4581cc5c,
        64'hf9200793_c7817c1c,
        64'h00f76f63_0c893783,
        64'h02093703_12048e63,
        64'h24818cfd_4c81485c,
        64'h07093483_3de030ef,
        64'h855685d2_0f200613,
        64'h86e20179_09630004,
        64'h3903b711_6f6000ef,
        64'hf5850513_00006517,
        64'hd5858593_00005597,
        64'h000b1d63_3b7d4200,
        64'h0bb78b4e_bd6100c4,
        64'he493bd85_41e030ef,
        64'hf6850513_00006517,
        64'hf5858593_00006597,
        64'h14900613_d7468693,
        64'h00005697_b7654701,
        64'h47812585_e31c9746,
        64'h93818375_17821702,
        64'h00be873b_8fd98fe9,
        64'h01076733_0087d79b,
        64'h01c87833_0087981b,
        64'h01076733_0187971b,
        64'h0187d81b_f2e50067,
        64'h036316fd_06052781,
        64'h0107e7b3_01e8183b,
        64'h07050037_1f1b0006,
        64'h4803ec06_89e36e89,
        64'hf0050513_00ff0e37,
        64'h43114701_47814581,
        64'h63900107_e6836541,
        64'h00043883_603cee07,
        64'h9be38b85_449cdf3f,
        64'hf0ef8522_488cdb7f,
        64'hf0efe024_852244cc,
        64'h80826165_45016ce2,
        64'h7c027ba2_7b427ae2,
        64'h6a0669a6_694664e6,
        64'h740670a6_efe9485c,
        64'h038a8a93_00006a97,
        64'h68198993_eb7ff0ef,
        64'h25810015_e5930098,
        64'h99b78522_0d89b583,
        64'hcd1ff0ef_85224585,
        64'he93ff0ef_85222405,
        64'h8593000f_45b7d27f,
        64'hf0ef8522_45814605,
        64'h46854705_cf5ff0ef,
        64'h85224581_cbdff0ef,
        64'h852285a6_c81ff0ef,
        64'h078a0a13_00006a17,
        64'h85220009_5583c4ff,
        64'hf0efed2c_0c130000,
        64'h5c178522_00892583,
        64'hbe1ff0ef_85224581,
        64'hd71ff0ef_85224581,
        64'h46054681_47050144,
        64'he4931607_86638b85,
        64'h008a2783_000a0963,
        64'h8cdd0324_3c234c1c,
        64'h4485e391_448d8b89,
        64'hc7090017_f7134481,
        64'h00492783_16f99a63,
        64'h04043a03_420007b7,
        64'h00043983_bf5ff0ef,
        64'h45856008_0e049c63,
        64'h6ca020ef_00c90513,
        64'h45814611_d01ce030,
        64'h84b2892e_0005d783,
        64'h020408a3_ec66f062,
        64'hf45ef85a_fc56e0d2,
        64'he4cef486_e8caeca6,
        64'h7100f0a2_71598082,
        64'h61056902_64a26442,
        64'h60e2c844_04993c23,
        64'h612030ef_15c50513,
        64'h00006517_14c58593,
        64'h00006597_07600613,
        64'hf5868693_00005697,
        64'h02f90263_84ae842a,
        64'h420007b7_ec06e426,
        64'he8220005_3903e04a,
        64'h11018082_610564a2,
        64'h644260e2_e4246580,
        64'h30ef1a25_05130000,
        64'h65171925_85930000,
        64'h659706f0_0613f8e6,
        64'h86930000_569702f4,
        64'h026384ae_420007b7,
        64'hec06e426_6100e822,
        64'h11018082_610564a2,
        64'h644260e2_e0a08c7d,
        64'h17fd6785_69e030ef,
        64'h1e850513_00006517,
        64'h1d858593_00006597,
        64'h06800613_fc468693,
        64'h00005697_02f48263,
        64'h842e4200_07b7ec06,
        64'he8226104_e4261101,
        64'h80826105_64a26442,
        64'h60e2fc80_90411442,
        64'h6e2030ef_22c50513,
        64'h00006517_21c58593,
        64'h00006597_06100613,
        64'hff868693_00005697,
        64'h02f48263_842e4200,
        64'h07b7ec06_e8226104,
        64'he4261101_d4dff06f,
        64'h01414581_60a26402,
        64'h6008f23f_f0ef4605,
        64'h46854705_45818522,
        64'hef1ff0ef_45818522,
        64'hf39ff0ef_842a4581,
        64'h04053023_02053c23,
        64'h46054681_4705e022,
        64'he4061141_80820141,
        64'h45016402_60a2d97f,
        64'hf0ef4581_6008f67f,
        64'hf0ef4581_46054685,
        64'h47058522_f35ff0ef,
        64'h45818522_f7dff0ef,
        64'he4064581_85224605,
        64'h46814705_7100e022,
        64'h11418082_612169e2,
        64'h790274a2_02b9b823,
        64'h8dc57442_70e288a1,
        64'h0125e5b3_0034949b,
        64'h8dd90049_79130029,
        64'h191b8b05_89890014,
        64'h159b6722_7c6030ef,
        64'he43a3125_05130000,
        64'h65173025_85930000,
        64'h659705a0_06130ce6,
        64'h86930000_569702f9,
        64'h84638436_893284ae,
        64'h420007b7_fc06f04a,
        64'hf426f822_00053983,
        64'hec4e7139_80826105,
        64'h64a26442_60e2f404,
        64'h013030ef_35c50513,
        64'h00006517_34c58593,
        64'h00006597_05300613,
        64'h10868693_00005697,
        64'h02f40263_84ae4200,
        64'h07b7ec06_e4266100,
        64'he8221101_80826105,
        64'h64a26442_60e2f004,
        64'h053030ef_39c50513,
        64'h00006517_38c58593,
        64'h00006597_04c00613,
        64'h13868693_00005697,
        64'h02f40263_84ae4200,
        64'h07b7ec06_e4266100,
        64'he8221101_80826105,
        64'h64a26442_60e2ec80,
        64'h90011402_097030ef,
        64'h3e050513_00006517,
        64'h3d058593_00006597,
        64'h04500613_04c68693,
        64'h00007697_02f48263,
        64'h842e4200_07b7ec06,
        64'he8226104_e4261101,
        64'h80826105_64a26442,
        64'h60e2e880_90011402,
        64'h0db030ef_42450513,
        64'h00006517_41458593,
        64'h00006597_03e00613,
        64'h09868693_00007697,
        64'h02f48263_842e4200,
        64'h07b7ec06_e8226104,
        64'he4261101_80826105,
        64'h64a26442_60e2e404,
        64'h11b030ef_46450513,
        64'h00006517_45458593,
        64'h00006597_03600613,
        64'h1f068693_00005697,
        64'h02f40263_84ae4200,
        64'h07b7ec06_e4266100,
        64'he8221101_80826105,
        64'h64a26442_60e2e004,
        64'h15b030ef_4a450513,
        64'h00006517_49458593,
        64'h00006597_02f00613,
        64'h22068693_00005697,
        64'h02f40263_84ae4200,
        64'h07b7ec06_e4266100,
        64'he8221101_80826105,
        64'h64a26442_60e2fc24,
        64'h19b030ef_4e450513,
        64'h00006517_4d458593,
        64'h00006597_08800613,
        64'h24868693_00005697,
        64'h02f50263_84ae842a,
        64'h420007b7_ec06e426,
        64'he8221101_8082556d,
        64'hbfe50007_ac238082,
        64'h4501cf98_02000713,
        64'h00d71763_469100d7,
        64'h0d63711c_46a15958,
        64'h80826149_640a60aa,
        64'hf83ff0ef_0808f01f,
        64'hf0ef0808_e85ff0ef,
        64'h080885a2_6622f71f,
        64'hf0efe42e_e5060808,
        64'h842ae122_71758082,
        64'h610531a5_05130000,
        64'h751760e2_fca71de3,
        64'hfef68fa3_fec68f23,
        64'h0007c783_97ae0006,
        64'h46038bbd_962e0047,
        64'hd6130705_06890007,
        64'hc78300e1_07b34541,
        64'h57058593_00006597,
        64'h35868693_00007697,
        64'h47013bf0_20efec06,
        64'h850a4641_05050593,
        64'h11018082_e13cb6c7,
        64'h87930000_0797ed3c,
        64'h639c13a7_87930000,
        64'h7797e93c_04053423,
        64'h639c1427_87930000,
        64'h77978082_614569a2,
        64'h694264e2_740270a2,
        64'hfd24fde3_45019782,
        64'h8522603c_fc1c078e,
        64'h643c0124_f5633c90,
        64'h20ef9522_45819201,
        64'h16020006_091b40a9,
        64'h863b449d_04000993,
        64'h00e78023_97a2f800,
        64'h07130017_8513e84a,
        64'hf406e44e_ec26842a,
        64'h03f7f793_f0227179,
        64'h653c8082_61616ba2,
        64'h6b426ae2_7a0279a2,
        64'h794274e2_640660a6,
        64'hb7c99782_44018526,
        64'h60bc0174_176399d6,
        64'h41590933_481020ef,
        64'h0144043b_86560084,
        64'h853385ce_020ada93,
        64'h020a1a93_00090a1b,
        64'h00f97463_93811782,
        64'h00078a1b_408b07bb,
        64'h04000b93_04000b13,
        64'he53c8932_89ae84aa,
        64'h97b203f7_f413ec56,
        64'hf052e486_e45ee85a,
        64'hf44ef84a_fc26e0a2,
        64'h715d653c_80826105,
        64'h692264c2_cd70cd34,
        64'hc97c0505_282300c8,
        64'h863b00d3_06bb00fe,
        64'h07bb010e_883b6462,
        64'hf3ef9de3_00e587bb,
        64'h0005869b_0003861b,
        64'h0f118f5d_0157171b,
        64'h00b7579b_9f3d0077,
        64'h47339fa1_8f4dfff7,
        64'h47130007_081b00b3,
        64'h85bb4080_9fa18dd5,
        64'h0115d59b_94aa00f5,
        64'h969b048a_9db5ffc2,
        64'ha4038db9_02c10075,
        64'he5b3fff7_c593023f,
        64'h44839ead_00c703bb,
        64'h00c3e633_400c9ead,
        64'h0166561b_00a6139b,
        64'h0082a583_9e2d8e3d,
        64'h8e59fff6_c6139db1,
        64'h00f8073b_01076833,
        64'h01a8581b_0003a583,
        64'h9e2d0068_171b0107,
        64'h083b0042_a5839f2d,
        64'h942a040a_418c95aa,
        64'h058a93aa_038a020f,
        64'h45839f2d_022f4403,
        64'h021f4383_0002a703,
        64'h00d745b3_8f5dfff6,
        64'h471349a2_82930000,
        64'h5297f5f5_92e300e4,
        64'h07bb0004_069b0002,
        64'h861b0f91_8f5d0177,
        64'h171b0097_579b9f3d,
        64'h8f219fa5_00574733,
        64'h0007081b_00d2843b,
        64'h8ec10009_24830106,
        64'hd69b9fa5_0106941b,
        64'h992a9ea1_090a0056,
        64'hc6b300e7_c6b3ffc3,
        64'ha4839c35_00c702bb,
        64'h03c100c2_e6330156,
        64'h561b013f_c90300b6,
        64'h129b4080_00c2863b,
        64'h9ea194aa_00e2c2b3,
        64'h048a00f8_073b0083,
        64'ha4039e21_01076833,
        64'h01c8581b_0048171b,
        64'h012fc483_0107083b,
        64'h40809e21_94aa048a,
        64'h0043a403_9f21011f,
        64'hc4839f25_400000c2,
        64'hc4b3942a_040a00d7,
        64'hc2b30003_a703010f,
        64'hc4035223_83930000,
        64'h53978ffa_5acf0f13,
        64'h00005f17_f25599e3,
        64'h00e407bb_0004069b,
        64'h0003861b_000f081b,
        64'h8f5d0147_171b00c7,
        64'h579b9f3d_00774733,
        64'h01e77733_0083c733,
        64'h9fb900d3_843b8ec1,
        64'h40980126_d69b9fb9,
        64'h00e6941b_94aa048a,
        64'hffcfa703_9eb90fc1,
        64'h01e6c6b3_fff5c483,
        64'h8efd007f_46b30591,
        64'h9f3500cf_03bb00c3,
        64'he6334018_9eb90176,
        64'h561b0096_139b008f,
        64'ha7039e39_8e3d8e75,
        64'h01e7c633_9f3100f8,
        64'h0f3b010f_68330003,
        64'ha70301b8_581b9e39,
        64'h00581f1b_010f083b,
        64'h004fa703_00ef0f3b,
        64'h942a040a_4318972a,
        64'h070a93aa_038a0005,
        64'hc70300ef_0f3b0025,
        64'hc4030015_c383000f,
        64'haf0301e6_c73300cf,
        64'h7f3300d7_cf336962,
        64'h82930000_52975cef,
        64'h8f930000_5f976965,
        64'h85930000_5597f45f,
        64'h17e300e3_87bb0003,
        64'h869b0005_881b0f41,
        64'h8f5d0167_171b00a7,
        64'h579b9f3d_8f2d9fa1,
        64'h00777733_8f2d0007,
        64'h061b00d7_03bbffcf,
        64'ha4039fa1_00d3e6b3,
        64'h0116969b_00f6d39b,
        64'h007686bb_8ebd00cf,
        64'h24038ef9_00b7c6b3,
        64'h00d383bb_00c5873b,
        64'h008383bb_8e590146,
        64'h561b00c6_171b9e39,
        64'h008f2383_8e358e6d,
        64'h00f6c633_9f3100f8,
        64'h05bb0077_073b0105,
        64'he8330198_581b0078,
        64'h159b0105_883b004f,
        64'h2703ff4f_a3839db9,
        64'h007585bb_0fc1008f,
        64'ha403000f_2583000f,
        64'ha38300b6_47338dfd,
        64'h00c6c5b3_654f8f93,
        64'h00005f97_887687f2,
        64'h869a8646_04050293,
        64'h8f2ae44a_e826ec22,
        64'h110105c5_28830585,
        64'h23030545_2e030505,
        64'h2e83bf89_eaf71de3,
        64'h0e500793_01814703,
        64'hf8d771e3_0007869b,
        64'h02000613_47299381,
        64'h1782f4c7_e5e30585,
        64'h068500e5_8023f917,
        64'h80e3b751_842abf19,
        64'h00e785a3_47216786,
        64'hae5fd0ef_082c462d,
        64'h6506b07f_d0ef4581,
        64'h02000613_6506f445,
        64'h0005041b_a55fe0ef,
        64'h1028dbd5_01814783,
        64'h02f51b63_4791b7c1,
        64'h0005041b_8fefe0ef,
        64'h00f50223_47857522,
        64'h00f50023_5795a885,
        64'h078500c6_802300fe,
        64'h06b3b7cd_ffe81be3,
        64'h06080563_00054803,
        64'h0505bfcd_f36d8082,
        64'h61256446_60e68522,
        64'h441900ee_f863a821,
        64'h00070f1b_adc50513,
        64'h00007517_93411742,
        64'h370100a3_6c639141,
        64'h1542f9f7_051b2785,
        64'h0006c703_48b107f0,
        64'h0e934365_8e2e4781,
        64'h082cfeb7_06e30007,
        64'h47039736_93010207,
        64'h9713fff6_079bbf45,
        64'h863eb74d_2605a061,
        64'h00e78ca3_00078ba3,
        64'h00078b23_04600713,
        64'h00e78c23_02100713,
        64'h6786bc7f_d0ef082c,
        64'h462dc3dd_65060181,
        64'h4783e179_2501abbf,
        64'he0ef1028_4585e841,
        64'h0005041b_bd6fe0ef,
        64'hda021028_4581ea29,
        64'h02000593_eba10007,
        64'hc78397b6_93810206,
        64'h17934601_00010c23,
        64'h66a2ec55_0005041b,
        64'hee3fd0ef_ec86e8a2,
        64'h1028002c_4605e42a,
        64'h711db7d5_842abf55,
        64'h00048023_00f51563,
        64'h47918082_61256906,
        64'h64a66446_60e68522,
        64'h00a92023_c29fd0ef,
        64'h953e0347_87930270,
        64'h079300e6_84630005,
        64'h46830430_0793470d,
        64'h6562e015_0005041b,
        64'he69fd0ef_510c6562,
        64'h02090a63_fec783e3,
        64'h177d0007_c78397a6,
        64'h93811782_0007869b,
        64'hfff6879b_ce890007,
        64'h00230200_061346ad,
        64'h00b48713_ca1fd0ef,
        64'h8526462d_75c2e93d,
        64'h2501b8ff_e0ef0828,
        64'h4585e559_2501ca8f,
        64'he0efd202_08284581,
        64'hc4b9e051_0005041b,
        64'hf9bfd0ef_ec86e8a2,
        64'h08284601_002c8932,
        64'h84aee42a_e0cae4a6,
        64'h711d8082_61256446,
        64'h60e62501_ad6fe0ef,
        64'h00f50223_478500e7,
        64'h8ca30087_571b00e7,
        64'h8c230044_570300e7,
        64'h8ba30087_571b00e7,
        64'h8b237522_00645703,
        64'hcb856786_eb950207,
        64'hf79300b7_c7834519,
        64'h67a6e129_25019abf,
        64'he0efe4be_1028083c,
        64'h65a2e929_2501810f,
        64'he0efec86_1028002c,
        64'h4605842e_e42ae8a2,
        64'h711dbfcd_47a18082,
        64'h614d853e_64ea740a,
        64'h70aa0005_079bb50f,
        64'he0ef6506_e7910005,
        64'h079be24f_e0ef0088,
        64'h00f70223_06d707a3,
        64'h478506f7_04a30086,
        64'hd69b0106_d69b0087,
        64'hd79b0107_d79b0107,
        64'h979b06f7_04232781,
        64'h0107d79b_06f70723,
        64'h0107969b_57d602f6,
        64'h9d630557_468302e0,
        64'h07936706_efb10005,
        64'h079bfc3f_d0ef8522,
        64'hc5a54789_0005059b,
        64'hcaefe0ef_85220005,
        64'h059bf2df_d0ef85a6,
        64'h00044503_06f70863,
        64'h57d64736_cbbd8bc1,
        64'h00b4c783_00f40223,
        64'h478500f4_85a30207,
        64'he7936406_02814783,
        64'he0dfd0ef_00d48513,
        64'h02a10593_464d648a,
        64'hefc50005_079bdc5f,
        64'he0ef10a8_0ce79363,
        64'h4711cbf9_0005079b,
        64'haadfe0ef_10a86582,
        64'h0c054d63_47adf05f,
        64'hd0ef850a_e49fd0ef,
        64'h10a8008c_02800613,
        64'he55fd0ef_102805ad,
        64'h46550e05_8e634791,
        64'h65e61007_12630207,
        64'h77134799_00b7c703,
        64'h77861007_9a630005,
        64'h079baf7f_e0eff0be,
        64'h083cf4be_008865a2,
        64'h67861207_96630005,
        64'h079b964f_e0efed26,
        64'hf122f506_0088002c,
        64'h4605e02e_e42a7171,
        64'h80826165_64e67406,
        64'h70a62501_c9efe0ef,
        64'h00f50223_47850087,
        64'h05a38c3d_02747413,
        64'h8c658cbd_752200b7,
        64'h4783c30d_6706e39d,
        64'h0207f793_00b7c783,
        64'h451967a6_e9152501,
        64'hb65fe0ef_e4be1028,
        64'h083c65a2_e1312501,
        64'h9cafe0ef_f4861028,
        64'h4605002c_843284ae,
        64'he42aeca6_f0a27159,
        64'hb7c54421_8082614d,
        64'h6d466ce6_7c067ba6,
        64'h7b467ae6_6a0a69aa,
        64'h694a64ea_740a70aa,
        64'h8522f25f_e0ef85ca,
        64'h7522441d_b7498c6a,
        64'h0ffbfb93_f61fd0ef,
        64'h3bfd8552_45812000,
        64'h0613ec09_0005041b,
        64'h8dcfe0ef_01950223,
        64'h03852823_001c0d1b,
        64'h7522a82d_0005041b,
        64'hd5afe0ef_00f50223,
        64'h47850097_8aa30167,
        64'h8a230137_8da30157,
        64'h8d2300e7_8ca30007,
        64'h8ba30007_8b230460,
        64'h071300e7_8c230210,
        64'h071300e7_85a37522,
        64'h47416786_e8350005,
        64'h041bf59f_e0ef1028,
        64'h040b9963_4c850027,
        64'h4b8306f4_04a306d4,
        64'h07a30087_d79b0086,
        64'hd69b0107_d79b0106,
        64'hd69b0107_979b06f4,
        64'h04232781_0107d79b,
        64'h0107969b_06f40723,
        64'h478100f6_93635714,
        64'h00d61663_57d20007,
        64'h4603468d_05740aa3,
        64'h772280ef_e0ef0544,
        64'h051385d2_049404a3,
        64'h05640423_053407a3,
        64'h05540723_040405a3,
        64'h04040523_03740a23,
        64'h02000613_04f406a3,
        64'h0084d49b_0089d99b,
        64'h04600793_0ff97a93,
        64'h04f40623_02e00b93,
        64'h0104d49b_02100793,
        64'h0109d99b_02f40fa3,
        64'h0104949b_0109199b,
        64'h0ff4fb13_47c12481,
        64'h88cfe0ef_85520200,
        64'h0593462d_898fe0ef,
        64'h85520005_0c1b4581,
        64'h20000613_03440a13,
        64'hf6efe0ef_85220109,
        64'h549b85ca_74221604,
        64'h14630005_041ba98f,
        64'he0ef7522_16f90b63,
        64'h440557fd_16f90f63,
        64'h44094785_18090263,
        64'h0005091b_b45fe0ef,
        64'h45817522_18079f63,
        64'h0207f793_00b7c783,
        64'h441967a6_1af41763,
        64'h47911c04_09630005,
        64'h041bd67f_e0efe4be,
        64'h1028083c_65a21c04,
        64'h14630005_041bbd0f,
        64'he0efe8ea_ece6f0e2,
        64'hf4def8da_fcd6e152,
        64'he54ee94a_ed26f506,
        64'hf1221028_002c4605,
        64'he42a7171_b769d575,
        64'h250191cf_f0ef85a2,
        64'h7502bf61_2501f20f,
        64'he0ef7502_e411f155,
        64'h25019f5f_e0ef1008,
        64'hfaf518e3_4791d94d,
        64'h2501836f_f0ef00a8,
        64'h4581f161_2501951f,
        64'he0efcaa2_00a84589,
        64'h96cfe0ef_00a8100c,
        64'h02800613_fc878de3,
        64'h01492783_c89d88c1,
        64'hcc0d0005_041bad8f,
        64'he0ef0009_45037902,
        64'h80826149_794674e6,
        64'h640a60aa_451dcb81,
        64'h0014f793_00b5c483,
        64'hc59975e2_eb890207,
        64'hf79300b7_c7834519,
        64'h6786e105_2501e3bf,
        64'he0efe0be_1008081c,
        64'h65a2e905_2501ca0f,
        64'he0eff8ca_fca6e122,
        64'he5061008_002c4605,
        64'he42a7175_b7b100f4,
        64'h0523fbf7_f79300a4,
        64'h4783f55d_25016ec0,
        64'h40ef0304_05930017,
        64'hc5034685_4c50601c,
        64'hdba50407_f79300a4,
        64'h4783fcf9_6ae34d1c,
        64'h6008fcf9_00e34509,
        64'h4785b769_449db7e1,
        64'h2501a1cf_f0ef85ca,
        64'h6008f979_2501b37f,
        64'he0ef167d_10000637,
        64'h4c0cb7dd_450502f9,
        64'h146357fd_0005091b,
        64'h94dfe0ef_4c0cbf7d,
        64'h84aa00a4_05a3c539,
        64'h00042a23_2501a58f,
        64'hf0ef484c_ef016008,
        64'h00f40523_c8180207,
        64'he793fed7_72e34814,
        64'h4458cf39_0027f713,
        64'h00a44783_80826105,
        64'h64a26902_85266442,
        64'h60e20007_849bcb91,
        64'h00b44783_e4910005,
        64'h049bbc4f_e0ef842a,
        64'he04aec06_e426e822,
        64'h1101bfad_8a2abfbd,
        64'h4a09b749_4a05b7c5,
        64'h39f10911_2485e111,
        64'h65820155_75332501,
        64'habcfe0ef_e02e854a,
        64'hb745fc0c_94e33cfd,
        64'h39f90909_2485e391,
        64'h8fd90087_979b0009,
        64'h47030019_4783038b,
        64'h91632000_09930344,
        64'h091385ce_e9212501,
        64'hd10fe0ef_0015899b,
        64'h85220009_9e631afd,
        64'h4c094481_49814901,
        64'h10000ab7_504cb74d,
        64'h009b2023_00f402a3,
        64'h0017e793_c8040054,
        64'h4783fef9_63e32905,
        64'h4c1c2485_e1110955,
        64'h08630935_08632501,
        64'ha55fe0ef_852285ca,
        64'h4a8559fd_44814909,
        64'h02fb9f63_47850004,
        64'h4b838082_61656ce2,
        64'h7c027ba2_7b427ae2,
        64'h6a0669a6_694664e6,
        64'h85527406_70a600fb,
        64'h202302f7_6263ffec,
        64'h871b481c_01842c83,
        64'h6000000a_1c630005,
        64'h0a1be7cf_e0efec66,
        64'hf062f45e_fc56e4ce,
        64'he8caeca6_f486e0d2,
        64'h8522002c_46018b2e,
        64'he42af85a_8432f0a2,
        64'h7159bfcd_44198082,
        64'h616564e6_740670a6,
        64'h8522c10f_e0ef1028,
        64'h85a6c489_cf816786,
        64'he8010005_041b872f,
        64'hf0efe4be_1028083c,
        64'h65a2e00d_0005041b,
        64'hedafe0ef_f486f0a2,
        64'h1028002c_460184ae,
        64'he42aeca6_7159bf65,
        64'h84aad16d_bf7d0004,
        64'h2a2300f5_16634791,
        64'h2501f8bf_e0ef8522,
        64'h4581c68f_e0ef8522,
        64'h85ca0004_2a2302f5,
        64'h13634791_2501b32f,
        64'hf0ef8522_45810224,
        64'h30238082_614564e2,
        64'h69428526_740270a2,
        64'h0005049b_c5ffe0ef,
        64'h85224581_00091f63,
        64'he8890005_049bd98f,
        64'he0ef892e_842af406,
        64'he84aec26_f0227179,
        64'h80820141_640260a2,
        64'h00043023_e1192501,
        64'hdbafe0ef_842ae406,
        64'he0221141_b7c1fcf5,
        64'h01e34791_bfdd4525,
        64'h80826121_744270e2,
        64'hf971fcf5_0be34791,
        64'h2501cbdf_e0ef00f4,
        64'h14230067_d7838522,
        64'h458167e2_c448e30f,
        64'he0ef0007_c50367e2,
        64'ha02d0004_30234515,
        64'he7898bc1_00b5c783,
        64'hcd996c0c_e5292501,
        64'h97cff0ef_f01c101c,
        64'he01c8522_65a267e2,
        64'he1152501_fe6fe0ef,
        64'h0828002c_4601842a,
        64'hc52de42e_f822fc06,
        64'h7139b7bd_c45c0137,
        64'h87bb4134_84bbcc0c,
        64'h445cfaf5_fae34f9c,
        64'h601cfaba_fee3fd45,
        64'h88e30005_059bc4bf,
        64'he0efbf69_84cee599,
        64'h0005059b_fddfe0ef,
        64'hcb818b89_600800a4,
        64'h4783b765_cc0cc84c,
        64'hb5ed4905_00f405a3,
        64'h478500f5_976357fd,
        64'hbded4909_00f405a3,
        64'h478900f5_97634785,
        64'h0005059b_814ff0ef,
        64'he595484c_bfb19ca9,
        64'h0094d49b_cd112501,
        64'hc87fe0ef_6008d7b5,
        64'h1ff4f793_c45c9fa5,
        64'h445c0499_ea634a85,
        64'h5a7dd1c1_9c9dc45c,
        64'h27814c0c_8ff94130,
        64'h07bb02c6_ed630337,
        64'h563b0336_d6bbfff4,
        64'h869b377d_c7290097,
        64'h999b0025_47836008,
        64'hbf59cc44_ed352501,
        64'h2bd040ef_85ce0017,
        64'hc5038626_4685601c,
        64'h00f40523_fbf7f793,
        64'h00a44783_ed512501,
        64'h30f040ef_0017c503,
        64'h85ce4685_601cc385,
        64'h0407f793_03040993,
        64'h00a44783_fc960ee3,
        64'h4c50d3e5_1ff7f793,
        64'h445c4481_bf7d00f4,
        64'h05230207_e79300a4,
        64'h4783c81c_fcf778e3,
        64'h4818445c_e4bd0004,
        64'h26234458_84bae391,
        64'h8b8900a4_47830097,
        64'h77634818_80826121,
        64'h6aa26a42_69e27902,
        64'h74a2854a_744270e2,
        64'h0007891b_cf8900b4,
        64'h47830009_17630005,
        64'h091bfb4f_e0ef84ae,
        64'h842ae456_e852ec4e,
        64'hfc06f04a_f426f822,
        64'h7139b709_fe9465e3,
        64'hfee78fa3_24050785,
        64'h00074703_97369281,
        64'h02041693_67220789,
        64'hbddd4545_b7e900c6,
        64'h8023377d_fc964603,
        64'h962a1088_92010207,
        64'h1613b7c1_2785b731,
        64'h9c3d0136_8023fff7,
        64'hc7930127_1a6396b2,
        64'h920166a2_02069613,
        64'h00e586bb_40f405bb,
        64'hfff7871b_04e46263,
        64'h0037871b_eb05fc97,
        64'h47039736_10949301,
        64'h02079713_4781f5cf,
        64'he0ef1828_100cb759,
        64'h4509f8e5_16e367a2,
        64'h4711dd61_2501a9ef,
        64'hf0ef1828_45810145,
        64'h0e632501_8a7fe0ef,
        64'h0007c503_65c677e2,
        64'he1052501_e48ff0ef,
        64'h18284581_f9492501,
        64'hf63fe0ef_18284581,
        64'hc2aa8cdf_e0ef0007,
        64'hc50365c6_77e2f555,
        64'h2501e6ef_f0ef1828,
        64'h4581fd45_2501f89f,
        64'he0ef1828_45858082,
        64'h61497a06_79a67946,
        64'h74e6640a_60aa0007,
        64'h8023078d_00e78123,
        64'h02f00713_0e941863,
        64'h00e780a3_03a00713,
        64'h00e78023_0307071b,
        64'h53874703_00008717,
        64'he50567a2_4501040a,
        64'h12634a16_c2be02f0,
        64'h09934bdc_597d8426,
        64'h77e2ecbe_081ce529,
        64'h2501acdf_e0ef1828,
        64'h002c4601_84ae0005,
        64'h0023f0d2_f4cef8ca,
        64'he122e506_e42afca6,
        64'h7175bfd9_4415fcf4,
        64'h1ee34791_b7c5c8c8,
        64'h97bfe0ef_0004c503,
        64'h74a2cb99_8bc100b5,
        64'hc7838082_616564e6,
        64'h740670a6_8522cbd8,
        64'h575277a2_e9916586,
        64'he41d0005_041bcd2f,
        64'hf0efe4be_1028083c,
        64'h65a2ec19_0005041b,
        64'hb3bfe0ef_eca6f486,
        64'hf0a21028_002c4601,
        64'he42a7159_bfe5452d,
        64'h80826105_60e24501,
        64'h5ea78823_00008797,
        64'h00054a63_95bfe0ef,
        64'hec060028_e42a1101,
        64'h80820141_640260a2,
        64'h00043023_e1192501,
        64'h9cbfe0ef_8522e901,
        64'h2501efff_f0ef842a,
        64'he406e022_11418082,
        64'h01416402_60a24505,
        64'hebbfe06f_014160a2,
        64'h640200f5_02234785,
        64'h00f40523_fdf7f793,
        64'h600800a4_47830007,
        64'h89a30007_892300e7,
        64'h8ca300d7_8da30460,
        64'h07130086_d69b00e7,
        64'h8c230210_07130106,
        64'hd69b00e7_8aa30087,
        64'h571b0107_571b0107,
        64'h171b00e7_8a232701,
        64'h0107571b_0107169b,
        64'h00e78d23_00078ba3,
        64'h00078b23_485800e7,
        64'h8fa300d7_8f230187,
        64'h571b0107_569b00d7,
        64'h8ea300e7_8e230086,
        64'hd69b0106_d69b0107,
        64'h169b4818_00e785a3,
        64'h02076713_00b7c703,
        64'h741ce15d_2501b77f,
        64'he0ef6008_500c00f4,
        64'h0523fbf7_f79300a4,
        64'h4783ed55_25016850,
        64'h40ef0304_05930017,
        64'hc5034685_4c50601c,
        64'hc3950407_f793cf69,
        64'h0207f713_00a44783,
        64'he1752501_acffe0ef,
        64'h842ae406_e0221141,
        64'hbd2d499d_b5f9c81c,
        64'hbf4100f4_05230407,
        64'he79300a4_47839dbf,
        64'he0ef9522_85d28626,
        64'h03050513_0007849b,
        64'h0127f463_40ab87bb,
        64'h1ff57513_0009049b,
        64'h444801a4_2e23fd09,
        64'h25016c70_40ef85da,
        64'h4685001d_c50300e7,
        64'hfa63445c_481800c7,
        64'h8e634c5c_bdd100fa,
        64'ha0239fa5_000aa783,
        64'hc45c9fa5_4099093b,
        64'h445c9a3e_93810204,
        64'h97930094_949b00f4,
        64'h0523fbf7_f79300a4,
        64'h4783a4ff_e0ef855a,
        64'h95d22000_06139181,
        64'h15820097_959b0297,
        64'hf26341a5_87bb4c4c,
        64'hf1512501_763040ef,
        64'h85d286a6_001dc503,
        64'h419704bb_00f77463,
        64'h9fb5002d_c703c4b5,
        64'h8d320007_849b00a6,
        64'h863b0099_579b000c,
        64'h869bd159_250197cf,
        64'hf0ef856e_4c0c0004,
        64'h3d8300f4_0523fbf7,
        64'hf79300a4_4783f969,
        64'h25017b10_40ef85da,
        64'h0017c503_46854c50,
        64'h601cc38d_0407f793,
        64'h00a44783_c85ce311,
        64'hcc1c4858_bf994985,
        64'h00f405a3_47850187,
        64'h9763b795_00f40523,
        64'h0207e793_00a44783,
        64'h12f76a63_4818445c,
        64'hf3fd0005_079bd86f,
        64'hf0ef4c0c_b7594989,
        64'h00f405a3_478902e7,
        64'h98634705_cb914581,
        64'h485cef01_040c9a63,
        64'h0ffcfc93_0197fcb3,
        64'h37fd0025_47830097,
        64'h5c9b6008_14079363,
        64'h1ff77793_04090463,
        64'h44585c7d_03040b13,
        64'h20000b93_04f76c63,
        64'h0127873b_445c1807,
        64'h8f638b89_00a44783,
        64'h80826165_6da26d42,
        64'h6ce27c02_7ba27b42,
        64'h7ae26a06_69a66946,
        64'h64e6854e_740670a6,
        64'h0007899b_c39d00b4,
        64'h47830009_97630005,
        64'h099bcb5f_e0ef8ab6,
        64'h89328a2e_842a0006,
        64'ha023e46e_e86aec66,
        64'hf062f45e_f85aeca6,
        64'hf486fc56_e0d2e4ce,
        64'he8caf0a2_7159b59d,
        64'h499dbf9d_bd1fe0ef,
        64'h855295a2_86260305,
        64'h85930007_849b0127,
        64'hf46340bb_87bb1ff5,
        64'hf5930009_049b444c,
        64'h01a42e23_f1152501,
        64'h0bc050ef_85da0017,
        64'hc503863a_4685601c,
        64'h00f40523_fbf7f793,
        64'h672200a4_4783f139,
        64'h25011100_50efe43a,
        64'h85da4685_001dc503,
        64'hc38d0407_f79300a4,
        64'h478304e6_01634c50,
        64'hb70500fa_a0239fa5,
        64'h000aa783_c45c9fa5,
        64'h4099093b_445c9a3e,
        64'h93810204_97930094,
        64'h949bc5ff_e0ef9552,
        64'h85da2000_06139101,
        64'h15020097_951b0097,
        64'hfc6341a5_07bb4c48,
        64'hc3850407_f79300a4,
        64'h4783f94d_250114a0,
        64'h50ef85d2_863a86a6,
        64'h001dc503_419684bb,
        64'h00f6f463_9fb1002d,
        64'hc683c4b5_8d3a0007,
        64'h849b00a6_073b0099,
        64'h579b000c_861bd579,
        64'h2501b98f_f0ef856e,
        64'h4c0c0004_3d83cc08,
        64'hb7a54985_00f405a3,
        64'h47850185_1763b7e5,
        64'h2501bd6f_f0ef4c0c,
        64'hb7414989_00f405a3,
        64'h478900a7_ec634785,
        64'h4848eb11_020c9963,
        64'h0ffcfc93_0197fcb3,
        64'h37fd0025_47830097,
        64'h5c9b6008_12079063,
        64'h1ff77793_4458fa09,
        64'h0ce35c7d_03040b13,
        64'h20000b93_0006091b,
        64'h00f67463_893e40f9,
        64'h07bb445c_01042903,
        64'h16078963_8b8500a4,
        64'h47838082_61096de2,
        64'h7d027ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_854e7446,
        64'h70e60007_899bc39d,
        64'h662200b4_47830009,
        64'h98630005_099be91f,
        64'he0ef8ab6_e4328a2e,
        64'h842a0006_a023ec6e,
        64'hf06af466_f862fc5e,
        64'he0daf0ca_f4a6fc86,
        64'he4d6e8d2_eccef8a2,
        64'h7119b7d5_491db7e5,
        64'h49118082_61496b46,
        64'h6ae67a06_79a67946,
        64'h74e6854a_640a60aa,
        64'h00f49423_0134b023,
        64'h0004ae23_0004a623,
        64'hc8880069_d783dbbf,
        64'he0ef01c4_0513c8c8,
        64'hf33fe0ef_0009c503,
        64'h000485a3_d09c0144,
        64'h8523f480_0309a783,
        64'h85a279a2_020a6a13,
        64'hc399008a_7793e3ad,
        64'h8b850009_84630029,
        64'hf993e72d_0107f713,
        64'h00b44783_f565a085,
        64'h4921f609_81e30049,
        64'hf993e3d9_8bc500b4,
        64'h4783a895_892ac90d,
        64'h250183af_f0ef0135,
        64'h262385da_39fd7522,
        64'he9112501_e3fff0ef,
        64'h030aab03_855685ce,
        64'h04098b63_00fa8223,
        64'h0005099b_00040aa3,
        64'h00040a23_00040da3,
        64'h00040d23_4785fc9f,
        64'he0ef85a2_000ac503,
        64'h00040fa3_00040f23,
        64'h00040ea3_00040e23,
        64'h000405a3_00e40c23,
        64'h00040ba3_00040b23,
        64'h00e40823_000407a3,
        64'h00040723_00f40ca3,
        64'h00f408a3_02100713,
        64'h04600793_7aa2cfcd,
        64'h008a7793_6406e949,
        64'h008a6a13_2501e75f,
        64'hf0ef1028_00f51663,
        64'h4791c54d_c3e101f9,
        64'hfa1301c9_f7934519,
        64'he011e119_64062501,
        64'hb6dff0ef_e4be1028,
        64'h083c65a2_14091063,
        64'h0005091b_9d6ff0ef,
        64'h1028002c_8a7984aa,
        64'h89b20005_30231405,
        64'h0d634925_e42ee8da,
        64'hecd6f0d2_f4cefca6,
        64'he122e506_f8ca7175,
        64'hbfe5452d_80826121,
        64'h70e22501_a0eff0ef,
        64'h0828080c_460100f6,
        64'h18634785_cb114501,
        64'he39897aa_00070023,
        64'hc3196762_00070023,
        64'hc3196622_631800a7,
        64'h8733050e_cc478793,
        64'h00009797_04054263,
        64'h83eff0ef_f42ee432,
        64'he82efc06_1028ec2a,
        64'h7139b759_4505bf5d,
        64'h0009049b_00f402a3,
        64'h0017e793_00544783,
        64'hc81c2785_01378a63,
        64'h481cf15d_25018aff,
        64'hf0ef8522_85a64601,
        64'h03390763_fb490ce3,
        64'hbf754501_00091463,
        64'h0005091b_ec8ff0ef,
        64'h852285a6_00f4fa63,
        64'h4c1c59fd_4a05fcf5,
        64'hfde384ae_842ae052,
        64'he44ee84a_f406ec26,
        64'hf0227179_4d1c8082,
        64'h61456a02_69a26942,
        64'h64e27402_70a24509,
        64'h80824509_00b7ed63,
        64'h47858082_610564a2,
        64'h85266442_60e200e7,
        64'h82234705_601c82af,
        64'hf0ef462d_6c08700c,
        64'h84cff0ef_45810200,
        64'h06136c08_e0850005,
        64'h049ba42f_f0ef6008,
        64'h484ce49d_0005049b,
        64'hfa9ff0ef_842aec06,
        64'he426e822_11018082,
        64'h610564a2_644260e2,
        64'h451d00f5_13634791,
        64'hdd792501_bcdff0ef,
        64'h85224585_cb990097,
        64'h8d630007_c7836c1c,
        64'hed092501_a8cff0ef,
        64'h6008484c_0e500493,
        64'he50d2501_88fff0ef,
        64'h842ae426_ec06e822,
        64'h45811101_bfe54511,
        64'hb7cd0004_2a23d945,
        64'h2501c13f_f0ef8522,
        64'h45818082_614569a2,
        64'h694264e2_740270a2,
        64'h45010097_9a630017,
        64'hb79317e1_8bfd0337,
        64'h80630327_026303f7,
        64'hf79300b7_c783c321,
        64'h0007c703_6c1ce129,
        64'h2501afaf_f0ef6008,
        64'ha0b1c90d_e199484c,
        64'h49bd0e50_09134511,
        64'h84aef406_842ae44e,
        64'he84aec26_f0227179,
        64'hbdf90ff7_77130017,
        64'he7933701_eea866e3,
        64'h0ff57513_f9f7051b,
        64'heea87ae3_0ff57513,
        64'hfbf7051b_bd6d4519,
        64'hf11710e3_00088663,
        64'h00054883_0c450513,
        64'h00008517_00054c63,
        64'h4185551b_0187151b,
        64'h02b6f263_fd370ae3,
        64'hf95704e3_f94706e3,
        64'hf4e374e3_00074703,
        64'h97229301_17020017,
        64'h061b8732_45ad46a1,
        64'h0ff7f793_0027979b,
        64'h05659a63_bdb9c4c8,
        64'haf2ff0ef_0007c503,
        64'h609cdbe5_8bc100b5,
        64'hc7836c8c_fbf58b91,
        64'hb73d4515_fb0dbf15,
        64'h4501e807_03e30004,
        64'hbc230004_a623cb89,
        64'h0207f793_0047f713,
        64'hf4e518e3_4711c505,
        64'h00b7c783_709c4511,
        64'hbf654701_bdfd00e9,
        64'h05a39432_92011602,
        64'h00876713_00d79463,
        64'h46918bb1_01076713,
        64'h00b69463_45850037,
        64'hf6930ff7_f7930027,
        64'h979b0165_966300d9,
        64'h00234695_00d51563,
        64'h0e500693_00094503,
        64'hc6ed4711_a06d2685,
        64'h00e50023_954a9101,
        64'h02069513_0027e793,
        64'ha8dd0505_a0d14865,
        64'h02000313_478145a1,
        64'h47014681_b7ad0240,
        64'h0793943a_12f6e063,
        64'h02000693_f7578be3,
        64'hbf954709_bf1d0405,
        64'h80826121_6b026aa2,
        64'h6a4269e2_790274a2,
        64'h744270e2_0004bc23,
        64'h2501a85f_f0ef8526,
        64'h4581b791_c55c4bdc,
        64'h611cbf75_dfdff0ef,
        64'h85264581_fed608e3,
        64'hfff7c683_fff74603,
        64'h07850705_0cb78d63,
        64'h00b78593_709cef91,
        64'h8ba100b7_4783c7e5,
        64'h00074783_6c98e96d,
        64'h2501cdaf_f0ef6088,
        64'h48cc1005_10632501,
        64'hadbff0ef_85264581,
        64'h00f905a3_02000793,
        64'h943a0947_9763470d,
        64'h1b378e63_00244783,
        64'h00f900a3_02e00793,
        64'h0b379063_00144783,
        64'h01390023_0d379263,
        64'h00044783_b40ff0ef,
        64'h854a0200_0593462d,
        64'h0204b903_0d578063,
        64'h0d478263_00044783,
        64'h4b2102e0_099305c0,
        64'h0a9302f0_0a130ae7,
        64'hfc6347fd_00044703,
        64'h0004a623_04050ce7,
        64'h906305c0_071300e7,
        64'h8663842e_84aa02f0,
        64'h07130005_c783e05a,
        64'he456e852_ec4ef04a,
        64'hfc06f426_f8227139,
        64'hb7e9db1c_27855b1c,
        64'h2a856018_f1412501,
        64'hd1cff0ef_01450223,
        64'hb7b9c848_a83ff0ef,
        64'h85a6c804_6008d91c,
        64'h415787bb_591c00fa,
        64'hed630025_47836008,
        64'h4a0502aa_2823aa5f,
        64'hf0ef8552_85a60004,
        64'h3a03beef_f0ef0345,
        64'h05134581_20000613,
        64'h6008f579_2501dd8f,
        64'hf0ef6008_fcf48de3,
        64'h57fdfcf4_8be34785,
        64'hd4bd451d_0005049b,
        64'he81ff0ef_480cf60a,
        64'h0ee306f4_e0634d1c,
        64'h6008b761_450500f4,
        64'h946357fd_bf494509,
        64'h0097e463_47850005,
        64'h049bb27f_f0effc0a,
        64'h9fe30157_fab337fd,
        64'h00495a9b_00254783,
        64'hbf5d4501_ec1c97ce,
        64'h03478793_01241523,
        64'h0996601c_fcf775e3,
        64'h0009071b_00855783,
        64'he18dc85c_61082785,
        64'h480c0009_9d63842a,
        64'h8a2e00f9_7993d7ed,
        64'h495c8082_61216aa2,
        64'h6a4269e2_790274a2,
        64'h744270e2_4511eb99,
        64'h93c1e456_e852ec4e,
        64'hf4260309_17932905,
        64'hf822fc06_00a55903,
        64'hf04a7139_bfad4405,
        64'hf6f50fe3_4785dd61,
        64'h2501dbbf_f0ef8526,
        64'h85ce8622_bf4900f4,
        64'h82a30017_e7930054,
        64'hc783c89c_37fdfae7,
        64'h83e3577d_c4c0489c,
        64'h02099063_e9052501,
        64'hde9ff0ef_852685a2,
        64'h167d1000_0637b76d,
        64'hfb2411e3_05450863,
        64'hfd5507e3_c9012501,
        64'hc05ff0ef_852685a2,
        64'h4409bf55_4905b7d5,
        64'hfaf47ee3_894e4c9c,
        64'h80826121_6aa26a42,
        64'h69e27902_74a27442,
        64'h70e28522_547d00f4,
        64'h1d6357fd_0887f863,
        64'h47850005_041bc43f,
        64'hf0efa821_4401052a,
        64'h606304f4_63632405,
        64'h4c9c5afd_4a05844a,
        64'h04f97763_4d1c0409,
        64'h0a6300c5_2903e19d,
        64'h89ae84aa_e456e852,
        64'hf04af822_fc06ec4e,
        64'hf4267139_bf3d4989,
        64'hb745012a_81a300fa,
        64'h81230189_591b0109,
        64'h579b00fa_80a30087,
        64'hd79b0324_0a230107,
        64'hd79b9426_0109179b,
        64'h01256933_8d71f000,
        64'h06372501_da0ff0ef,
        64'h85569aa6_03440a93,
        64'h1fc47413_0024141b,
        64'hf80996e3_0005099b,
        64'hfd8ff0ef_9dbd0075,
        64'hd59b515c_bf790144,
        64'h82230324_0aa30089,
        64'h591b0109_591b0109,
        64'h191b0324_0a239426,
        64'h1fe47413_0014141b,
        64'hfc0992e3_0005099b,
        64'h811ff0ef_9dbd0085,
        64'hd59b515c_b7e90127,
        64'he9339bc1_00f97913,
        64'h0089591b_0347c783,
        64'h015487b3_80826121,
        64'h6aa26a42_69e27902,
        64'h74a2854e_744270e2,
        64'h00f48223_4785032a,
        64'h8a239aa6_0ff97913,
        64'h0049591b_c40d1ffa,
        64'hfa930009_9f630005,
        64'h099b86bf_f0ef9dbd,
        64'h8526009a_d59b50dc,
        64'h00f48223_478502fa,
        64'h0a239a26_0ff7f793,
        64'h8fd98ff5_0049179b,
        64'h00f7f713_16c16685,
        64'h0347c783_014487b3,
        64'hcc191ffa_7a130ff9,
        64'h7793001a_0a9b8805,
        64'h06099663_0005099b,
        64'h8b9ff0ef_9dbd009a,
        64'h559b00ba_0a3b515c,
        64'h0015da1b_15479463,
        64'h0ee78863_470d0ae7,
        64'h8f63842e_89324709,
        64'h00054783_0af5f063,
        64'h498984aa_4d1c16ba,
        64'h75634a05_e456ec4e,
        64'hf04af426_f822fc06,
        64'he8527139_80826105,
        64'h64a28526_644260e2,
        64'h00e78223_4705601c,
        64'h00e78023_57156c1c,
        64'hf3cff0ef_45810200,
        64'h06136c08_ec990005,
        64'h049b933f_f0ef6008,
        64'h484ce495_0005049b,
        64'hf33ff0ef_842aec06,
        64'he426e822_110100a5,
        64'h5583b78d_4505bfc1,
        64'h413484bb_f6f476e3,
        64'h4f9c0009_3783f68a,
        64'hfbe30144_0c630005,
        64'h041be6ff_f0efbf75,
        64'h2501e59f_f0ef0134,
        64'hf66385a2_00093503,
        64'h4a850992_5a7d843a,
        64'h0027c983_8722b75d,
        64'h45010099_3c2300a9,
        64'h2a2394be_03478793,
        64'h049688bd_00093783,
        64'h9d3d0044_d79bd171,
        64'h00892823_5788fce4,
        64'hf7e30087_d703eb15,
        64'h579800e6_9463470d,
        64'h0007c683_e02184ae,
        64'hfee474e3_4f98611c,
        64'h80826121_6aa26a42,
        64'h69e27902_74a27442,
        64'h70e24509_00f41c63,
        64'h892a4785_00b51523,
        64'he456e852_ec4ef426,
        64'hfc06f04a_4540f822,
        64'h71398082_853e4785,
        64'hb76517fd_25011000,
        64'h07b7807f_f0ef954a,
        64'h03450513_1fc57513,
        64'h0024151b_f9352501,
        64'ha39ff0ef_9dbd0075,
        64'hd59b515c_b7598fc9,
        64'h0087979b_03494503,
        64'h03594783_99221fe4,
        64'h74130014_141bfd59,
        64'h2501a63f_f0ef9dbd,
        64'h0085d59b_515cbf45,
        64'h8fe9157d_6505bf65,
        64'h8391c019_8fc50087,
        64'h979b8805_03494783,
        64'h994e1ff9_f993f579,
        64'h2501a93f_f0ef0344,
        64'hc483854a_9dbd94ca,
        64'h1ff4f493_0099d59b,
        64'h0014899b_02492783,
        64'h80826145_853e69a2,
        64'h694264e2_740270a2,
        64'h57fdc911_2501ac7f,
        64'hf0ef9dbd_0094d59b,
        64'h9cad515c_0015d49b,
        64'h00f71e63_08d70e63,
        64'h468d06d7_0c63842e,
        64'h46890005_470302e5,
        64'hf963892a_e44eec26,
        64'hf022f406_e84a7179,
        64'h4d180eb7_f7634785,
        64'h80824501_80829d2d,
        64'h02d585bb_55480025,
        64'h458300f6_f96337f9,
        64'hffe5869b_4d1c8082,
        64'h610564a2_644260e2,
        64'h00a03533_25016310,
        64'h50ef4581_46010014,
        64'h45030004_02a363d0,
        64'h50ef85a6_4685d810,
        64'h22f401a3_22e40123,
        64'h20d40ca3_20d40c23,
        64'h0187d79b_0107d71b,
        64'h260522e4_00a322f4,
        64'h00230720_06930014,
        64'h45030087_571b0107,
        64'h571b0107_971b5010,
        64'h20e40f23_445c20f4,
        64'h0fa30187_d79b0107,
        64'hd71b20e4_0ea320f4,
        64'h0e230087_571b0107,
        64'h571b0107_971b20e4,
        64'h0d2302e4_0ba30410,
        64'h0713481c_20f40da3,
        64'h02f40b23_06100793,
        64'h02f40aa3_02f40a23,
        64'h05200793_22f409a3,
        64'hfaa00793_22f40923,
        64'h05500793_a01ff0ef,
        64'h85264581_20000613,
        64'h03440493_0af71b63,
        64'h47850054_47030cf7,
        64'h1063478d_00044703,
        64'hed692501_bffff0ef,
        64'h842ae426_ec06e822,
        64'h1101bdc5_9cbd0017,
        64'hd79b8885_029787bb,
        64'h478db701_0014949b,
        64'h00f91563_4789d41c,
        64'h9fb5e00a_05e3b545,
        64'ha25ff0ef_05440513,
        64'hb5b90005_099ba33f,
        64'hf0ef0584_0513b351,
        64'h47810004_2a230124,
        64'h002300f4_13237cf7,
        64'h18230000_971793c1,
        64'h17c22785_7de7d783,
        64'h00009797_c448a63f,
        64'hf0ef2204_0513c808,
        64'ha6dff0ef_21c40513,
        64'h00f51c63_27278793,
        64'h25016141_77b7a83f,
        64'hf0ef2184_051302f5,
        64'h17632527_87932501,
        64'h416157b7_a99ff0ef,
        64'h03440513_04f71263,
        64'ha5570713_4107d79b,
        64'h776d0107_979b8fd9,
        64'h0087979b_000402a3,
        64'h23244703_23344783,
        64'he13d2501_ce5ff0ef,
        64'h8522001a_859b06f7,
        64'h1b634705_4107d79b,
        64'h0107979b_8fd90087,
        64'h979b0644_47030654,
        64'h478308f9_1963478d,
        64'h00f402a3_f8000793,
        64'hc45cc81c_57fdee99,
        64'he7e32481_0094d49b,
        64'h1ff4849b_0024949b,
        64'hd408b17f_f0ef0604,
        64'h0513f00a_15e310e9,
        64'h1263470d_d05c0354,
        64'h2023cc04_d4580157,
        64'h87bb2489_00ea873b,
        64'h490d00b6_73630905,
        64'h165500b9_39336641,
        64'h19556905_dd8d84ae,
        64'h0364d5bb_40c504bb,
        64'hf4c564e3_873200d7,
        64'h063b9f3d_004a571b,
        64'h27810339_06bbdfb1,
        64'h8fd90087_979b2501,
        64'h04244703_04344783,
        64'h14050e63_8d450085,
        64'h151b0474_44830484,
        64'h4503f3c1_00fa7793,
        64'h01441423_00fa6a33,
        64'h008a1a1b_04544783,
        64'h04644a03_ffc900fb,
        64'h77b3fffb_079bfa0b,
        64'h03e30164_01230414,
        64'h4b03faf7_69e30ff7,
        64'hf7930124_01a3fff9,
        64'h079b4705_01342e23,
        64'h04444903_29811a09,
        64'h866300f9_e9b30089,
        64'h999b04a4_478304b4,
        64'h4983fef7_11e32000,
        64'h07134107_d79b0107,
        64'h979b8fd9_0087979b,
        64'h03f44703_04044783,
        64'hbfb947b5_c1194a81,
        64'hf6e504e3_4785470d,
        64'hb7bd00e5_19634785,
        64'h470dfe99_15e30491,
        64'hc10de9df_f0ef8522,
        64'h85d6000a_87634509,
        64'h0004aa83_01048913,
        64'hff2a14e3_09910941,
        64'h00a9a023_2501c5bf,
        64'hf0ef854a_c7894501,
        64'hffc94783_89a623a4,
        64'h0a131fa4_0913848a,
        64'h04f51a63_4785ee1f,
        64'hf0ef8522_4581f569,
        64'h89110009_0463fb71,
        64'h478d0015_77130f40,
        64'h60ef00a4_00a30004,
        64'h00230ff4_f5138082,
        64'h6161853e_6b426ae2,
        64'h7a0279a2_794274e2,
        64'h640660a6_47a9c111,
        64'h89110009_0563e38d,
        64'h00157793_1e2060ef,
        64'h00144503_cb850004,
        64'h47830089_b023c015,
        64'h47b184aa_638097ba,
        64'ha5878793_0000a797,
        64'h00351713_02054e63,
        64'h47addd9f_f0ef8932,
        64'h852e89aa_00053023,
        64'he85aec56_f052fc26,
        64'he0a2e486_f44ef84a,
        64'h715dbfcd_450d8082,
        64'h61056902_64a26442,
        64'h60e200a0_35338d05,
        64'h01257533_2501d33f,
        64'hf0ef0864_05130097,
        64'h8c634501_0127f7b3,
        64'h14650493_00544537,
        64'hfff50913_01000537,
        64'h0005079b_d59ff0ef,
        64'h06a40513_02f71f63,
        64'ha5570713_4107d79b,
        64'h776d0107_979b8fd9,
        64'h0087979b_45092324,
        64'h47032334_4783e52d,
        64'h2501fa3f_f0ef842a,
        64'hd91c0005_022357fd,
        64'he04ae426_ec06e822,
        64'h11018082_61056902,
        64'h64a26442_60e28522,
        64'h0324a823_597d4405,
        64'hc1192501_298060ef,
        64'h03448593_864a4685,
        64'h0014c503_ec190005,
        64'h041bfddf_f0ef892e,
        64'h84aa02b7_87634401,
        64'he04ae426_ec06e822,
        64'h1101591c_80824501,
        64'hf8dff06f_c3990045,
        64'h4783b7f9_4505b7e5,
        64'h397d3100_60ef85ce,
        64'h86269cbd_46850014,
        64'h45034c5c_ff2a74e3,
        64'h4a050034_49038082,
        64'h61456a02_69a26942,
        64'h64e27402_70a24501,
        64'h00e7eb63_40f487bb,
        64'h00040223_4c58505c,
        64'he1312501_352060ef,
        64'h85ce8626_46850015,
        64'h4503842a_03450993,
        64'he052e84a_f4065904,
        64'he44eec26_f0227179,
        64'h8082853e_27818fd9,
        64'h0107979b_8fd50087,
        64'h979b0145_c6830155,
        64'hc78300d5_1d630007,
        64'h079b8f5d_0087979b,
        64'h468d01a5_c70301b5,
        64'hc7838082_45258082,
        64'h014160a2_4525c391,
        64'h45010015_77933c40,
        64'h60ef0017_c503e406,
        64'h114102e6_90630085,
        64'h57030067_d683c70d,
        64'h0007c703_cb85611c,
        64'hc915bfd5_c5474703,
        64'h0000a717_8082853a,
        64'he11c0006_871b0789,
        64'h00b66663_0ff6f593,
        64'hfd06869b_577d4605,
        64'h0007c683_b7dd0705,
        64'ha00d577d_00d70663,
        64'h00178693_00c69863,
        64'h02d5fc63_00074683,
        64'h03a00613_02000593,
        64'hcf99873e_611c8082,
        64'h61056902_64a26442,
        64'h60e20004_002300f4,
        64'h93238fd9_0087979b,
        64'h01694703_01794783,
        64'h00f49223_8fd90087,
        64'h979b0189_47030199,
        64'h4783c088_f59ff0ef,
        64'h00f58423_84ae01c9,
        64'h051300b9_4783fcc7,
        64'h9ee30685_040500e4,
        64'h00230405_00640023,
        64'h01179563_0e500713,
        64'h01071463_00a70e63,
        64'h27850006_c703462d,
        64'h02e00313_48a54815,
        64'h86ca0200_05134781,
        64'h01853903_cfa50095,
        64'h8413e04a_e426ec06,
        64'he8221101_495cbfcd,
        64'h050500b5_00238082,
        64'h00f61363_367d57fd,
        64'hb7f5fee5_0fa30585,
        64'h05050005_c7038082,
        64'h00f61363_367d57fd,
        64'h80822501_8d5d0562,
        64'h8fd907c2_00354503,
        64'h00254783_8f5d07a2,
        64'h00054703_00154783,
        64'hb7d914fd_b7e9b9ff,
        64'hf0efbfc1_710a8493,
        64'h77d050ef_4501dff1,
        64'h54fd000a_2783bfc5,
        64'hbb9ff0ef_fc075de3,
        64'h03379713_83093783,
        64'h02074563_03379713,
        64'h83093783_5a0b0493,
        64'hedbfe0ef_8522e78d,
        64'h0009a783_e4a9d807,
        64'ha7230000_a797d807,
        64'had230000_a797da07,
        64'ha3230000_a797d807,
        64'haf230000_a797da07,
        64'h95230000_a797dcf7,
        64'h09a30000_a7170054,
        64'h4783dcf7_0f230000,
        64'ha7170044_4783def7,
        64'h04a30000_a7170034,
        64'h4783def7_0a230000,
        64'ha7174300_19370026,
        64'h2b370024_4783e0f7,
        64'h03a30000_a7176a89,
        64'hdf8a0a13_0000aa17,
        64'h00144783_e0f70e23,
        64'h0000a717_e0498993,
        64'h0000a997_44810004,
        64'h4783e2a4_04130000,
        64'ha41707d0_30ef0465,
        64'h05130000_9517e3e5,
        64'hc5830000_a597e476,
        64'h46030000_a617e506,
        64'hc6830000_a697e5b8,
        64'h48030000_a817e627,
        64'hc7830000_a797e697,
        64'h47030000_a7170b90,
        64'h30ef0725_05130000,
        64'h951780e7_b423e05a,
        64'he456e852_ec4ef04a,
        64'hf426f822_fc068f4d,
        64'h91c115c2_00800737,
        64'h71398087_b5838007,
        64'hb6034300_17b7bf91,
        64'hff3410e3_0f7030ef,
        64'hfec48fa3_0ff67613,
        64'h00c95633_0286061b,
        64'h04852405_855285a2,
        64'h028a863b_49990b6a,
        64'h0a130000_9a175ae1,
        64'h4401eda4_84930000,
        64'ha4978082_61616ae2,
        64'h7a0279a2_794274e2,
        64'h82f6b423_47a16406,
        64'h60a68086_b7838006,
        64'hb78380f6_b42393c1,
        64'h80a6b023_17c29101,
        64'h430016b7_8fd91502,
        64'h0ff77713_8ff18321,
        64'h0087179b_f0060613,
        64'h01000637_4722f2ff,
        64'hf0ef4512_7d0050ef,
        64'h0028f3a5_85930000,
        64'ha5974609_7e0050ef,
        64'h0048f4c5_85930000,
        64'ha5974611_f4a78ca3,
        64'h0000a797_fe056513,
        64'h893d0030_70eff6f7,
        64'h05230000_a7175791,
        64'hf6f709a3_0000a717,
        64'h578df6f7_0e230000,
        64'ha7175789_f8f702a3,
        64'h0000a717_5785f8f7,
        64'h07230000_a71757b9,
        64'h0a091d63_c3190107,
        64'h9713fff9_47931f10,
        64'h30ef1825_05130000,
        64'h9517892a_077070ef,
        64'hec56f052_f44efc26,
        64'he0a2f84a_e486c63e,
        64'h04b00513_45854601,
        64'h00740207_879b0700,
        64'h07b7715d_80822501,
        64'h8d5d8d79_00ff0737,
        64'h0085151b_8fd98f75,
        64'h0085571b_f0068693,
        64'h8fd966c1_0185579b,
        64'h0185171b_80829141,
        64'h15428d5d_05220085,
        64'h579b8082_614564e2,
        64'h740270a2_85228d4f,
        64'hf0ef0225_05130000,
        64'ha5170450_069301a7,
        64'h57030000_a7170168,
        64'h88930000_a89785a6,
        64'h862247b2_0007a803,
        64'h03078793_0000a797,
        64'h0ed050ef_f4060068,
        64'h07858593_0000a597,
        64'h461184ae_8432ec26,
        64'hf0227179_bfc14785,
        64'heb9ff0ef_80826105,
        64'h64a26442_60e2c3c0,
        64'h0c2007b7_2cf030ef,
        64'h24850513_00009517,
        64'he7990206_c1630337,
        64'h16938304_b7034300,
        64'h14b74781_2401ec06,
        64'he42643c0_e8220c20,
        64'h07b71101_b7e1ff06,
        64'hbc2306a1_26050008,
        64'h380300d7_88338082,
        64'h61010113_5f813483,
        64'h85266001_34036081,
        64'h30838287_b8234300,
        64'h17b70405_aa1ff0ef,
        64'h862602e6_446397c2,
        64'h85b64300_08378f95,
        64'h868a83f5_02d7473b,
        64'h17822705_46a10077,
        64'h67139fad_377d8005,
        64'h859b6585_02d51a63,
        64'h80668693_6685c691,
        64'h8005069b_00015503,
        64'h00d10023_0086d69b,
        64'h0106d69b_0106969b,
        64'h00d100a3_872646d4,
        64'h96aa068e_9ebd8006,
        64'h869b7007_f7930084,
        64'h179bea25_439014e7,
        64'h87930000_a797cfb5,
        64'h27818ff1_fff7c793,
        64'h00c5963b_10100593,
        64'h8a1d08b8_696335b9,
        64'h5f200813_ffc5849b,
        64'h25816011_34235e91,
        64'h3c23630c_8387b783,
        64'h972a4300_05379f2d,
        64'h8406871b_03877593,
        64'h66850034_171b00f6,
        64'h74132601_60813023,
        64'h9f010113_8307b603,
        64'h430017b7_bba54601,
        64'h40b030ef_36c50513,
        64'h00009517_85aab369,
        64'h00f41623_60800793,
        64'h00f41f23_0024d783,
        64'h00f41e23_0004d783,
        64'h02f41423_01e45783,
        64'h02f41323_02a00613,
        64'h01c45783_299050ef,
        64'h852285ca_46192a30,
        64'h50ef0064_05132165,
        64'h85930000_a5974619,
        64'h2b5050ef_854e2265,
        64'h85930000_a5974619,
        64'h2c5050ef_854a85ce,
        64'h461900f5_9a230165,
        64'h89930205_89132000,
        64'h0793eaf7_19e32687,
        64'hd7830000_a7970285,
        64'hd703ecf7_11e32764,
        64'h84930000_a49727e7,
        64'hd7830000_a7970265,
        64'hd703b1e1_3e450513,
        64'h00009517_b9c93d65,
        64'h05130000_9517b9f1,
        64'h3b050513_00009517,
        64'hb1dd39a5_05130000,
        64'h9517b9c5_38c50513,
        64'h00009517_b9ed36e5,
        64'h05130000_9517b311,
        64'h36850513_00009517,
        64'hb3393525_05130000,
        64'h9517bb21_34450513,
        64'h00009517_b30d32e5,
        64'h05130000_9517b335,
        64'h32850513_00009517,
        64'hb7993770_50ef0868,
        64'h30058593_0000a597,
        64'h4611f4f7_0de30204,
        64'h5703f6f7_01e317fd,
        64'h67c101e4_5703f6e7,
        64'h87e35fe0_0713bf95,
        64'hcc6ff0ef_02a40513,
        64'h85ca55d0_30ef34e5,
        64'h05130000_9517cdcf,
        64'hf0ef8522_85a65710,
        64'h30ef3525_05130000,
        64'h951702e7_98634d20,
        64'h0713b765_d6dfe0ef,
        64'h02a40513_34458593,
        64'h0000a597_34060613,
        64'h0000a617_34468693,
        64'h0000a697_f7e9439c,
        64'h35078793_0000a797,
        64'hc799439c_36078793,
        64'h0000a797_34f72e23,
        64'h0000a717_47e204e6,
        64'h94630430_07138082,
        64'h616179a2_794274e2,
        64'h640660a6_55c060ef,
        64'h450102a4_0593ff89,
        64'h061b3727_87930000,
        64'ha79766a2_476244b0,
        64'h50efe436_38f72e23,
        64'h0000a717_39c50513,
        64'h0000a517_39458593,
        64'h0000a597_461947e2,
        64'h3ad79e23_0000a797,
        64'h04e79b63_01c15683,
        64'h04500713_00e10e23,
        64'h02344703_00e10ea3,
        64'h01c11903_02244703,
        64'h00e10e23_27810274,
        64'h470300e1_0ea301c1,
        64'h178300f1_0e230254,
        64'h478300f1_0ea30264,
        64'h47030244_4783bdb5,
        64'h43850513_00009517,
        64'hb55942a5_05130000,
        64'h9517bd41_41c50513,
        64'h00009517_a06ddcbf,
        64'he0ef4501_85a202f4,
        64'h12238626_01c15783,
        64'h00a10e23_812100a1,
        64'h0ea3db9f_f0ef00f4,
        64'h1e230029_d78300f4,
        64'h1d230009_d78302f4,
        64'h10230224_0513fde4,
        64'h859b01c4_578300f4,
        64'h1f230204_12230204,
        64'h012301a4_578352b0,
        64'h50ef854a_49c58593,
        64'h0000a597_461953b0,
        64'h50ef8522_85ca4619,
        64'h10f71c63_4ce7d783,
        64'h0000a797_02045703,
        64'h12f71463_4dc98993,
        64'h0000a997_4e47d783,
        64'h0000a797_01e45703,
        64'hb73d61a5_05130000,
        64'h9517f0f5_9ce30880,
        64'h079326f5_89630ff0,
        64'h079326f5_88630890,
        64'h0793b73d_f4f58ae3,
        64'h61050513_00009517,
        64'h06c00793_26f58b63,
        64'h06700793_00b7ef63,
        64'h28f58663_08400793,
        64'hbf91f6f5_8de35fe5,
        64'h05130000_951705e0,
        64'h079328f5_846305c0,
        64'h0793b7bd_f8f58ae3,
        64'h5e850513_00009517,
        64'h03200793_28f58763,
        64'h02f00793_00b7ef63,
        64'h2af58263_03300793,
        64'h04b7e263_2cf58263,
        64'h06200793_b7c95e65,
        64'h05130000_9517faf5,
        64'h96e30290_07932af5,
        64'h86630210_0793bf6d,
        64'hfef580e3_5cc50513,
        64'h00009517_47d916f5,
        64'h8a6347c5_00b7ed63,
        64'h2cf58263_47f5a431,
        64'h7eb030ef_fef591e3,
        64'h5b050513_00009517,
        64'h47a118f5_82634799,
        64'ha41d0040_40ef7465,
        64'h05130000_951702f5,
        64'h83635aa5_05130000,
        64'h95174789_10f58463,
        64'h478502b7_e3631af5,
        64'h83634791_04b7e563,
        64'h1cf58263_47b108b7,
        64'he76332f5_896302e0,
        64'h07930174_458369b0,
        64'h50ef5d25_05130000,
        64'ha5174619_85ca0064,
        64'h09136af0_50ef4611,
        64'h082884b2_05e94407,
        64'h9a638005_079b0af5,
        64'h0e636dd7_879367a1,
        64'h3cf50563_842e8067,
        64'h8793f44e_f84afc26,
        64'he486e0a2_6785715d,
        64'hbf55943e_00e15783,
        64'h00f10723_00d14783,
        64'h00f107a3_34f90909,
        64'h00c14783_701050ef,
        64'h00684609_85ca8082,
        64'h61459141_694264e2,
        64'h1542fff5_45137402,
        64'h70a29522_01045513,
        64'h942a9041_14420104,
        64'h55130290_44634401,
        64'h84ae892a_f406e84a,
        64'hec26f022_71798082,
        64'h62050513_00009517,
        64'hbf7566a5_05130000,
        64'h95178407_8793fce6,
        64'h08e366a5_05130000,
        64'h95178387_8713bfe9,
        64'h65850513_00009517,
        64'h82878793_00c74963,
        64'hfee609e3_67c50513,
        64'h00009517_83078713,
        64'h8082faf6_12e365e5,
        64'h05130000_95178187,
        64'h879300e6_0a6365e5,
        64'h05130000_95178107,
        64'h87138082_01416ce5,
        64'h05130000_a51760a2,
        64'h146040ef_e4066de5,
        64'h05130000_a5176fe5,
        64'h85930000_95979e3d,
        64'h11417c07_879b77fd,
        64'h04c7c963_70c50513,
        64'h00009517_87f78793,
        64'h6785c3ad_68c50513,
        64'h00009517_8006079b,
        64'h04c74963_06e60b63,
        64'h6b050513_00009517,
        64'h80878713_08a74463,
        64'h862a0ce5_07638207,
        64'h87136785_8082953e,
        64'h057e4505_97aa2000,
        64'h0537e308_95360017,
        64'h86930075_6513157d,
        64'h631c77a7_07130000,
        64'ha7178082_40000537,
        64'h8082057e_4505bfb1,
        64'h24050040_60ef854a,
        64'h45818626_20e040ef,
        64'h855e85ca_993e8626,
        64'h8c9d7902_0097ff63,
        64'h77a274c2_99828526,
        64'h0009061b_45c22300,
        64'h40ef856a_86ca85a6,
        64'h66428082_612d6d0a,
        64'h6caa6c4a_6bea7b0a,
        64'h7aaa7a4a_79ea690e,
        64'h64ae644e_60ee5575,
        64'h25a040ef_70450513,
        64'h00009517_85a60397,
        64'he8630184_87b37482,
        64'h04090863_79222780,
        64'h40ef855a_85a2cfbd,
        64'h77c20957_926347a2,
        64'h99829dbd_00280380,
        64'h06137786_028a05bb,
        64'ha0916566_00f46463,
        64'h07815783_764d0d13,
        64'h00009d17_08000cb7,
        64'h80000c37_78cb8b93,
        64'h00009b97_754b0b13,
        64'h00009b17_4a850380,
        64'h0a134401_06e79d63,
        64'h55796318_67470713,
        64'h0000a717_8ff98361,
        64'h577d6786_9982e16a,
        64'he566e962_ed5ef15a,
        64'hf556f952_e1cae5a6,
        64'he9a2ed86_00884581,
        64'h89aa0400_0613fd4e,
        64'h7115bfd5_8f8d2505,
        64'h8082e21c_00b7f463,
        64'h45019181_87aa1582,
        64'hbf390705_01070023,
        64'h0005d463_4185d59b,
        64'h0185959b_c5190975,
        64'h75130005_450300bc,
        64'h05330007_4583bfdd,
        64'h4701bf1d_3cfdfe97,
        64'h6ae32705_67220ee0,
        64'h70efe43a_855eb75d,
        64'h00c58023_0ff67613,
        64'h00ea85b3_0006c603,
        64'hbf6500c5_90239241,
        64'h164295d6_00171593,
        64'h0006d603_006d1c63,
        64'hbfc1e190_95d60037,
        64'h15936290_011d1863,
        64'hbf856862_78820705,
        64'h96d27322_674266a2,
        64'h3aa040ef_e436e83a,
        64'hec42f046_f41a855a,
        64'h65829201_1602c190,
        64'h260195d6_00271593,
        64'h4290030d_1b63b795,
        64'h557dd135_0c2070ef,
        64'h99369281_168241b4,
        64'h043b66a2_3e6040ef,
        64'hfa060c23_e43687e5,
        64'h05130000_a51785d6,
        64'h963e011c_0ac5ed63,
        64'h415705bb_0006861b,
        64'h02e00813_875603bd,
        64'h06bb0d9d_e66399ba,
        64'h03470733_9301020d,
        64'h971305b6_6c630007,
        64'h061b4309_48a14811,
        64'h470186ce_000c8d9b,
        64'h008cf463_00040d9b,
        64'h442040ef_8c450513,
        64'h0000a517_85ca8082,
        64'h616d6daa_6d4a6cea,
        64'h7c0a7baa_7b4a7aea,
        64'h6a0e69ae_694e64ee,
        64'h740e70ae_4501e00d,
        64'h7d8c0c13_00008c17,
        64'h870b8b93_0000ab97,
        64'h908b0b13_0000ab17,
        64'h03810a93_020a5a13,
        64'h0017849b_e03e020d,
        64'h1a13001d_179b03ac,
        64'hdcbb4cc1_000c9563,
        64'h02ccdcbb_04000c93,
        64'h00e7f663_84368d32,
        64'h89ae892a_04000793,
        64'he56ef162_f55ef95a,
        64'hfd56e1d2_eda6f586,
        64'he96ae5ce_e9caf1a2,
        64'h02c7073b_8cbaed66,
        64'h71514e40_406f6105,
        64'h96050513_0000a517,
        64'h64a26902_85a6864a,
        64'h60e26442_4fe040ef,
        64'h95850513_0000a517,
        64'h85a2c801_50e040ef,
        64'h89329625_05130000,
        64'ha5170585_14590087,
        64'hf46300e4_5433942a,
        64'h47a500d4_14334405,
        64'h03b6869b_02f50533,
        64'h47a9c10d_44018d7d,
        64'hfff7c793_00e797b3,
        64'h57fdb7f5_9b450513,
        64'h0000a517_85aafb07,
        64'h9de32785_55e0406f,
        64'h61059ca5_05130000,
        64'ha51785aa_690264a2,
        64'h60e26442_e495e04a,
        64'he822ec06_0007c483,
        64'he42697c2_11019f68,
        64'h08130000_b8179381,
        64'h1782cd85_00e555b3,
        64'h03c6871b_02f886bb,
        64'h481958d9_4781862e,
        64'hb78d9ea5_05130000,
        64'ha51785aa_5b60406f,
        64'h6105a1a5_05130000,
        64'ha5176902_64a285ca,
        64'h862660e2_64425d00,
        64'h40efa2a5_05130000,
        64'ha51785a2_c8015e00,
        64'h40ef84b2_a3450513,
        64'h0000a517_f86102f4,
        64'h5433bfc1_02e45433,
        64'ha039943e_00144413,
        64'h03243413_02e47433,
        64'h02f457b3_06400713,
        64'h02877463_06300713,
        64'hc70502f4_773347a9,
        64'h0287e663_47293e80,
        64'h0793c021_02f555b3,
        64'h02f57433_bf7d2407,
        64'h87934685_b7d9a007,
        64'h87934681_6460406f,
        64'h6105a8a5_05130000,
        64'ha51785aa_690264a2,
        64'h60e26442_02091663,
        64'he426e822_ec060007,
        64'h4903e04a_97361101,
        64'hae870713_0000b717,
        64'h3e800793_46890ca7,
        64'hf7633e70_079304a7,
        64'h676323f7_8713000f,
        64'h47b704a7_6963862e,
        64'h9ff78713_3b9ad7b7,
        64'h8082612d_450160ee,
        64'h6aa040ef_ae450513,
        64'h0000a517_002cfebf,
        64'hf0efed86_45050c80,
        64'h0613002c_7115f73f,
        64'hf06f4581_862e86b2,
        64'h80826145_69a26942,
        64'h64e2854a_740270a2,
        64'h278060ef_afc58593,
        64'h0000a597_00890533,
        64'hffd4841b_00f44463,
        64'hffe4879b_9c296c00,
        64'h40ef954a_b2c60613,
        64'h0000a617_86ce40a4,
        64'h85bb0095_5d630009,
        64'h8f63842a_6de040ef,
        64'h854a85a6_b4460613,
        64'h0000a617_ffc70713,
        64'h00009717_b4c68693,
        64'h0000a697_c50939e6,
        64'h86930000_a6978932,
        64'h89ae84b6_f022f406,
        64'he44ee84a_ec267179,
        64'hbfdd75c0_40ef8562,
        64'hb7e90905_766040ef,
        64'h856600fb_e7630ff7,
        64'hf793fe05_879b0007,
        64'hc583012a_07b3b781,
        64'h04852405_786040ef,
        64'h71850513_0000a517,
        64'h00f45b63_0009079b,
        64'hff047913_79e040ef,
        64'h855aff2d_cce32d85,
        64'h7aa040ef_8556a029,
        64'h00f97913_4d81fffd,
        64'h4913028d_1d637c00,
        64'h40efbd25_05130000,
        64'ha5170104_c583dbe5,
        64'hb7c57d40_40ef8562,
        64'ha0317dc0_40ef8556,
        64'h7e2040ef_77450513,
        64'h0000a517_ffb912e3,
        64'h09057f40_40ef8566,
        64'h02fbe263_0ff7f793,
        64'hfe05879b_0007c583,
        64'h012487b3_4dc14901,
        64'h013040ef_855ae7a9,
        64'hc42900f4_77938082,
        64'h61656da2_6d426ce2,
        64'h7c027ba2_7b427ae2,
        64'h6a0669a6_694664e6,
        64'h740670a6_03344163,
        64'hfff58d1b_c44c8c93,
        64'h0000ac97_c54c0c13,
        64'h0000ac17_06000b93,
        64'hc48b0b13_0000ab17,
        64'h918a8a93_0000ba97,
        64'h4401ff05_049389ae,
        64'h8a2ae46e_e8caf486,
        64'he86aec66_f062f45e,
        64'hf85afc56_e0d2e4ce,
        64'heca6f0a2_7159b7cd,
        64'h093040ef_de07ae23,
        64'h0000b797_c7450513,
        64'h0000a517_80826151,
        64'h641260b2_85220b10,
        64'h40efc5a5_05130000,
        64'ha517c325_85930000,
        64'ha597860a_c10d842a,
        64'hdedff0ef_85220d10,
        64'h40efc525_05130000,
        64'ha517c525_85930000,
        64'ha597842a_00054603,
        64'h00154683_00254703,
        64'h00354783_00454803,
        64'h00554883_e222e606,
        64'h716d8082_7f010113,
        64'h7c813983_7d013903,
        64'h7d813483_7e013403,
        64'h45017e81_30836165,
        64'h8cfff0ef_86c685a6,
        64'h18085632_6882fbaf,
        64'hf0ef03e1_0513863e,
        64'h86c285a2_67c26822,
        64'hf8aff0ef_d64e0521,
        64'h051385a2_864a86ba,
        64'h943e7fc4_04136762,
        64'h747d97ba_81078793,
        64'h10186785_7b8060ef,
        64'hd602e83e_ec3ae442,
        64'h893689b2_e04605a1,
        64'h051384aa_71597d31,
        64'h34237d21_38237c91,
        64'h3c237e81_30237e11,
        64'h34238101_01131990,
        64'h406fd025_05130000,
        64'ha51785aa_80826125,
        64'h7aa27a42_79e26906,
        64'h64a66446_450160e6,
        64'h911a6305_96bff0ef,
        64'h85ce86a6_10084652,
        64'h855ff0ef_460156fd,
        64'h02e10513_85a2821f,
        64'hf0ef0440_06130430,
        64'h06930421_051385a2,
        64'h943e1451_978a020a,
        64'h879312f1_1c233537,
        64'h87936799_12f11b23,
        64'h26378793_77e105b0,
        64'h60ef04f1_06230661,
        64'h05134641_479985ce,
        64'h04f11523_10100793,
        64'h023060ef_ca3e04a1,
        64'h05134581_0f000613,
        64'h0fc00793_089060ef,
        64'h000107a3_15410223,
        64'h14f101a3_14510513,
        64'h460585ca_57fd0a30,
        64'h60ef13f1_05134611,
        64'h95beff04_0593978a,
        64'h020a8793_12f10f23,
        64'h479112f1_0ea30370,
        64'h07930c70_60ef0141,
        64'h07a31a68_460585ca,
        64'h993e978a_020a8793,
        64'h12f11d23_13500793,
        64'hc83e4a05_fef40913,
        64'h439cf027_87930000,
        64'hb7970a50_60ef8526,
        64'h55fd4619_94beff84,
        64'h0493978a_020a8793,
        64'h747d2bd0_40efca02,
        64'h6a85e125_05130000,
        64'ha517911a_89aaf456,
        64'hf852fc4e_e0cae4a6,
        64'he8a2ec86_711d737d,
        64'hb35d2e50_40efdfe5,
        64'h05130000_a517bf45,
        64'hdf850513_0000a517,
        64'h95be978a_d0040593,
        64'h35078793_67853090,
        64'h40efdf25_05130000,
        64'ha5173150_40efdee5,
        64'h05130000_a51700fa,
        64'h20234785_de0796e3,
        64'h000a2783_bbcd3310,
        64'h40efdfa5_05130000,
        64'ha517b501_33f040ef,
        64'hdf050513_0000a517,
        64'h95be978a_f0040593,
        64'h35048793_357040ef,
        64'hdf850513_0000a517,
        64'h95bee004_0593978a,
        64'h35048793_36f040ef,
        64'h02f5d5bb_e107879b,
        64'h678502f6_763b02f5,
        64'hf6bb02f5_d63b03c0,
        64'h079314f7_1e230000,
        64'hb7170121_578316f7,
        64'h13230000_b717e1e5,
        64'h05130000_a51755c2,
        64'h01015783_3af040ef,
        64'he1050513_0000a517,
        64'h01014583_01114603,
        64'h01214683_01314703,
        64'h3cb040ef_e0c50513,
        64'h0000a517_01814583,
        64'h01914603_01a14683,
        64'h01b14703_3e7040ef,
        64'h00b14703_1cf71323,
        64'h0000b717_e0c50513,
        64'h0000a517_00814583,
        64'h35215783_1cf71e23,
        64'h0000b717_00914603,
        64'h00a14683_35015783,
        64'h41b040ef_e0c50513,
        64'h0000a517_35014583,
        64'h35114603_35214683,
        64'h35314703_289060ef,
        64'h01490593_4611953e,
        64'hcb840513_978a3504,
        64'h87936485_2a1060ef,
        64'h0e880109_05934611,
        64'h45b040ef_e3c50513,
        64'h0000a517_00fa2023,
        64'h47851207_9a63000a,
        64'h2783b311_d00d0023,
        64'h2cd060ef_9d228562,
        64'h866ab759_cc048513,
        64'hbb29cef4_2023401c,
        64'h00f40023_ce344783,
        64'h00f400a3_ce244783,
        64'h00f40123_ce144783,
        64'h00f401a3_ce044783,
        64'h305060ef_4611953e,
        64'hce048513_978a3507,
        64'h87936785_bfdd855a,
        64'h4611bbb1_321060ef,
        64'h85564611_b39df00d,
        64'h002332f0_60ef9d22,
        64'h953e866a_f0048513,
        64'h978a3507_87936785,
        64'ha00d953e_978a3507,
        64'h87936785_4611cd04,
        64'h85138082_3b010113,
        64'h35013d03_35813c83,
        64'h36013c03_36813b83,
        64'h37013b03_37813a83,
        64'h38013a03_38813983,
        64'h39013903_39813483,
        64'h3a013403_3a813083,
        64'h911a6305_cebff0ef,
        64'h0e8885de_86ca5672,
        64'hbd5ff0ef_35e10513,
        64'h85a24601_56fdba1f,
        64'hf0ef3721_051385a2,
        64'h04400613_04300693,
        64'h943ecec4_0413978a,
        64'h350a8793_46f11423,
        64'h35378793_679946f1,
        64'h13232637_879377e1,
        64'h3dd060ef_36f10e23,
        64'h39610513_85de4799,
        64'h464136f1_1d231010,
        64'h07933a50_60efde3e,
        64'h37a10513_45810f00,
        64'h06131020_079340b0,
        64'h60ef4731_0d230001,
        64'h03a346f1_0ca347b1,
        64'h051385a6_460557fd,
        64'h425060ef_47410a23,
        64'h47510513_461195be,
        64'hcf440593_978a350a,
        64'h879346f1_09a30360,
        64'h07934470_60ef4741,
        64'h072346f1_05134611,
        64'h4a1195be_cf040593,
        64'h978a350a_879346f1,
        64'h06a30320_079346b0,
        64'h60efc0d2_46c10513,
        64'h85a64605_94becb74,
        64'h0493c2a6_978a350a,
        64'h879346f1_15231350,
        64'h079300f1_03a3478d,
        64'h443060ef_854a55fd,
        64'h4619993e_cf840913,
        64'h978a350a_87936590,
        64'h40efde02_54e25a52,
        64'h02850513_0000a517,
        64'h4bd060ef_953e4611,
        64'h01490593_ce840513,
        64'h978a350a_87934d30,
        64'h60ef013c_a023953e,
        64'h46110109_0593ce44,
        64'h05134985_978a350a,
        64'h87936a85_16079263,
        64'h000ca783_3ae79d63,
        64'h470938e7_81634719,
        64'h24e78163_0007859b,
        64'h747d4715_00614783,
        64'hf8e79ce3_0ff00713,
        64'h24e78563_03800713,
        64'haad94605_cb648513,
        64'hfae798e3_03500713,
        64'h22e78063_03300713,
        64'h00f76e63_22e78363,
        64'h03600713_b759e00d,
        64'h002354f0_60ef9d22,
        64'h953e866a_e0048513,
        64'h978a3507_87936785,
        64'hfee794e3_473d22e7,
        64'h85634731_b77d7210,
        64'h40ef2525_05130000,
        64'ha51785b6_22e78963,
        64'hcc848513_470d2ae7,
        64'h89634705_02f76263,
        64'h24e78163_471904f7,
        64'h6b6326e7_8d630007,
        64'h869b01a9_89bb0589,
        64'h02a00713_29890f07,
        64'hc7830015_cd030139,
        64'h07b395ca_0f098593,
        64'h9c3a9b3a_49818a36,
        64'h8cb28bae_d0048c13,
        64'hcb848b13_970a3507,
        64'h87139aba_cd848a93,
        64'h970a3507_871374fd,
        64'h678526f7_11634789,
        64'h00054703_a0017a90,
        64'h40ef1525_05130000,
        64'ha51785aa_00e7ea63,
        64'h892a5800_073797aa,
        64'hd0040023_f0040023,
        64'he0040023_ca040b23,
        64'hce042023_d00007b7,
        64'h943e747d_978a911a,
        64'h35078793_35a13823,
        64'h35913c23_37813023,
        64'h37713423_37613823,
        64'h37513c23_39413023,
        64'h39313423_38913c23,
        64'h3a113423_39213823,
        64'h3a813023_6785737d,
        64'hc5010113_fadff06f,
        64'h614564e2_00e4859b,
        64'h70a27402_852200f4,
        64'h162347a1_689060ef,
        64'h85b64619_852266a2,
        64'h695060ef_e436f406,
        64'h46190519_84b2842a,
        64'hec26f022_71798082,
        64'h01416402_60a28522,
        64'hfa5ff0ef_e4064501,
        64'h85aa8622_0005841b,
        64'he0221141_bff105a1,
        64'h25050116_b02396ba,
        64'h010686bb_0035169b,
        64'h0005b883_808280c7,
        64'h3823973e_678500f5,
        64'h47636805_450102d7,
        64'hc7bb2785_0077e793,
        64'hfff6079b_8007bc23,
        64'h97ba46a1_67856398,
        64'h53878793_0000b797,
        64'h80826145_740270a2,
        64'h00f41523_fff7c793,
        64'h9fb94107_d71b9fb9,
        64'h93411742_4107579b,
        64'hfed79ce3_9f31ffe7,
        64'hd6030789_470187a2,
        64'h01440693_749060ef,
        64'h01040513_002c4611,
        64'h755060ef_00c40513,
        64'h00041523_006c4611,
        64'h00f404a3_47c576b0,
        64'h60efec3e_00840513,
        64'h00041323_082c4621,
        64'h47c177f0_60ef0044,
        64'h05130161_05934609,
        64'h78d060ef_00f11b23,
        64'hc4360509_084c57fd,
        64'h460900f1_1a238fd9,
        64'h0087979b_0ff77713,
        64'h0087d713_c632842a,
        64'h419c00f5_10230457,
        64'h879b6785_c19c27d1,
        64'hf022f406_7179419c,
        64'h80820005_132300f5,
        64'h122300d5_112300c5,
        64'h10238fd9_0087979b,
        64'h0ff77713_c19c0087,
        64'hd7138ed9_06a20086,
        64'hd71b8e59_27a10622,
        64'h0086571b_419cc19c,
        64'h2785c319_0017f713,
        64'h419cbfcd_fda00513,
        64'h80826121_74a27442,
        64'h70e29782_85a66562,
        64'h701ce509_c39ff0ef,
        64'h842a0830_65a2c105,
        64'hc7dff0ef_84b2e42e,
        64'hf822fc06_f4267139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2655c,
        64'h862686ca_6562e519,
        64'hc75ff0ef_083065a2,
        64'hc115cb7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2615c,
        64'h862686ca_6562e519,
        64'hcb5ff0ef_083065a2,
        64'hc115cf7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hb7e16522_f569cdbf,
        64'hf0ef8526_85ce0030,
        64'hbfc90284_8493c501,
        64'h69f060ef_854a608c,
        64'h292050ef_855285ca,
        64'h60908082_61216a42,
        64'h69e27902_74a27442,
        64'h70e24501_00849b63,
        64'h942602f4_043344ea,
        64'h0a130000_aa1789ae,
        64'h892afc06_e852ec4e,
        64'hf04a0280_079302f4,
        64'h043b840d_8c057a24,
        64'h84930000_b4977aa4,
        64'h04130000_b417f426,
        64'hf822639c_68478793,
        64'h0000b797_7139bfdd,
        64'h45018082_61056442,
        64'h60e2fda0_05138302,
        64'h610560e2_65a26442,
        64'h85220003_0e630205,
        64'h3303c919_db9ff0ef,
        64'he42eec06_4108842a,
        64'he8221101_bfc56562,
        64'hf96dd97f_f0ef0830,
        64'h80826145_70a24501,
        64'he50965a2_de1ff0ef,
        64'hf406e42e_7179bfc1,
        64'h5479fcf7_1be30ff0,
        64'h079300c7_c70367a2,
        64'h0ee080ef_6522f565,
        64'h842adcff_f0ef85a6,
        64'h00308522_80826145,
        64'h64e27402_70a28522,
        64'h543511a0_80ef50e5,
        64'h05130000_a51700f4,
        64'hcf63445c_396050ef,
        64'h51050513_0000a517,
        64'h85a6842a_c11dfda0,
        64'h0413e47f_f0ef84ae,
        64'hf406ec26_f0227179,
        64'h80826145_694264e2,
        64'h740270a2_85221540,
        64'h80ef6522_3ce050ef,
        64'h53850513_0000a517,
        64'h864a608c_ed01842a,
        64'he45ff0ef_84aa85ca,
        64'h0030c11d_fda00413,
        64'he8dff0ef_892eec26,
        64'hf406e84a_f0227179,
        64'hb7d92405_192080ef,
        64'h652240c0_50ef854e,
        64'h85a20127_896300c7,
        64'hc78367a2_ed09e83f,
        64'hf0ef8526_85a20030,
        64'h80826121_69e27902,
        64'h74a27442_70e200f4,
        64'h496344dc_59498993,
        64'h0000a997_0ff00913,
        64'h440184aa_cd01eebf,
        64'hf0efec4e_f04af426,
        64'hf822fc06_7139bfd5,
        64'h54798082_61457402,
        64'h70a28522_1f8080ef,
        64'h00f70963_00c54703,
        64'h0ff00793_6562e911,
        64'h842aee7f_f0ef0830,
        64'h65a2c105_fda00413,
        64'hf2dff0ef_e42ef406,
        64'hf0227179_b7c1fda0,
        64'h0513bf65_24052320,
        64'h80ef4981_65224b00,
        64'h50ef8552_00099563,
        64'h2485cb99_0087c783,
        64'h67a2ed19_f29ff0ef,
        64'h854a85a2_00308082,
        64'h61216a42_69e27902,
        64'h74a27442_70e24501,
        64'hc0915535_00f44d63,
        64'h00c92783_47ca0a13,
        64'h0000ba17_44014481,
        64'h4985892a_cd31f9bf,
        64'hf0efe852_ec4ef04a,
        64'hf426f822_fc067139,
        64'hbfe54501_80820141,
        64'h60a26108_c509fbbf,
        64'hf0efe406_1141b7f5,
        64'h02870713_fea68de3,
        64'h47148082_853a4701,
        64'h00e79563_97ba02d7,
        64'h87b30280_069302d7,
        64'h87bb878d_8f99a1a7,
        64'h87930000_c7976294,
        64'ha2470713_0000c717,
        64'h8f868693_0000c697,
        64'hb7edfda0_07138302,
        64'h853e85b2_00030563,
        64'h01853303_8082853a,
        64'he21c97b6_470102a7,
        64'h87b30a00_051300b7,
        64'hd963454c_0005cc63,
        64'h5735c285_87ae6914,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h000a2e2e_2e746e65,
        64'h6d6f6d20_61207469,
        64'h61772065_7361656c,
        64'h50202165_6e616972,
        64'h41206d6f_7266206f,
        64'h6c6c6548_ffdff06f,
        64'h10500073_34102373,
        64'h342022f3_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_015090ef,
        64'hfec5c6e3_02058593,
        64'h0005bc23_0005b823,
        64'h0005b423_0005b023,
        64'h3b860613_0000c617,
        64'hc2058593_0000c597,
        64'h30579073_09078793,
        64'h00000797_00078067,
        64'h40b787b3_00d787b3,
        64'h01478793_00000797,
        64'hfcc5cce3_02068693,
        64'h02058593_00e6bc23,
        64'h0185b703_00e6b823,
        64'h0105b703_00e6b423,
        64'h0085b703_00e6b023,
        64'h0005b703_0006b703,
        64'hff810113_01b11113,
        64'h0110011b_fe0e9ae3,
        64'h0085b703_fffe8e93,
        64'h0005b703_240e8e9b,
        64'h000f4eb7_01169693,
        64'h3ff6869b_000046b7,
        64'hc0c60613_0000c617,
        64'hfb058593_00000597,
        64'h000280e7_13050513,
        64'h00000517_0b228293,
        64'h00008297_000280e7,
        64'h08c28293_00008297,
        64'h01111113_3ff1011b,
        64'h00004137_fe0e9ee3,
        64'hfffe8e93_710e8e9b,
        64'h00002eb7_11249c63,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
