/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'h011111133ff1011b0000413711249463, /*    1 */
128'h00008297000280e708c2829300008297, /*    2 */
128'h000280e713050513000005170b228293, /*    3 */
128'ha1c606130000c617fc05859300000597, /*    4 */
128'h000f4eb7011696933ff6869b000046b7, /*    5 */
128'h0085b703fffe8e930005b703240e8e9b, /*    6 */
128'hff81011301b111130110011bfe0e9ae3, /*    7 */
128'h0085b70300e6b0230005b7030006b703, /*    8 */
128'h0185b70300e6b8230105b70300e6b423, /*    9 */
128'hfcc5cce3020686930205859300e6bc23, /*   10 */
128'h40b787b300d787b30147879300000797, /*   11 */
128'h30579073090787930000079700078067, /*   12 */
128'h1c8606130000c617a30585930000c597, /*   13 */
128'h0005bc230005b8230005b4230005b023, /*   14 */
128'h020004b7694090effec5c6e302058593, /*   15 */
128'h02000937004484930124a02300100913, /*   16 */
128'h3440297310500073ff24c6e34009091b, /*   17 */
128'hf1402973020004b7fe090ae300897913, /*   18 */
128'h0004a903000920230099093300291913, /*   19 */
128'h4009091b0200093700448493fe091ee3, /*   20 */
128'h1050007334102373342022f3ff24c6e3, /*   21 */
128'h41206d6f7266206f6c6c6548ffdff06f, /*   22 */
128'h617720657361656c502021656e616972, /*   23 */
128'h000a2e2e2e746e656d6f6d2061207469, /*   24 */
128'h00000000000000000000000000000000, /*   25 */
128'h00000000000000000000000000000000, /*   26 */
128'h00000000000000000000000000000000, /*   27 */
128'h00000000000000000000000000000000, /*   28 */
128'h00000000000000000000000000000000, /*   29 */
128'h00000000000000000000000000000000, /*   30 */
128'h00000000000000000000000000000000, /*   31 */
128'hd963454c0005cc635735c28587ae6914, /*   32 */
128'he21c97b6470102a787b30a00051300b7, /*   33 */
128'h853e85b200030563018533038082853a, /*   34 */
128'h6f8686930000b697b7edfda007138302, /*   35 */
128'h87930000c7976294824707130000c717, /*   36 */
128'h87b30280069302d787bb878d8f9981a7, /*   37 */
128'h47148082853a470100e7956397ba02d7, /*   38 */
128'hf0efe4061141b7f502870713fea68de3, /*   39 */
128'hbfe545018082014160a26108c509fbbf, /*   40 */
128'hf0efe852ec4ef04af426f822fc067139, /*   41 */
128'h0000ba17440144814985892acd31f9bf, /*   42 */
128'hc091553500f44d6300c9278327ca0a13, /*   43 */
128'h61216a4269e2790274a2744270e24501, /*   44 */
128'h67a2ed19f29ff0ef854a85a200308082, /*   45 */
128'h50ef8552000995632485cb990087c783, /*   46 */
128'h0513bf652405222080ef498165224a00, /*   47 */
128'hf2dff0efe42ef406f0227179b7c1fda0, /*   48 */
128'h842aee7ff0ef083065a2c105fda00413, /*   49 */
128'h00f7096300c547030ff007936562e911, /*   50 */
128'h547980826145740270a285221e8080ef, /*   51 */
128'hf0efec4ef04af426f822fc067139bfd5, /*   52 */
128'h0000a9970ff00913440184aacd01eebf, /*   53 */
128'h74a2744270e200f4496344dc39498993, /*   54 */
128'hf0ef852685a200308082612169e27902, /*   55 */
128'h85a20127896300c7c78367a2ed09e83f, /*   56 */
128'hb7d92405182080ef65223fc050ef854e, /*   57 */
128'he8dff0ef892eec26f406e84af0227179, /*   58 */
128'he45ff0ef84aa85ca0030c11dfda00413, /*   59 */
128'h338505130000a517864a608ced01842a, /*   60 */
128'h740270a28522144080ef65223be050ef, /*   61 */
128'hf406ec26f022717980826145694264e2, /*   62 */
128'h85a6842ac11dfda00413e47ff0ef84ae, /*   63 */
128'hcf63445c386050ef310505130000a517, /*   64 */
128'h543510a080ef30e505130000a51700f4, /*   65 */
128'h003085228082614564e2740270a28522, /*   66 */
128'h0de080ef6522f565842adcfff0ef85a6, /*   67 */
128'h5479fcf71be30ff0079300c7c70367a2, /*   68 */
128'he50965a2de1ff0eff406e42e7179bfc1, /*   69 */
128'hf96dd97ff0ef08308082614570a24501, /*   70 */
128'he42eec064108842ae8221101bfc56562, /*   71 */
128'h852200030e6302053303c919db9ff0ef, /*   72 */
128'h60e2fda005138302610560e265a26442, /*   73 */
128'h0000b7977139bfdd4501808261056442, /*   74 */
128'h04130000b417f426f822639c48478793, /*   75 */
128'h043b840d8c055a2484930000b4975aa4, /*   76 */
128'h892afc06e852ec4ef04a0280079302f4, /*   77 */
128'h942602f4043324ea0a130000aa1789ae, /*   78 */
128'h69e2790274a2744270e2450100849b63, /*   79 */
128'h282050ef855285ca6090808261216a42, /*   80 */
128'hbfc902848493c50168f060ef854a608c, /*   81 */
128'hb7e16522f569cdbff0ef852685ce0030, /*   82 */
128'h84b68432e42efc06f04af426f8227139, /*   83 */
128'hcb5ff0ef083065a2c115cf7ff0ef893a, /*   84 */
128'h70e2978285a2615c862686ca6562e519, /*   85 */
128'hbfc5fda0051380826121790274a27442, /*   86 */
128'h84b68432e42efc06f04af426f8227139, /*   87 */
128'hc75ff0ef083065a2c115cb7ff0ef893a, /*   88 */
128'h70e2978285a2655c862686ca6562e519, /*   89 */
128'hbfc5fda0051380826121790274a27442, /*   90 */
128'hc7dff0ef84b2e42ef822fc06f4267139, /*   91 */
128'h701ce509c39ff0ef842a083065a2c105, /*   92 */
128'h8082612174a2744270e2978285a66562, /*   93 */
128'h2785c3190017f713419cbfcdfda00513, /*   94 */
128'hd71b8e5927a106220086571b419cc19c, /*   95 */
128'h0ff77713c19c0087d7138ed906a20086, /*   96 */
128'h122300d5112300c510238fd90087979b, /*   97 */
128'hf022f4067179419c80820005132300f5, /*   98 */
128'h419c00f510230457879b6785c19c27d1, /*   99 */
128'h0087979b0ff777130087d713c632842a, /*  100 */
128'hc4360509084c57fd460900f11a238fd9, /*  101 */
128'h051301610593460977d060ef00f11b23, /*  102 */
128'h00041323082c462147c176f060ef0044, /*  103 */
128'h00f404a347c575b060efec3e00840513, /*  104 */
128'h745060ef00c4051300041523006c4611, /*  105 */
128'h01440693739060ef01040513002c4611, /*  106 */
128'hfed79ce39f31ffe7d6030789470187a2, /*  107 */
128'h9fb94107d71b9fb9934117424107579b, /*  108 */
128'h80826145740270a200f41523fff7c793, /*  109 */
128'h97ba46a167856398338787930000b797, /*  110 */
128'hc7bb27850077e793fff6079b8007bc23, /*  111 */
128'h3823973e678500f547636805450102d7, /*  112 */
128'h010686bb0035169b0005b883808280c7, /*  113 */
128'he0221141bff105a125050116b02396ba, /*  114 */
128'hfa5ff0efe406450185aa86220005841b, /*  115 */
128'hec26f022717980820141640260a28522, /*  116 */
128'h685060efe436f4064619051984b2842a, /*  117 */
128'h162347a1679060ef85b64619852266a2, /*  118 */
128'h614564e200e4859b70a27402852200f4, /*  119 */
128'h3a8130236785737dc5010113fadff06f, /*  120 */
128'h3931342338913c233a11342339213823, /*  121 */
128'h377134233761382337513c2339413023, /*  122 */
128'h3507879335a1382335913c2337813023, /*  123 */
128'hce042023d00007b7943e747d978a911a, /*  124 */
128'hd0040023f0040023e0040023ca040b23, /*  125 */
128'ha51785aa00e7ea63892a5800073797aa, /*  126 */
128'h00054703a001799040eff52505130000, /*  127 */
128'h970a3507871374fd678526f711634789, /*  128 */
128'hcb848b13970a350787139abacd848a93, /*  129 */
128'h9c3a9b3a49818a368cb28baed0048c13, /*  130 */
128'hc7830015cd03013907b395ca0f098593, /*  131 */
128'h869b01a989bb058902a0071329890f07, /*  132 */
128'h24e78163471904f76b6326e78d630007, /*  133 */
128'hcc848513470d2ae78963470502f76263, /*  134 */
128'h40ef052505130000a51785b622e78963, /*  135 */
128'hfee794e3473d22e785634731b77d7110, /*  136 */
128'h953e866ae0048513978a350787936785, /*  137 */
128'h03600713b759e00d002353f060ef9d22, /*  138 */
128'h22e780630330071300f76e6322e78363, /*  139 */
128'haad94605cb648513fae798e303500713, /*  140 */
128'hf8e79ce30ff0071324e7856303800713, /*  141 */
128'h24e781630007859b747d471500614783, /*  142 */
128'h000ca7833ae79d63470938e781634719, /*  143 */
128'h05134985978a350a87936a8516079263, /*  144 */
128'h60ef013ca023953e461101090593ce44, /*  145 */
128'h01490593ce840513978a350a87934c30, /*  146 */
128'he28505130000a5174ad060ef953e4611, /*  147 */
128'h978a350a8793649040efde0254e25a52, /*  148 */
128'h433060ef854a55fd4619993ecf840913, /*  149 */
128'h879346f115231350079300f103a3478d, /*  150 */
128'h85a6460594becb740493c2a6978a350a, /*  151 */
128'h06a30320079345b060efc0d246c10513, /*  152 */
128'h4a1195becf040593978a350a879346f1, /*  153 */
128'h0793437060ef4741072346f105134611, /*  154 */
128'hcf440593978a350a879346f109a30360, /*  155 */
128'h415060ef47410a2347510513461195be, /*  156 */
128'h03a346f10ca347b1051385a6460557fd, /*  157 */
128'h0613102007933fb060ef47310d230001, /*  158 */
128'h0793395060efde3e37a1051345810f00, /*  159 */
128'h3961051385de4799464136f11d231010, /*  160 */
128'h13232637879377e13cd060ef36f10e23, /*  161 */
128'h350a879346f1142335378793679946f1, /*  162 */
128'h0440061304300693943ecec40413978a, /*  163 */
128'h85a2460156fdba1ff0ef3721051385a2, /*  164 */
128'h0e8885de86ca5672bd5ff0ef35e10513, /*  165 */
128'h3a0134033a813083911a6305cebff0ef, /*  166 */
128'h38013a03388139833901390339813483, /*  167 */
128'h36013c0336813b8337013b0337813a83, /*  168 */
128'h851380823b01011335013d0335813c83, /*  169 */
128'ha00d953e978a3507879367854611cd04, /*  170 */
128'h953e866af0048513978a350787936785, /*  171 */
128'h85564611b39df00d002331f060ef9d22, /*  172 */
128'h87936785bfdd855a4611bbb1311060ef, /*  173 */
128'h2f5060ef4611953ece048513978a3507, /*  174 */
128'h00f40123ce14478300f401a3ce044783, /*  175 */
128'h00f40023ce34478300f400a3ce244783, /*  176 */
128'h866ab759cc048513bb29cef42023401c, /*  177 */
128'h2783b311d00d00232bd060ef9d228562, /*  178 */
128'h0000a51700fa2023478512079a63000a, /*  179 */
128'h0e8801090593461144b040efc3c50513, /*  180 */
128'hcb840513978a350487936485291060ef, /*  181 */
128'h35314703279060ef014905934611953e, /*  182 */
128'h0000a517350145833511460335214683, /*  183 */
128'h00a146833501578340b040efc0c50513, /*  184 */
128'h35215783fcf71e230000b71700914603, /*  185 */
128'h0000b717c0c505130000a51700814583, /*  186 */
128'h01b147033d7040ef00b14703fcf71323, /*  187 */
128'h0000a517018145830191460301a14683, /*  188 */
128'h01214683013147033bb040efc0c50513, /*  189 */
128'hc10505130000a5170101458301114603, /*  190 */
128'h05130000a51755c20101578339f040ef, /*  191 */
128'hb71701215783f6f713230000b717c1e5, /*  192 */
128'hf6bb02f5d63b03c00793f4f71e230000, /*  193 */
128'h02f5d5bbe107879b678502f6763b02f5, /*  194 */
128'h95bee0040593978a3504879335f040ef, /*  195 */
128'h35048793347040efbf8505130000a517, /*  196 */
128'hbf0505130000a51795be978af0040593, /*  197 */
128'h40efbfa505130000a517b50132f040ef, /*  198 */
128'h20234785de0796e3000a2783bbcd3210, /*  199 */
128'ha517305040efbee505130000a51700fa, /*  200 */
128'h3507879367852f9040efbf2505130000, /*  201 */
128'hbf8505130000a51795be978ad0040593, /*  202 */
128'hb35d2d5040efbfe505130000a517bf45, /*  203 */
128'hf852fc4ee0cae4a6e8a2ec86711d737d, /*  204 */
128'h6a85c12505130000a517911a89aaf456, /*  205 */
128'h0493978a020a8793747d2ad040efca02, /*  206 */
128'hb797095060ef852655fd461994beff84, /*  207 */
128'hc83e4a05fef40913439cd02787930000, /*  208 */
128'h993e978a020a879312f11d2313500793, /*  209 */
128'h07930b7060ef014107a31a68460585ca, /*  210 */
128'h020a879312f10f23479112f10ea30370, /*  211 */
128'h60ef13f10513461195beff040593978a, /*  212 */
128'h14f101a314510513460585ca57fd0930, /*  213 */
128'h0fc00793079060ef000107a315410223, /*  214 */
128'h013060efca3e04a1051345810f000613, /*  215 */
128'h05134641479985ce04f1152310100793, /*  216 */
128'h2637879377e104b060ef04f106230661, /*  217 */
128'h879312f11c2335378793679912f11b23, /*  218 */
128'h06930421051385a2943e1451978a020a, /*  219 */
128'h02e1051385a2821ff0ef044006130430, /*  220 */
128'h85ce86a610084652855ff0ef460156fd, /*  221 */
128'h64a66446450160e6911a630596bff0ef, /*  222 */
128'ha51785aa808261257aa27a4279e26906, /*  223 */
128'h3423810101131890406fb02505130000, /*  224 */
128'h34237d2138237c913c237e8130237e11, /*  225 */
128'h893689b2e04605a1051384aa71597d31, /*  226 */
128'h101867857a8060efd602e83eec3ae442, /*  227 */
128'h943e7fc404136762747d97ba81078793, /*  228 */
128'hf8aff0efd64e0521051385a2864a86ba, /*  229 */
128'hf0ef03e10513863e86c285a267c26822, /*  230 */
128'h8cfff0ef86c685a6180856326882fbaf, /*  231 */
128'h7d8134837e01340345017e8130836165, /*  232 */
128'h716d80827f0101137c8139837d013903, /*  233 */
128'h003547830045480300554883e222e606, /*  234 */
128'ha597842a000546030015468300254703, /*  235 */
128'h40efa52505130000a517a52585930000, /*  236 */
128'ha597860ac10d842adedff0ef85220c10, /*  237 */
128'h40efa5a505130000a517a32585930000, /*  238 */
128'h0000a51780826151641260b285220a10, /*  239 */
128'h083040efbe07ae230000b797a7450513, /*  240 */
128'hf85afc56e0d2e4ceeca6f0a27159b7cd, /*  241 */
128'h8a2ae46ee8caf486e86aec66f062f45e, /*  242 */
128'h718a8a930000aa974401ff05049389ae, /*  243 */
128'h0000ac1706000b93a48b0b130000ab17, /*  244 */
128'hfff58d1ba44c8c930000ac97a54c0c13, /*  245 */
128'h6a0669a6694664e6740670a603344163, /*  246 */
128'h61656da26d426ce27c027ba27b427ae2, /*  247 */
128'h003040ef855ae7a9c42900f477938082, /*  248 */
128'hfe05879b0007c583012487b34dc14901, /*  249 */
128'h09057e4040ef856602fbe2630ff7f793, /*  250 */
128'h7d2040ef574505130000a517ffb912e3, /*  251 */
128'hb7c57c4040ef8562a0317cc040ef8556, /*  252 */
128'h40ef9d2505130000a5170104c583dbe5, /*  253 */
128'h00f979134d81fffd4913028d1d637b00, /*  254 */
128'h855aff2dcce32d8579a040ef8556a029, /*  255 */
128'h00f45b630009079bff04791378e040ef, /*  256 */
128'h04852405776040ef518505130000a517, /*  257 */
128'hf793fe05879b0007c583012a07b3b781, /*  258 */
128'hb7e90905756040ef856600fbe7630ff7, /*  259 */
128'he44ee84aec267179bfdd74c040ef8562, /*  260 */
128'h86930000a697893289ae84b6f022f406, /*  261 */
128'h0000971794c686930000a697c50919e6, /*  262 */
128'h854a85a6944606130000a617dfc70713, /*  263 */
128'h85bb00955d6300098f63842a6ce040ef, /*  264 */
128'h40ef954a92c606130000a61786ce40a4, /*  265 */
128'hffd4841b00f44463ffe4879b9c296b00, /*  266 */
128'h268060ef8fc585930000a59700890533, /*  267 */
128'h8082614569a2694264e2854a740270a2, /*  268 */
128'h0613002c7115f73ff06f4581862e86b2, /*  269 */
128'h0000a517002cfebff0efed8645050c80, /*  270 */
128'h8082612d450160ee69a040ef8e450513, /*  271 */
128'h47b704a76963862e9ff787133b9ad7b7, /*  272 */
128'hf7633e70079304a7676323f78713000f, /*  273 */
128'h8e8707130000b7173e80079346890ca7, /*  274 */
128'he426e822ec0600074903e04a97361101, /*  275 */
128'ha51785aa690264a260e2644202091663, /*  276 */
128'h879346816360406f610588a505130000, /*  277 */
128'h02f57433bf7d240787934685b7d9a007, /*  278 */
128'h0287e66347293e800793c02102f555b3, /*  279 */
128'h0287746306300713c70502f4773347a9, /*  280 */
128'h0324341302e4743302f457b306400713, /*  281 */
128'h5433bfc102e45433a039943e00144413, /*  282 */
128'h40ef84b2834505130000a517f86102f4, /*  283 */
128'h40ef82a505130000a51785a2c8015d00, /*  284 */
128'ha517690264a285ca862660e264425c00, /*  285 */
128'h951785aa5a60406f610581a505130000, /*  286 */
128'h481958d94781862eb78d7ea505130000, /*  287 */
128'h1782cd8500e555b303c6871b02f886bb, /*  288 */
128'he42697c211017f6808130000a8179381, /*  289 */
128'h60e26442e495e04ae822ec060007c483, /*  290 */
128'h61057ca505130000951785aa690264a2, /*  291 */
128'h0000951785aafb079de3278554e0406f, /*  292 */
128'hfff7c79300e797b357fdb7f57b450513, /*  293 */
128'h03b6869b02f5053347a9c10d44018d7d, /*  294 */
128'hf46300e45433942a47a500d414334405, /*  295 */
128'h89327625051300009517058514590087, /*  296 */
128'h758505130000951785a2c8014fe040ef, /*  297 */
128'h64a2690285a6864a60e264424ee040ef, /*  298 */
128'h71514d40406f61057605051300009517, /*  299 */
128'he96ae5cee9caf1a202c7073b8cbaed66, /*  300 */
128'he56ef162f55ef95afd56e1d2eda6f586, /*  301 */
128'h00e7f66384368d3289ae892a04000793, /*  302 */
128'hdcbb4cc1000c956302ccdcbb04000c93, /*  303 */
128'h0017849be03e020d1a13001d179b03ac, /*  304 */
128'h708b0b1300009b1703810a93020a5a13, /*  305 */
128'h5d8c0c1300008c17670b8b9300009b97, /*  306 */
128'h6a0e69ae694e64ee740e70ae4501e00d, /*  307 */
128'h616d6daa6d4a6cea7c0a7baa7b4a7aea, /*  308 */
128'h432040ef6c4505130000951785ca8082, /*  309 */
128'h470186ce000c8d9b008cf46300040d9b, /*  310 */
128'h971305b66c630007061b430948a14811, /*  311 */
128'h06bb0d9de66399ba034707339301020d, /*  312 */
128'h415705bb0006861b02e00813875603bd, /*  313 */
128'h05130000951785d6963e011c0ac5ed63, /*  314 */
128'h043b66a23d6040effa060c23e43667e5, /*  315 */
128'h557dd1350b2070ef99369281168241b4, /*  316 */
128'h260195d6002715934290030d1b63b795, /*  317 */
128'hec42f046f41a855a658292011602c190, /*  318 */
128'h96d27322674266a239a040efe436e83a, /*  319 */
128'h15936290011d1863bf85686278820705, /*  320 */
128'h0006d603006d1c63bfc1e19095d60037, /*  321 */
128'hbf6500c590239241164295d600171593, /*  322 */
128'h00c580230ff6761300ea85b30006c603, /*  323 */
128'h6ae3270567220de070efe43a855eb75d, /*  324 */
128'h053300074583bfdd4701bf1d3cfdfe97, /*  325 */
128'h0185959bc519097575130005450300bc, /*  326 */
128'hbf390705010700230005d4634185d59b, /*  327 */
128'h8082e21c00b7f4634501918187aa1582, /*  328 */
128'h89aa04000613fd4e7115bfd58f8d2505, /*  329 */
128'hf556f952e1cae5a6e9a2ed8600884581, /*  330 */
128'h577d67869982e16ae566e962ed5ef15a, /*  331 */
128'h55796318474707130000a7178ff98361, /*  332 */
128'h00009b174a8503800a13440106e79d63, /*  333 */
128'h80000c3758cb8b9300009b97554b0b13, /*  334 */
128'h07815783564d0d1300009d1708000cb7, /*  335 */
128'h06137786028a05bba091656600f46463, /*  336 */
128'h77c20957926347a299829dbd00280380, /*  337 */
128'h040908637922268040ef855a85a2cfbd, /*  338 */
128'h0000951785a60397e863018487b37482, /*  339 */
128'h64ae644e60ee557524a040ef50450513, /*  340 */
128'h6caa6c4a6bea7b0a7aaa7a4a79ea690e, /*  341 */
128'h40ef856a86ca85a666428082612d6d0a, /*  342 */
128'h77a274c2998285260009061b45c22200, /*  343 */
128'h855e85ca993e86268c9d79020097ff63, /*  344 */
128'h24057f5050ef854a458186261fe040ef, /*  345 */
128'ha7178082400005378082057e4505bfb1, /*  346 */
128'h869300756513157d631c57a707130000, /*  347 */
128'h057e450597aa20000537e30895360017, /*  348 */
128'h862a0ce507638207871367858082953e, /*  349 */
128'h4b050513000095178087871308a74463, /*  350 */
128'h000095178006079b04c7496306e60b63, /*  351 */
128'h0000951787f787936785c3ad48c50513, /*  352 */
128'h11417c07879b77fd04c7c96350c50513, /*  353 */
128'h05130000a5174fe58593000095979e3d, /*  354 */
128'h05130000a51760a2136040efe4064de5, /*  355 */
128'h05130000951781078713808201414ce5, /*  356 */
128'h0513000095178187879300e60a6345e5, /*  357 */
128'h00009517830787138082faf612e345e5, /*  358 */
128'h8287879300c74963fee609e347c50513, /*  359 */
128'h951783878713bfe94585051300009517, /*  360 */
128'h951784078793fce608e346a505130000, /*  361 */
128'h4205051300009517bf7546a505130000, /*  362 */
128'h84ae892af406e84aec26f02271798082, /*  363 */
128'h942a9041144201045513029044634401, /*  364 */
128'h1542fff54513740270a2952201045513, /*  365 */
128'h0068460985ca808261459141694264e2, /*  366 */
128'h00f107a334f9090900c147836f1050ef, /*  367 */
128'hbf55943e00e1578300f1072300d14783, /*  368 */
128'h8793f44ef84afc26e486e0a26785715d, /*  369 */
128'h0e636dd7879367a13cf50563842e8067, /*  370 */
128'h082884b205e944079a638005079b0af5, /*  371 */
128'ha517461985ca0064091369f050ef4611, /*  372 */
128'h07930174458368b050ef3d2505130000, /*  373 */
128'h1cf5826347b108b7e76332f5896302e0, /*  374 */
128'h478502b7e3631af58363479104b7e563, /*  375 */
128'h83633aa5051300009517478910f58463, /*  376 */
128'ha41d7f5030ef546505130000951702f5, /*  377 */
128'h3b0505130000951747a118f582634799, /*  378 */
128'h2cf5826347f5a4317db030effef591e3, /*  379 */
128'h0000951747d916f58a6347c500b7ed63, /*  380 */
128'h866302100793bf6dfef580e33cc50513, /*  381 */
128'h051300009517faf596e3029007932af5, /*  382 */
128'h04b7e2632cf5826306200793b7c93e65, /*  383 */
128'h02f0079300b7ef632af5826303300793, /*  384 */
128'h3e850513000095170320079328f58763, /*  385 */
128'h079328f5846305c00793b7bdf8f58ae3, /*  386 */
128'hbf91f6f58de33fe505130000951705e0, /*  387 */
128'h0670079300b7ef6328f5866308400793, /*  388 */
128'h410505130000951706c0079326f58b63, /*  389 */
128'h079326f5886308900793b73df4f58ae3, /*  390 */
128'h9517f0f59ce30880079326f589630ff0, /*  391 */
128'h0000a79701e45703b73d41a505130000, /*  392 */
128'h12f714632dc989930000a9972e47d783, /*  393 */
128'h10f71c632ce7d7830000a79702045703, /*  394 */
128'h0000a597461952b050ef852285ca4619, /*  395 */
128'h012301a4578351b050ef854a29c58593, /*  396 */
128'h859b01c4578300f41f23020412230204, /*  397 */
128'h1d230009d78302f4102302240513fde4, /*  398 */
128'h0ea3db9ff0ef00f41e230029d78300f4, /*  399 */
128'h1223862601c1578300a10e23812100a1, /*  400 */
128'h00009517a06ddcbfe0ef450185a202f4, /*  401 */
128'hb55922a5051300009517bd4121c50513, /*  402 */
128'h470302444783bdb52385051300009517, /*  403 */
128'h178300f10e230254478300f10ea30264, /*  404 */
128'h00e10e2327810274470300e10ea301c1, /*  405 */
128'h0234470300e10ea301c1190302244703, /*  406 */
128'h04e79b6301c156830450071300e10e23, /*  407 */
128'h0000a597461947e21ad79e230000a797, /*  408 */
128'h0000a71719c505130000a51719458593, /*  409 */
128'ha79766a2476243b050efe43618f72e23, /*  410 */
128'h450102a40593ff89061b172787930000, /*  411 */
128'h616179a2794274e2640660a654c060ef, /*  412 */
128'h0000a71747e204e69463043007138082, /*  413 */
128'hc799439c160787930000a79714f72e23, /*  414 */
128'h0000a697f7e9439c150787930000a797, /*  415 */
128'h0000a597140606130000a61714468693, /*  416 */
128'h0713b765d6dfe0ef02a4051314458593, /*  417 */
128'h30ef152505130000951702e798634d20, /*  418 */
128'h051300009517cdcff0ef852285a65610, /*  419 */
128'hcc6ff0ef02a4051385ca54d030ef14e5, /*  420 */
128'h67c101e45703f6e787e35fe00713bf95, /*  421 */
128'h4611f4f70de302045703f6f701e317fd, /*  422 */
128'hb799367050ef0868100585930000a597, /*  423 */
128'h051300009517b3351285051300009517, /*  424 */
128'h9517bb211445051300009517b30d12e5, /*  425 */
128'h1685051300009517b339152505130000, /*  426 */
128'h00009517b9ed16e5051300009517b311, /*  427 */
128'hb1dd19a5051300009517b9c518c50513, /*  428 */
128'h051300009517b9f11b05051300009517, /*  429 */
128'hd703b1e11e45051300009517b9c91d65, /*  430 */
128'h84930000a49707e7d7830000a7970265, /*  431 */
128'hd7830000a7970285d703ecf711e30764, /*  432 */
128'h89930205891320000793eaf719e30687, /*  433 */
128'h2b5050ef854a85ce461900f59a230165, /*  434 */
128'h2a5050ef854e026585930000a5974619, /*  435 */
128'h50ef00640513016585930000a5974619, /*  436 */
128'h01c45783289050ef852285ca46192930, /*  437 */
128'h02f4142301e4578302f4132302a00613, /*  438 */
128'h00f41f230024d78300f41e230004d783, /*  439 */
128'h0000951785aab36900f4162360800793, /*  440 */
128'h300017b7bba546013fb030ef16c50513, /*  441 */
128'h74132601608130239f0101138307b603, /*  442 */
128'h8406871b0387759366850034171b00f6, /*  443 */
128'h3c23630c8387b783972a300005379f2d, /*  444 */
128'h5f200813ffc5849b2581601134235e91, /*  445 */
128'h00c5963b101005938a1d08b8696335b9, /*  446 */
128'h87930000a797cfb527818ff1fff7c793, /*  447 */
128'h869b7007f7930084179bea254390f4e7, /*  448 */
128'h00d100a3872646d496aa068e9ebd8006, /*  449 */
128'h00d100230086d69b0106d69b0106969b, /*  450 */
128'h806686936685c6918005069b00015503, /*  451 */
128'h67139fad377d8005859b658502d51a63, /*  452 */
128'h868a83f502d7473b1782270546a10077, /*  453 */
128'h862602e6446397c285b6300008378f95, /*  454 */
128'h30838287b823300017b70405aa1ff0ef, /*  455 */
128'h610101135f8134838526600134036081, /*  456 */
128'hbc2306a126050008380300d788338082, /*  457 */
128'he42643c0e8220c2007b71101b7e1ff06, /*  458 */
128'h16938304b703300014b747812401ec06, /*  459 */
128'h0485051300009517e7990206c1630337, /*  460 */
128'h64a2644260e2c3c00c2007b72bf030ef, /*  461 */
128'hf0227179bfc14785eb9ff0ef80826105, /*  462 */
128'he78585930000a597461184ae8432ec26, /*  463 */
128'he30787930000a7970dd050eff4060068, /*  464 */
128'h88930000a89785a6862247b20007a803, /*  465 */
128'ha51704500693e1a757030000a717e168, /*  466 */
128'h740270a285228d4ff0efe22505130000, /*  467 */
128'h15428d5d05220085579b8082614564e2, /*  468 */
128'h8fd966c10185579b0185171b80829141, /*  469 */
128'h0085151b8fd98f750085571bf0068693, /*  470 */
128'h07b7715d808225018d5d8d7900ff0737, /*  471 */
128'h04b005134585460100740207879b0700, /*  472 */
128'hc63eec56f052f44efc26e0a2e486f84a, /*  473 */
128'h30eff825051300009517892a067070ef, /*  474 */
128'h47e1d8078d230000a7970a091a631e10, /*  475 */
128'h0000a71703e00793d8f708a30000a717, /*  476 */
128'h578dd6f70ea30000a7174789d8f70323, /*  477 */
128'h0000a71707f00793d6f70a230000a717, /*  478 */
128'h0048d5c585930000a5974611d6f704a3, /*  479 */
128'h0028d4a585930000a59746097e0050ef, /*  480 */
128'h010006374722f3fff0ef45127d0050ef, /*  481 */
128'h0ff777138ff183210087179bf0060613, /*  482 */
128'h80a6b02317c29101300016b78fd91502, /*  483 */
128'h60a68086b7838006b78380f6b42393c1, /*  484 */
128'h7a0279a2794274e282f6b42347a16406, /*  485 */
128'h4401cea484930000a497808261616ae2, /*  486 */
128'h028a863b4999ec6a0a1300009a175ae1, /*  487 */
128'h00c956330286061b04852405855285a2, /*  488 */
128'hff3410e30f7030effec48fa30ff67613, /*  489 */
128'h71398087b5838007b603300017b7bf91, /*  490 */
128'hf426f822fc068f4d91c115c200800737, /*  491 */
128'h951780e7b423e05ae456e852ec4ef04a, /*  492 */
128'h47030000a7170b9030efe82505130000, /*  493 */
128'h48030000a817c727c7830000a797c797, /*  494 */
128'h46030000a617c606c6830000a697c6b8, /*  495 */
128'h051300009517c4e5c5830000a597c576, /*  496 */
128'h4783c3a404130000a41707d030efe565, /*  497 */
128'h0000a717c14989930000a99744810004, /*  498 */
128'hc08a0a130000aa1700144783c2f70623, /*  499 */
128'h2b3700244783c0f70ba30000a7176a89, /*  500 */
128'h4783c0f702230000a717300019370026, /*  501 */
128'ha71700444783bef70ca30000a7170034, /*  502 */
128'h01a30000a71700544783bef707230000, /*  503 */
128'ha7230000a797ba079d230000a797bef7, /*  504 */
128'ha5230000a797ba07ab230000a797ba07, /*  505 */
128'h0009a783e4a9b807af230000a797ba07, /*  506 */
128'h830937835a0b0493eebfe0ef8522e78d, /*  507 */
128'h03379713830937830207456303379713, /*  508 */
128'h54fd000a2783bfc5bc9ff0effc075de3, /*  509 */
128'hf0efbfc1710a849377d050ef4501dff1, /*  510 */
128'h0005470300154783b7d914fdb7e9baff, /*  511 */
128'h8fd907c200354503002547838f5d07a2, /*  512 */
128'h00f61363367d57fd808225018d5d0562, /*  513 */
128'hb7f5fee50fa3058505050005c7038082, /*  514 */
128'h050500b50023808200f61363367d57fd, /*  515 */
128'h8413e04ae426ec06e8221101495cbfcd, /*  516 */
128'h86ca02000513478101853903cfa50095, /*  517 */
128'h27850006c703462d02e0031348a54815, /*  518 */
128'h011795630e5007130107146300a70e63, /*  519 */
128'h9ee30685040500e40023040500640023, /*  520 */
128'h00f5842384ae01c9051300b94783fcc7, /*  521 */
128'h979b0189470301994783c088f59ff0ef, /*  522 */
128'h016947030179478300f492238fd90087, /*  523 */
128'h60e20004002300f493238fd90087979b, /*  524 */
128'hcf99873e611c80826105690264a26442, /*  525 */
128'h02d5fc630007468303a0061302000593, /*  526 */
128'ha00d577d00d706630017869300c69863, /*  527 */
128'hfd06869b577d46050007c683b7dd0705, /*  528 */
128'he11c0006871b078900b666630ff6f593, /*  529 */
128'hc915bfd5a64747030000a7178082853a, /*  530 */
128'h57030067d683c70d0007c703cb85611c, /*  531 */
128'h60ef0017c503e406114102e690630085, /*  532 */
128'h014160a24525c3914501001577933c40, /*  533 */
128'h468d01a5c70301b5c783808245258082, /*  534 */
128'hc78300d51d630007079b8f5d0087979b, /*  535 */
128'h0107979b8fd50087979b0145c6830155, /*  536 */
128'he44eec26f02271798082853e27818fd9, /*  537 */
128'h4503842a03450993e052e84af4065904, /*  538 */
128'he1312501352060ef85ce862646850015, /*  539 */
128'h00e7eb6340f487bb000402234c58505c, /*  540 */
128'h61456a0269a2694264e2740270a24501, /*  541 */
128'h45034c5cff2a74e34a05003449038082, /*  542 */
128'h397d310060ef85ce86269cbd46850014, /*  543 */
128'hf8dff06fc39900454783b7f94505b7e5, /*  544 */
128'he04ae426ec06e8221101591c80824501, /*  545 */
128'h041bfddff0ef892e84aa02b787634401, /*  546 */
128'h03448593864a46850014c503ec190005, /*  547 */
128'h0324a823597d4405c1192501298060ef, /*  548 */
128'h110180826105690264a2644260e28522, /*  549 */
128'hd91c0005022357fde04ae426ec06e822, /*  550 */
128'h470323344783e52d2501fa3ff0ef842a, /*  551 */
128'h776d0107979b8fd90087979b45092324, /*  552 */
128'h06a4051302f71f63a55707134107d79b, /*  553 */
128'hfff50913010005370005079bd59ff0ef, /*  554 */
128'h8c6345010127f7b31465049300544537, /*  555 */
128'h012575332501d33ff0ef086405130097, /*  556 */
128'h6105690264a2644260e200a035338d05, /*  557 */
128'he0a2e486f44ef84a715dbfcd450d8082, /*  558 */
128'h852e89aa00053023e85aec56f052fc26, /*  559 */
128'h0035171302054e6347addd9ff0ef8932, /*  560 */
128'h47b184aa638097ba868787930000a797, /*  561 */
128'h00144503cb85000447830089b023c015, /*  562 */
128'h891100090563e38d001577931e2060ef, /*  563 */
128'h7a0279a2794274e2640660a647a9c111, /*  564 */
128'h00230ff4f51380826161853e6b426ae2, /*  565 */
128'h478d001577130f4060ef00a400a30004, /*  566 */
128'hf0ef85224581f569891100090463fb71, /*  567 */
128'h0a131fa40913848a04f51a634785ee1f, /*  568 */
128'hf0ef854ac7894501ffc9478389a623a4, /*  569 */
128'hff2a14e30991094100a9a0232501c5bf, /*  570 */
128'h85d6000a876345090004aa8301048913, /*  571 */
128'h470dfe9915e30491c10de9dff0ef8522, /*  572 */
128'hf6e504e34785470db7bd00e519634785, /*  573 */
128'h03f4470304044783bfb947b5c1194a81, /*  574 */
128'h07134107d79b0107979b8fd90087979b, /*  575 */
128'h999b04a4478304b44983fef711e32000, /*  576 */
128'h0444490329811a09866300f9e9b30089, /*  577 */
128'hf793012401a3fff9079b470501342e23, /*  578 */
128'h03e30164012304144b03faf769e30ff7, /*  579 */
128'h04644a03ffc900fb77b3fffb079bfa0b, /*  580 */
128'h0144142300fa6a33008a1a1b04544783, /*  581 */
128'h151b0474448304844503f3c100fa7793, /*  582 */
128'h042447030434478314050e638d450085, /*  583 */
128'h2781033906bbdfb18fd90087979b2501, /*  584 */
128'hf4c564e3873200d7063b9f3d004a571b, /*  585 */
128'h19556905dd8d84ae0364d5bb40c504bb, /*  586 */
128'h490d00b673630905165500b939336641, /*  587 */
128'h2023cc04d458015787bb248900ea873b, /*  588 */
128'h0513f00a15e310e91263470dd05c0354, /*  589 */
128'h1ff4849b0024949bd408b17ff0ef0604, /*  590 */
128'hc45cc81c57fdee99e7e324810094d49b, /*  591 */
128'h478308f91963478d00f402a3f8000793, /*  592 */
128'h0107979b8fd90087979b064447030654, /*  593 */
128'h8522001a859b06f71b6347054107d79b, /*  594 */
128'h2324470323344783e13d2501ce5ff0ef, /*  595 */
128'h776d0107979b8fd90087979b000402a3, /*  596 */
128'h0344051304f71263a55707134107d79b, /*  597 */
128'h1763252787932501416157b7a99ff0ef, /*  598 */
128'h2501614177b7a83ff0ef2184051302f5, /*  599 */
128'ha6dff0ef21c4051300f51c6327278793, /*  600 */
128'h00009797c448a63ff0ef22040513c808, /*  601 */
128'h10230000971793c117c227855ee7d783, /*  602 */
128'h478100042a230124002300f413235ef7, /*  603 */
128'hb5b90005099ba33ff0ef05840513b351, /*  604 */
128'h9fb5e00a05e3b545a25ff0ef05440513, /*  605 */
128'h478db7010014949b00f915634789d41c, /*  606 */
128'h1101bdc59cbd0017d79b8885029787bb, /*  607 */
128'hed692501bffff0ef842ae426ec06e822, /*  608 */
128'h4785005447030cf71063478d00044703, /*  609 */
128'h8526458120000613034404930af71b63, /*  610 */
128'hfaa0079322f4092305500793a01ff0ef, /*  611 */
128'h02f40aa302f40a230520079322f409a3, /*  612 */
128'h0713481c20f40da302f40b2306100793, /*  613 */
128'h571b0107971b20e40d2302e40ba30410, /*  614 */
128'hd71b20e40ea320f40e230087571b0107, /*  615 */
128'h20e40f23445c20f40fa30187d79b0107, /*  616 */
128'h45030087571b0107571b0107971b5010, /*  617 */
128'h260522e400a322f40023072006930014, /*  618 */
128'h20d40ca320d40c230187d79b0107d71b, /*  619 */
128'h50ef85a64685d81022f401a322e40123, /*  620 */
128'h50ef4581460100144503000402a363d0, /*  621 */
128'h610564a2644260e200a0353325016310, /*  622 */
128'h458300f6f96337f9ffe5869b4d1c8082, /*  623 */
128'h8082450180829d2d02d585bb55480025, /*  624 */
128'hf022f406e84a71794d180eb7f7634785, /*  625 */
128'h46890005470302e5f963892ae44eec26, /*  626 */
128'h00f71e6308d70e63468d06d70c63842e, /*  627 */
128'hf0ef9dbd0094d59b9cad515c0015d49b, /*  628 */
128'h694264e2740270a257fdc9112501ac7f, /*  629 */
128'h0014899b0249278380826145853e69a2, /*  630 */
128'hc483854a9dbd94ca1ff4f4930099d59b, /*  631 */
128'h994e1ff9f993f5792501a93ff0ef0344, /*  632 */
128'h8391c0198fc50087979b880503494783, /*  633 */
128'h0085d59b515cbf458fe9157d6505bf65, /*  634 */
128'h74130014141bfd592501a63ff0ef9dbd, /*  635 */
128'h0087979b034945030359478399221fe4, /*  636 */
128'ha39ff0ef9dbd0075d59b515cb7598fc9, /*  637 */
128'h034505131fc575130024151bf9352501, /*  638 */
128'hb76517fd2501100007b7807ff0ef954a, /*  639 */
128'hfc06f04a4540f82271398082853e4785, /*  640 */
128'h892a478500b51523e456e852ec4ef426, /*  641 */
128'h69e2790274a2744270e2450900f41c63, /*  642 */
128'hfee474e34f98611c808261216aa26a42, /*  643 */
128'h579800e69463470d0007c683e02184ae, /*  644 */
128'h008928235788fce4f7e30087d703eb15, /*  645 */
128'h049688bd000937839d3d0044d79bd171, /*  646 */
128'h450100993c2300a92a2394be03478793, /*  647 */
128'h4a8509925a7d843a0027c9838722b75d, /*  648 */
128'h2501e59ff0ef0134f66385a200093503, /*  649 */
128'hfbe301440c630005041be6fff0efbf75, /*  650 */
128'h413484bbf6f476e34f9c00093783f68a, /*  651 */
128'he426e822110100a55583b78d4505bfc1, /*  652 */
128'h484ce4950005049bf33ff0ef842aec06, /*  653 */
128'h06136c08ec990005049b933ff0ef6008, /*  654 */
128'h00e7802357156c1cf3cff0ef45810200, /*  655 */
128'h64a28526644260e200e782234705601c, /*  656 */
128'hf04af426f822fc06e852713980826105, /*  657 */
128'h498984aa4d1c16ba75634a05e456ec4e, /*  658 */
128'h8f63842e89324709000547830af5f063, /*  659 */
128'h0015da1b154794630ee78863470d0ae7, /*  660 */
128'h8b9ff0ef9dbd009a559b00ba0a3b515c, /*  661 */
128'h7793001a0a9b8805060996630005099b, /*  662 */
128'h0347c783014487b3cc191ffa7a130ff9, /*  663 */
128'h8fd98ff50049179b00f7f71316c16685, /*  664 */
128'h00f48223478502fa0a239a260ff7f793, /*  665 */
128'h099b86bff0ef9dbd8526009ad59b50dc, /*  666 */
128'h0049591bc40d1ffafa9300099f630005, /*  667 */
128'h00f482234785032a8a239aa60ff97913, /*  668 */
128'h6aa26a4269e2790274a2854e744270e2, /*  669 */
128'h0089591b0347c783015487b380826121, /*  670 */
128'hd59b515cb7e90127e9339bc100f97913, /*  671 */
128'hfc0992e30005099b811ff0ef9dbd0085, /*  672 */
128'h191b03240a2394261fe474130014141b, /*  673 */
128'h822303240aa30089591b0109591b0109, /*  674 */
128'hfd8ff0ef9dbd0075d59b515cbf790144, /*  675 */
128'h1fc474130024141bf80996e30005099b, /*  676 */
128'h06372501da0ff0ef85569aa603440a93, /*  677 */
128'hd79b94260109179b012569338d71f000, /*  678 */
128'h579b00fa80a30087d79b03240a230107, /*  679 */
128'hb745012a81a300fa81230189591b0109, /*  680 */
128'hf04af822fc06ec4ef4267139bf3d4989, /*  681 */
128'h0a6300c52903e19d89ae84aae456e852, /*  682 */
128'h4c9c5afd4a05844a04f977634d1c0409, /*  683 */
128'hf0efa8214401052a606304f463632405, /*  684 */
128'h1d6357fd0887f86347850005041bc43f, /*  685 */
128'h69e2790274a2744270e28522547d00f4, /*  686 */
128'hfaf47ee3894e4c9c808261216aa26a42, /*  687 */
128'hc05ff0ef852685a24409bf554905b7d5, /*  688 */
128'hfb2411e305450863fd5507e3c9012501, /*  689 */
128'hde9ff0ef852685a2167d10000637b76d, /*  690 */
128'h83e3577dc4c0489c02099063e9052501, /*  691 */
128'h82a30017e7930054c783c89c37fdfae7, /*  692 */
128'h2501dbbff0ef852685ce8622bf4900f4, /*  693 */
128'hf04a7139bfad4405f6f50fe34785dd61, /*  694 */
128'hf426030917932905f822fc0600a55903, /*  695 */
128'h744270e24511eb9993c1e456e852ec4e, /*  696 */
128'h495c808261216aa26a4269e2790274a2, /*  697 */
128'h480c00099d63842a8a2e00f97993d7ed, /*  698 */
128'h0009071b00855783e18dc85c61082785, /*  699 */
128'h03478793012415230996601cfcf775e3, /*  700 */
128'h00495a9b00254783bf5d4501ec1c97ce, /*  701 */
128'h049bb27ff0effc0a9fe30157fab337fd, /*  702 */
128'h946357fdbf4945090097e46347850005, /*  703 */
128'h0ee306f4e0634d1c6008b761450500f4, /*  704 */
128'hd4bd451d0005049be81ff0ef480cf60a, /*  705 */
128'hf0ef6008fcf48de357fdfcf48be34785, /*  706 */
128'h05134581200006136008f5792501dd8f, /*  707 */
128'hf0ef855285a600043a03beeff0ef0345, /*  708 */
128'hed630025478360084a0502aa2823aa5f, /*  709 */
128'h85a6c8046008d91c415787bb591c00fa, /*  710 */
128'hd1cff0ef01450223b7b9c848a83ff0ef, /*  711 */
128'hb7e9db1c27855b1c2a856018f1412501, /*  712 */
128'he456e852ec4ef04afc06f426f8227139, /*  713 */
128'h8663842e84aa02f007130005c783e05a, /*  714 */
128'h0004a62304050ce7906305c0071300e7, /*  715 */
128'h0a9302f00a130ae7fc6347fd00044703, /*  716 */
128'h0d478263000447834b2102e0099305c0, /*  717 */
128'h854a02000593462d0204b9030d578063, /*  718 */
128'h013900230d37926300044783b40ff0ef, /*  719 */
128'h00f900a302e007930b37906300144783, /*  720 */
128'h943a09479763470d1b378e6300244783, /*  721 */
128'hadbff0ef8526458100f905a302000793, /*  722 */
128'h2501cdaff0ef608848cc100510632501, /*  723 */
128'h8ba100b74783c7e5000747836c98e96d, /*  724 */
128'h078507050cb78d6300b78593709cef91, /*  725 */
128'h85264581fed608e3fff7c683fff74603, /*  726 */
128'h4581b791c55c4bdc611cbf75dfdff0ef, /*  727 */
128'h744270e20004bc232501a85ff0ef8526, /*  728 */
128'h808261216b026aa26a4269e2790274a2, /*  729 */
128'h02000693f7578be3bf954709bf1d0405, /*  730 */
128'h47014681b7ad02400793943a12f6e063, /*  731 */
128'ha8dd0505a0d1486502000313478145a1, /*  732 */
128'h00e50023954a9101020695130027e793, /*  733 */
128'h0e50069300094503c6ed4711a06d2685, /*  734 */
128'h979b0165966300d90023469500d51563, /*  735 */
128'h00b6946345850037f6930ff7f7930027, /*  736 */
128'h0087671300d7946346918bb101076713, /*  737 */
128'hbf654701bdfd00e905a3943292011602, /*  738 */
128'hf4e518e34711c50500b7c783709c4511, /*  739 */
128'hbc230004a623cb890207f7930047f713, /*  740 */
128'hb73d4515fb0dbf154501e80703e30004, /*  741 */
128'h609cdbe58bc100b5c7836c8cfbf58b91, /*  742 */
128'h05659a63bdb9c4c8af2ff0ef0007c503, /*  743 */
128'h061b873245ad46a10ff7f7930027979b, /*  744 */
128'hf4e374e3000747039722930117020017, /*  745 */
128'h02b6f263fd370ae3f95704e3f94706e3, /*  746 */
128'h0000851700054c634185551b0187151b, /*  747 */
128'hf11710e30008866300054883ed450513, /*  748 */
128'heea87ae30ff57513fbf7051bbd6d4519, /*  749 */
128'he7933701eea866e30ff57513f9f7051b, /*  750 */
128'he84aec26f0227179bdf90ff777130017, /*  751 */
128'h49bd0e500913451184aef406842ae44e, /*  752 */
128'h2501afaff0ef6008a0b1c90de199484c, /*  753 */
128'hf79300b7c783c3210007c7036c1ce129, /*  754 */
128'hb79317e18bfd033780630327026303f7, /*  755 */
128'h694264e2740270a2450100979a630017, /*  756 */
128'h2501c13ff0ef852245818082614569a2, /*  757 */
128'h45811101bfe54511b7cd00042a23d945, /*  758 */
128'he50d250188fff0ef842ae426ec06e822, /*  759 */
128'hed092501a8cff0ef6008484c0e500493, /*  760 */
128'h85224585cb9900978d630007c7836c1c, /*  761 */
128'h451d00f513634791dd792501bcdff0ef, /*  762 */
128'he426e82211018082610564a2644260e2, /*  763 */
128'h484ce49d0005049bfa9ff0ef842aec06, /*  764 */
128'h06136c08e0850005049ba42ff0ef6008, /*  765 */
128'hf0ef462d6c08700c84cff0ef45810200, /*  766 */
128'h8526644260e200e782234705601c82af, /*  767 */
128'h8082450900b7ed6347858082610564a2, /*  768 */
128'h61456a0269a2694264e2740270a24509, /*  769 */
128'he44ee84af406ec26f02271794d1c8082, /*  770 */
128'h4c1c59fd4a05fcf5fde384ae842ae052, /*  771 */
128'h0005091bec8ff0ef852285a600f4fa63, /*  772 */
128'h03390763fb490ce3bf75450100091463, /*  773 */
128'h481cf15d25018afff0ef852285a64601, /*  774 */
128'h0017e79300544783c81c278501378a63, /*  775 */
128'h7139b7594505bf5d0009049b00f402a3, /*  776 */
128'h83eff0eff42ee432e82efc061028ec2a, /*  777 */
128'h8733050ead4787930000979704054263, /*  778 */
128'hc319676200070023c3196622631800a7, /*  779 */
128'h18634785cb114501e39897aa00070023, /*  780 */
128'h70e22501a0eff0ef0828080c460100f6, /*  781 */
128'he122e506f8ca7175bfe5452d80826121, /*  782 */
128'h0d634925e42ee8daecd6f0d2f4cefca6, /*  783 */
128'h1028002c8a7984aa89b2000530231405, /*  784 */
128'h083c65a2140910630005091b9d6ff0ef, /*  785 */
128'he011e11964062501b6dff0efe4be1028, /*  786 */
128'h4791c54dc3e101f9fa1301c9f7934519, /*  787 */
128'h008a6a132501e75ff0ef102800f51663, /*  788 */
128'h046007937aa2cfcd008a77936406e949, /*  789 */
128'h0004072300f40ca300f408a302100713, /*  790 */
128'h00040ba300040b2300e40823000407a3, /*  791 */
128'h00040ea300040e23000405a300e40c23, /*  792 */
128'he0ef85a2000ac50300040fa300040f23, /*  793 */
128'h00040a2300040da300040d234785fc9f, /*  794 */
128'h04098b6300fa82230005099b00040aa3, /*  795 */
128'he9112501e3fff0ef030aab03855685ce, /*  796 */
128'h250183aff0ef0135262385da39fd7522, /*  797 */
128'hf993e3d98bc500b44783a895892ac90d, /*  798 */
128'h00b44783f565a0854921f60981e30049, /*  799 */
128'h8b85000984630029f993e72d0107f713, /*  800 */
128'h85a279a2020a6a13c399008a7793e3ad, /*  801 */
128'h000485a3d09c01448523f4800309a783, /*  802 */
128'he0ef01c40513c8c8f33fe0ef0009c503, /*  803 */
128'h0004ae230004a623c8880069d783dbbf, /*  804 */
128'h74e6854a640a60aa00f494230134b023, /*  805 */
128'h4911808261496b466ae67a0679a67946, /*  806 */
128'he4d6e8d2eccef8a27119b7d5491db7e5, /*  807 */
128'hf06af466f862fc5ee0daf0caf4a6fc86, /*  808 */
128'he0ef8ab6e4328a2e842a0006a023ec6e, /*  809 */
128'h662200b44783000998630005099be91f, /*  810 */
128'h790674a6854e744670e60007899bc39d, /*  811 */
128'h7d027ca27c427be26b066aa66a4669e6, /*  812 */
128'h160789638b8500a44783808261096de2, /*  813 */
128'h00f67463893e40f907bb445c01042903, /*  814 */
128'h0ce35c7d03040b1320000b930006091b, /*  815 */
128'h5c9b6008120790631ff777934458fa09, /*  816 */
128'h0ffcfc930197fcb337fd002547830097, /*  817 */
128'h478900a7ec6347854848eb11020c9963, /*  818 */
128'h2501bd6ff0ef4c0cb741498900f405a3, /*  819 */
128'hb7a5498500f405a3478501851763b7e5, /*  820 */
128'h2501b98ff0ef856e4c0c00043d83cc08, /*  821 */
128'h849b00a6073b0099579b000c861bd579, /*  822 */
128'h00f6f4639fb1002dc683c4b58d3a0007, /*  823 */
128'h50ef85d2863a86a6001dc503419684bb, /*  824 */
128'hc3850407f79300a44783f94d250114a0, /*  825 */
128'h15020097951b0097fc6341a507bb4c48, /*  826 */
128'h949bc5ffe0ef955285da200006139101, /*  827 */
128'h4099093b445c9a3e9381020497930094, /*  828 */
128'hb70500faa0239fa5000aa783c45c9fa5, /*  829 */
128'hc38d0407f79300a4478304e601634c50, /*  830 */
128'h2501110050efe43a85da4685001dc503, /*  831 */
128'h00f40523fbf7f793672200a44783f139, /*  832 */
128'h0bc050ef85da0017c503863a4685601c, /*  833 */
128'hf5930009049b444c01a42e23f1152501, /*  834 */
128'h85930007849b0127f46340bb87bb1ff5, /*  835 */
128'h499dbf9dbd1fe0ef855295a286260305, /*  836 */
128'hf486fc56e0d2e4cee8caf0a27159b59d, /*  837 */
128'ha023e46ee86aec66f062f45ef85aeca6, /*  838 */
128'h099bcb5fe0ef8ab689328a2e842a0006, /*  839 */
128'h0007899bc39d00b44783000997630005, /*  840 */
128'h7ae26a0669a6694664e6854e740670a6, /*  841 */
128'h808261656da26d426ce27c027ba27b42, /*  842 */
128'h0127873b445c18078f638b8900a44783, /*  843 */
128'h44585c7d03040b1320000b9304f76c63, /*  844 */
128'h5c9b6008140793631ff7779304090463, /*  845 */
128'h0ffcfc930197fcb337fd002547830097, /*  846 */
128'h98634705cb914581485cef01040c9a63, /*  847 */
128'hf0ef4c0cb759498900f405a3478902e7, /*  848 */
128'h12f76a634818445cf3fd0005079bd86f, /*  849 */
128'h9763b79500f405230207e79300a44783, /*  850 */
128'hcc1c4858bf99498500f405a347850187, /*  851 */
128'h601cc38d0407f79300a44783c85ce311, /*  852 */
128'h25017b1040ef85da0017c50346854c50, /*  853 */
128'h3d8300f40523fbf7f79300a44783f969, /*  854 */
128'h869bd159250197cff0ef856e4c0c0004, /*  855 */
128'h8d320007849b00a6863b0099579b000c, /*  856 */
128'h419704bb00f774639fb5002dc703c4b5, /*  857 */
128'hf1512501763040ef85d286a6001dc503, /*  858 */
128'h15820097959b0297f26341a587bb4c4c, /*  859 */
128'h4783a4ffe0ef855a95d2200006139181, /*  860 */
128'h97930094949b00f40523fbf7f79300a4, /*  861 */
128'hc45c9fa54099093b445c9a3e93810204, /*  862 */
128'h8e634c5cbdd100faa0239fa5000aa783, /*  863 */
128'h4685001dc50300e7fa63445c481800c7, /*  864 */
128'h444801a42e23fd0925016c7040ef85da, /*  865 */
128'h0127f46340ab87bb1ff575130009049b, /*  866 */
128'he0ef952285d28626030505130007849b, /*  867 */
128'hbf4100f405230407e79300a447839dbf, /*  868 */
128'h842ae406e0221141bd2d499db5f9c81c, /*  869 */
128'h0207f71300a44783e1752501acffe0ef, /*  870 */
128'hc50346854c50601cc3950407f793cf69, /*  871 */
128'h4783ed552501685040ef030405930017, /*  872 */
128'he0ef6008500c00f40523fbf7f79300a4, /*  873 */
128'h0207671300b7c703741ce15d2501b77f, /*  874 */
128'hd69b0106d69b0107169b481800e785a3, /*  875 */
128'h571b0107569b00d78ea300e78e230086, /*  876 */
128'h00078b23485800e78fa300d78f230187, /*  877 */
128'h0107571b0107169b00e78d2300078ba3, /*  878 */
128'h571b0107571b0107171b00e78a232701, /*  879 */
128'h8c23021007130106d69b00e78aa30087, /*  880 */
128'h8ca300d78da3046007130086d69b00e7, /*  881 */
128'h600800a44783000789a30007892300e7, /*  882 */
128'h640200f50223478500f40523fdf7f793, /*  883 */
128'h0141640260a24505ebbfe06f014160a2, /*  884 */
128'h2501effff0ef842ae406e02211418082, /*  885 */
128'h00043023e11925019cbfe0ef8522e901, /*  886 */
128'hec060028e42a110180820141640260a2, /*  887 */
128'h40a780230000879700054a6395bfe0ef, /*  888 */
128'he42a7159bfe5452d8082610560e24501, /*  889 */
128'hb3bfe0efeca6f486f0a21028002c4601, /*  890 */
128'hf0efe4be1028083c65a2ec190005041b, /*  891 */
128'h575277a2e9916586e41d0005041bcd2f, /*  892 */
128'hc7838082616564e6740670a68522cbd8, /*  893 */
128'h97bfe0ef0004c50374a2cb998bc100b5, /*  894 */
128'h7175bfd94415fcf41ee34791b7c5c8c8, /*  895 */
128'h0023f0d2f4cef8cae122e506e42afca6, /*  896 */
128'h2501acdfe0ef1828002c460184ae0005, /*  897 */
128'h09934bdc597d842677e2ecbe081ce529, /*  898 */
128'he50567a24501040a12634a16c2be02f0, /*  899 */
128'h00e780230307071b3487470300008717, /*  900 */
128'h02f007130e94186300e780a303a00713, /*  901 */
128'h74e6640a60aa00078023078d00e78123, /*  902 */
128'he0ef18284585808261497a0679a67946, /*  903 */
128'h2501e6eff0ef18284581fd452501f89f, /*  904 */
128'hc2aa8cdfe0ef0007c50365c677e2f555, /*  905 */
128'h18284581f9492501f63fe0ef18284581, /*  906 */
128'h0007c50365c677e2e1052501e48ff0ef, /*  907 */
128'hf0ef1828458101450e6325018a7fe0ef, /*  908 */
128'h4509f8e516e367a24711dd612501a9ef, /*  909 */
128'h020797134781f5cfe0ef1828100cb759, /*  910 */
128'h0037871beb05fc974703973610949301, /*  911 */
128'h00e586bb40f405bbfff7871b04e46263, /*  912 */
128'hc79301271a6396b2920166a202069613, /*  913 */
128'h1613b7c12785b7319c3d01368023fff7, /*  914 */
128'h8023377dfc964603962a108892010207, /*  915 */
128'h0204169367220789bddd4545b7e900c6, /*  916 */
128'hfee78fa3240507850007470397369281, /*  917 */
128'hfc06f04af426f8227139b709fe9465e3, /*  918 */
128'h091bfb4fe0ef84ae842ae456e852ec4e, /*  919 */
128'h0007891bcf8900b44783000917630005, /*  920 */
128'h6aa26a4269e2790274a2854a744270e2, /*  921 */
128'h8b8900a4478300977763481880826121, /*  922 */
128'h4818445ce4bd00042623445884bae391, /*  923 */
128'h05230207e79300a44783c81cfcf778e3, /*  924 */
128'h4c50d3e51ff7f793445c4481bf7d00f4, /*  925 */
128'h0407f7930304099300a44783fc960ee3, /*  926 */
128'h30f040ef0017c50385ce4685601cc385, /*  927 */
128'h00f40523fbf7f79300a44783ed512501, /*  928 */
128'h2bd040ef85ce0017c50386264685601c, /*  929 */
128'h999b002547836008bf59cc44ed352501, /*  930 */
128'h563b0336d6bbfff4869b377dc7290097, /*  931 */
128'h27814c0c8ff9413007bb02c6ed630337, /*  932 */
128'h445c0499ea634a855a7dd1c19c9dc45c, /*  933 */
128'hc87fe0ef6008d7b51ff4f793c45c9fa5, /*  934 */
128'he595484cbfb19ca90094d49bcd112501, /*  935 */
128'h478900f5976347850005059b814ff0ef, /*  936 */
128'h478500f5976357fdbded490900f405a3, /*  937 */
128'h4783b765cc0cc84cb5ed490500f405a3, /*  938 */
128'h0005059bfddfe0efcb818b89600800a4, /*  939 */
128'h88e30005059bc4bfe0efbf6984cee599, /*  940 */
128'h445cfaf5fae34f9c601cfabafee3fd45, /*  941 */
128'h7139b7bdc45c013787bb413484bbcc0c, /*  942 */
128'h0828002c4601842ac52de42ef822fc06, /*  943 */
128'he01c852265a267e2e1152501fe6fe0ef, /*  944 */
128'hcd996c0ce529250197cff0eff01c101c, /*  945 */
128'ha02d000430234515e7898bc100b5c783, /*  946 */
128'h458167e2c448e30fe0ef0007c50367e2, /*  947 */
128'h2501cbdfe0ef00f414230067d7838522, /*  948 */
128'h80826121744270e2f971fcf50be34791, /*  949 */
128'he0221141b7c1fcf501e34791bfdd4525, /*  950 */
128'h00043023e1192501dbafe0ef842ae406, /*  951 */
128'he84aec26f022717980820141640260a2, /*  952 */
128'he8890005049bd98fe0ef892e842af406, /*  953 */
128'h0005049bc5ffe0ef8522458100091f63, /*  954 */
128'h30238082614564e269428526740270a2, /*  955 */
128'h136347912501b32ff0ef852245810224, /*  956 */
128'h4581c68fe0ef852285ca00042a2302f5, /*  957 */
128'h2a2300f5166347912501f8bfe0ef8522, /*  958 */
128'he42aeca67159bf6584aad16dbf7d0004, /*  959 */
128'hedafe0eff486f0a21028002c460184ae, /*  960 */
128'hf0efe4be1028083c65a2e00d0005041b, /*  961 */
128'h85a6c489cf816786e8010005041b872f, /*  962 */
128'h616564e6740670a68522c10fe0ef1028, /*  963 */
128'he42af85a8432f0a27159bfcd44198082, /*  964 */
128'he8caeca6f486e0d28522002c46018b2e, /*  965 */
128'h0a1be7cfe0efec66f062f45efc56e4ce, /*  966 */
128'h871b481c01842c836000000a1c630005, /*  967 */
128'h8552740670a600fb202302f76263ffec, /*  968 */
128'h7c027ba27b427ae26a0669a6694664e6, /*  969 */
128'h02fb9f63478500044b83808261656ce2, /*  970 */
128'ha55fe0ef852285ca4a8559fd44814909, /*  971 */
128'h4c1c2485e11109550863093508632501, /*  972 */
128'h0017e793c80400544783fef963e32905, /*  973 */
128'h10000ab7504cb74d009b202300f402a3, /*  974 */
128'h852200099e631afd4c09448149814901, /*  975 */
128'h091385cee9212501d10fe0ef0015899b, /*  976 */
128'h470300194783038b9163200009930344, /*  977 */
128'h39f909092485e3918fd90087979b0009, /*  978 */
128'habcfe0efe02e854ab745fc0c94e33cfd, /*  979 */
128'h39f109112485e1116582015575332501, /*  980 */
128'h1101bfad8a2abfbd4a09b7494a05b7c5, /*  981 */
128'h049bbc4fe0ef842ae04aec06e426e822, /*  982 */
128'h60e20007849bcb9100b44783e4910005, /*  983 */
128'h00a447838082610564a2690285266442, /*  984 */
128'he793fed772e348144458cf390027f713, /*  985 */
128'hf0ef484cef01600800f40523c8180207, /*  986 */
128'h84aa00a405a3c53900042a232501a58f, /*  987 */
128'h146357fd0005091b94dfe0ef4c0cbf7d, /*  988 */
128'he0ef167d100006374c0cb7dd450502f9, /*  989 */
128'h2501a1cff0ef85ca6008f9792501b37f, /*  990 */
128'h6008fcf900e345094785b769449db7e1, /*  991 */
128'hdba50407f79300a44783fcf96ae34d1c, /*  992 */
128'h40ef030405930017c50346854c50601c, /*  993 */
128'h0523fbf7f79300a44783f55d25016ec0, /*  994 */
128'he5061008002c4605e42a7175b7b100f4, /*  995 */
128'h65a2e9052501ca0fe0eff8cafca6e122, /*  996 */
128'h6786e1052501e3bfe0efe0be1008081c, /*  997 */
128'hc59975e2eb890207f79300b7c7834519, /*  998 */
128'h640a60aa451dcb810014f79300b5c483, /*  999 */
128'he0ef00094503790280826149794674e6, /* 1000 */
128'h01492783c89d88c1cc0d0005041bad8f, /* 1001 */
128'h96cfe0ef00a8100c02800613fc878de3, /* 1002 */
128'h4581f1612501951fe0efcaa200a84589, /* 1003 */
128'hfaf518e34791d94d2501836ff0ef00a8, /* 1004 */
128'he0ef7502e411f15525019f5fe0ef1008, /* 1005 */
128'h250191cff0ef85a27502bf612501f20f, /* 1006 */
128'hf1221028002c4605e42a7171b769d575, /* 1007 */
128'hf4def8dafcd6e152e54ee94aed26f506, /* 1008 */
128'h14630005041bbd0fe0efe8eaece6f0e2, /* 1009 */
128'h041bd67fe0efe4be1028083c65a21c04, /* 1010 */
128'h441967a61af4176347911c0409630005, /* 1011 */
128'h4581752218079f630207f79300b7c783, /* 1012 */
128'h44094785180902630005091bb45fe0ef, /* 1013 */
128'he0ef752216f90b63440557fd16f90f63, /* 1014 */
128'h549b85ca7422160414630005041ba98f, /* 1015 */
128'h2000061303440a13f6efe0ef85220109, /* 1016 */
128'h0593462d898fe0ef855200050c1b4581, /* 1017 */
128'h0ff4fb1347c1248188cfe0ef85520200, /* 1018 */
128'h0109d99b02f40fa30104949b0109199b, /* 1019 */
128'h04f4062302e00b930104d49b02100793, /* 1020 */
128'h0084d49b0089d99b046007930ff97a93, /* 1021 */
128'h0404052303740a230200061304f406a3, /* 1022 */
128'h05640423053407a305540723040405a3, /* 1023 */
128'h772280efe0ef0544051385d2049404a3, /* 1024 */
128'h00d6166357d200074603468d05740aa3, /* 1025 */
128'h0107969b06f40723478100f693635714, /* 1026 */
128'hd69b0107979b06f4042327810107d79b, /* 1027 */
128'h07a30087d79b0086d69b0107d79b0106, /* 1028 */
128'h040b99634c8500274b8306f404a306d4, /* 1029 */
128'h47416786e8350005041bf59fe0ef1028, /* 1030 */
128'h071300e78c230210071300e785a37522, /* 1031 */
128'h8d2300e78ca300078ba300078b230460, /* 1032 */
128'h478500978aa301678a2301378da30157, /* 1033 */
128'h7522a82d0005041bd5afe0ef00f50223, /* 1034 */
128'h8dcfe0ef0195022303852823001c0d1b, /* 1035 */
128'h3bfd8552458120000613ec090005041b, /* 1036 */
128'h7522441db7498c6a0ffbfb93f61fd0ef, /* 1037 */
128'h694a64ea740a70aa8522f25fe0ef85ca, /* 1038 */
128'h6d466ce67c067ba67b467ae66a0a69aa, /* 1039 */
128'he42aeca6f0a27159b7c544218082614d, /* 1040 */
128'h9cafe0eff48610284605002c843284ae, /* 1041 */
128'hb65fe0efe4be1028083c65a2e1312501, /* 1042 */
128'h0207f79300b7c783451967a6e9152501, /* 1043 */
128'h8c658cbd752200b74783c30d6706e39d, /* 1044 */
128'h00f502234785008705a38c3d02747413, /* 1045 */
128'h8082616564e6740670a62501c9efe0ef, /* 1046 */
128'hf122f5060088002c4605e02ee42a7171, /* 1047 */
128'h6786120796630005079b964fe0efed26, /* 1048 */
128'h079baf7fe0eff0be083cf4be008865a2, /* 1049 */
128'h7713479900b7c703778610079a630005, /* 1050 */
128'h46550e058e63479165e6100712630207, /* 1051 */
128'h10a8008c02800613e55fd0ef102805ad, /* 1052 */
128'h0c054d6347adf05fd0ef850ae49fd0ef, /* 1053 */
128'h4711cbf90005079baadfe0ef10a86582, /* 1054 */
128'hefc50005079bdc5fe0ef10a80ce79363, /* 1055 */
128'he0dfd0ef00d4851302a10593464d648a, /* 1056 */
128'h478500f485a30207e793640602814783, /* 1057 */
128'h57d64736cbbd8bc100b4c78300f40223, /* 1058 */
128'h059bf2dfd0ef85a60004450306f70863, /* 1059 */
128'hc5a547890005059bcaefe0ef85220005, /* 1060 */
128'h07936706efb10005079bfc3fd0ef8522, /* 1061 */
128'h0107969b57d602f69d630557468302e0, /* 1062 */
128'h979b06f7042327810107d79b06f70723, /* 1063 */
128'hd69b0106d69b0087d79b0107d79b0107, /* 1064 */
128'h00f7022306d707a3478506f704a30086, /* 1065 */
128'he0ef6506e7910005079be24fe0ef0088, /* 1066 */
128'h614d853e64ea740a70aa0005079bb50f, /* 1067 */
128'h4605842ee42ae8a2711dbfcd47a18082, /* 1068 */
128'h65a2e9292501810fe0efec861028002c, /* 1069 */
128'h67a6e12925019abfe0efe4be1028083c, /* 1070 */
128'hcb856786eb950207f79300b7c7834519, /* 1071 */
128'h8ba30087571b00e78b23752200645703, /* 1072 */
128'h8ca30087571b00e78c230044570300e7, /* 1073 */
128'h60e62501ad6fe0ef00f50223478500e7, /* 1074 */
128'h84aee42ae0cae4a6711d808261256446, /* 1075 */
128'hf9bfd0efec86e8a208284601002c8932, /* 1076 */
128'he0efd20208284581c4b9e0510005041b, /* 1077 */
128'h2501b8ffe0ef08284585e5592501ca8f, /* 1078 */
128'h00b48713ca1fd0ef8526462d75c2e93d, /* 1079 */
128'hfff6879bce89000700230200061346ad, /* 1080 */
128'h177d0007c78397a6938117820007869b, /* 1081 */
128'he69fd0ef510c656202090a63fec783e3, /* 1082 */
128'h468304300793470d6562e0150005041b, /* 1083 */
128'h953e034787930270079300e684630005, /* 1084 */
128'h64a6644660e6852200a92023c29fd0ef, /* 1085 */
128'h0004802300f515634791808261256906, /* 1086 */
128'h1028002c4605e42a711db7d5842abf55, /* 1087 */
128'h66a2ec550005041bee3fd0efec86e8a2, /* 1088 */
128'hc78397b6938102061793460100010c23, /* 1089 */
128'hda0210284581ea2902000593eba10007, /* 1090 */
128'he0ef10284585e8410005041bbd6fe0ef, /* 1091 */
128'h462dc3dd650601814783e1792501abbf, /* 1092 */
128'h00e78c23021007136786bc7fd0ef082c, /* 1093 */
128'h00e78ca300078ba300078b2304600713, /* 1094 */
128'h9713fff6079bbf45863eb74d2605a061, /* 1095 */
128'h082cfeb706e300074703973693010207, /* 1096 */
128'h0006c70348b107f00e9343658e2e4781, /* 1097 */
128'h370100a36c6391411542f9f7051b2785, /* 1098 */
128'h00070f1b8ec505130000751793411742, /* 1099 */
128'h6125644660e68522441900eef863a821, /* 1100 */
128'h06080563000548030505bfcdf36d8082, /* 1101 */
128'h078500c6802300fe06b3b7cdffe81be3, /* 1102 */
128'h00f502234785752200f500235795a885, /* 1103 */
128'h02f51b634791b7c10005041b8fefe0ef, /* 1104 */
128'h0005041ba55fe0ef1028dbd501814783, /* 1105 */
128'h6506b07fd0ef4581020006136506f445, /* 1106 */
128'h00e785a347216786ae5fd0ef082c462d, /* 1107 */
128'h068500e58023f91780e3b751842abf19, /* 1108 */
128'h02000613472993811782f4c7e5e30585, /* 1109 */
128'h0e50079301814703f8d771e30007869b, /* 1110 */
128'h230305452e0305052e83bf89eaf71de3, /* 1111 */
128'h8f2ae44ae826ec22110105c528830585, /* 1112 */
128'h00005f97887687f2869a864604050293, /* 1113 */
128'ha38300b647338dfd00c6c5b3464f8f93, /* 1114 */
128'h007585bb0fc1008fa403000f2583000f, /* 1115 */
128'h159b0105883b004f2703ff4fa3839db9, /* 1116 */
128'h05bb0077073b0105e8330198581b0078, /* 1117 */
128'h008f23838e358e6d00f6c6339f3100f8, /* 1118 */
128'h008383bb8e590146561b00c6171b9e39, /* 1119 */
128'h24038ef900b7c6b300d383bb00c5873b, /* 1120 */
128'h0116969b00f6d39b007686bb8ebd00cf, /* 1121 */
128'h061b00d703bbffcfa4039fa100d3e6b3, /* 1122 */
128'h579b9f3d8f2d9fa1007777338f2d0007, /* 1123 */
128'h869b0005881b0f418f5d0167171b00a7, /* 1124 */
128'h859300005597f45f17e300e387bb0003, /* 1125 */
128'h8293000052973def8f9300005f974a65, /* 1126 */
128'haf0301e6c73300cf7f3300d7cf334a62, /* 1127 */
128'hc70300ef0f3b0025c4030015c383000f, /* 1128 */
128'h942a040a4318972a070a93aa038a0005, /* 1129 */
128'h00581f1b010f083b004fa70300ef0f3b, /* 1130 */
128'h0f3b010f68330003a70301b8581b9e39, /* 1131 */
128'ha7039e398e3d8e7501e7c6339f3100f8, /* 1132 */
128'he63340189eb90176561b0096139b008f, /* 1133 */
128'h8efd007f46b305919f3500cf03bb00c3, /* 1134 */
128'hffcfa7039eb90fc101e6c6b3fff5c483, /* 1135 */
128'h40980126d69b9fb900e6941b94aa048a, /* 1136 */
128'h01e777330083c7339fb900d3843b8ec1, /* 1137 */
128'h8f5d0147171b00c7579b9f3d00774733, /* 1138 */
128'h00e407bb0004069b0003861b000f081b, /* 1139 */
128'h53978ffa3bcf0f1300005f17f25599e3, /* 1140 */
128'hc2b30003a703010fc403332383930000, /* 1141 */
128'hc4839f25400000c2c4b3942a040a00d7, /* 1142 */
128'h40809e2194aa048a0043a4039f21011f, /* 1143 */
128'h01c8581b0048171b012fc4830107083b, /* 1144 */
128'h048a00f8073b0083a4039e2101076833, /* 1145 */
128'h129b408000c2863b9ea194aa00e2c2b3, /* 1146 */
128'h03c100c2e6330156561b013fc90300b6, /* 1147 */
128'hc6b300e7c6b3ffc3a4839c3500c702bb, /* 1148 */
128'hd69b9fa50106941b992a9ea1090a0056, /* 1149 */
128'h0007081b00d2843b8ec1000924830106, /* 1150 */
128'h171b0097579b9f3d8f219fa500574733, /* 1151 */
128'h07bb0004069b0002861b0f918f5d0177, /* 1152 */
128'h47132aa2829300005297f5f592e300e4, /* 1153 */
128'h021f43830002a70300d745b38f5dfff6, /* 1154 */
128'h058a93aa038a020f45839f2d022f4403, /* 1155 */
128'h083b0042a5839f2d942a040a418c95aa, /* 1156 */
128'h01a8581b0003a5839e2d0068171b0107, /* 1157 */
128'h8e59fff6c6139db100f8073b01076833, /* 1158 */
128'h0166561b00a6139b0082a5839e2d8e3d, /* 1159 */
128'h44839ead00c703bb00c3e633400c9ead, /* 1160 */
128'ha4038db902c10075e5b3fff7c593023f, /* 1161 */
128'h0115d59b94aa00f5969b048a9db5ffc2, /* 1162 */
128'h47130007081b00b385bb40809fa18dd5, /* 1163 */
128'h00b7579b9f3d007747339fa18f4dfff7, /* 1164 */
128'h0005869b0003861b0f118f5d0157171b, /* 1165 */
128'h07bb010e883b6462f3ef9de300e587bb, /* 1166 */
128'hc97c0505282300c8863b00d306bb00fe, /* 1167 */
128'h715d653c80826105692264c2cd70cd34, /* 1168 */
128'hf052e486e45ee85af44ef84afc26e0a2, /* 1169 */
128'he53c893289ae84aa97b203f7f413ec56, /* 1170 */
128'h00078a1b408b07bb04000b9304000b13, /* 1171 */
128'h020a1a9300090a1b00f9746393811782, /* 1172 */
128'h0144043b86560084853385ce020ada93, /* 1173 */
128'h60bc0174176399d641590933481020ef, /* 1174 */
128'h794274e2640660a6b7c9978244018526, /* 1175 */
128'h653c808261616ba26b426ae27a0279a2, /* 1176 */
128'hf406e44eec26842a03f7f793f0227179, /* 1177 */
128'h00e7802397a2f800071300178513e84a, /* 1178 */
128'h16020006091b40a9863b449d04000993, /* 1179 */
128'h643c0124f5633c9020ef952245819201, /* 1180 */
128'hfd24fde3450197828522603cfc1c078e, /* 1181 */
128'h77978082614569a2694264e2740270a2, /* 1182 */
128'h7797e93c04053423639cf52787930000, /* 1183 */
128'h879300000797ed3c639cf4a787930000, /* 1184 */
128'h850a46410505059311018082e13cb6c7, /* 1185 */
128'h168686930000769747013bf020efec06, /* 1186 */
128'hc78300e107b345413805859300006597, /* 1187 */
128'h46038bbd962e0047d613070506890007, /* 1188 */
128'hfef68fa3fec68f230007c78397ae0006, /* 1189 */
128'h610512a505130000751760e2fca71de3, /* 1190 */
128'hf0efe42ee5060808842ae12271758082, /* 1191 */
128'hf0ef0808e85ff0ef080885a26622f71f, /* 1192 */
128'h80826149640a60aaf83ff0ef0808f01f, /* 1193 */
128'h00d71763469100d70d63711c46a15958, /* 1194 */
128'hbfe50007ac2380824501cf9802000713, /* 1195 */
128'h200007b7ec06e426e82211018082556d, /* 1196 */
128'h058686930000569702f5026384ae842a, /* 1197 */
128'h000065172e4585930000659708800613, /* 1198 */
128'h64a2644260e2fc2419b030ef2f450513, /* 1199 */
128'h07b7ec06e4266100e822110180826105, /* 1200 */
128'h030686930000569702f4026384ae2000, /* 1201 */
128'h000065172a4585930000659702f00613, /* 1202 */
128'h64a2644260e2e00415b030ef2b450513, /* 1203 */
128'h07b7ec06e4266100e822110180826105, /* 1204 */
128'h000686930000569702f4026384ae2000, /* 1205 */
128'h00006517264585930000659703600613, /* 1206 */
128'h64a2644260e2e40411b030ef27450513, /* 1207 */
128'h07b7ec06e8226104e426110180826105, /* 1208 */
128'hea8686930000769702f48263842e2000, /* 1209 */
128'h00006517224585930000659703e00613, /* 1210 */
128'h60e2e880900114020db030ef23450513, /* 1211 */
128'he8226104e42611018082610564a26442, /* 1212 */
128'h0000769702f48263842e200007b7ec06, /* 1213 */
128'h1e0585930000659704500613e5c68693, /* 1214 */
128'h90011402097030ef1f05051300006517, /* 1215 */
128'he82211018082610564a2644260e2ec80, /* 1216 */
128'h02f4026384ae200007b7ec06e4266100, /* 1217 */
128'h0000659704c00613f486869300005697, /* 1218 */
128'h053030ef1ac505130000651719c58593, /* 1219 */
128'he82211018082610564a2644260e2f004, /* 1220 */
128'h02f4026384ae200007b7ec06e4266100, /* 1221 */
128'h0000659705300613f186869300005697, /* 1222 */
128'h013030ef16c505130000651715c58593, /* 1223 */
128'hec4e71398082610564a2644260e2f404, /* 1224 */
128'h200007b7fc06f04af426f82200053983, /* 1225 */
128'h86930000569702f984638436893284ae, /* 1226 */
128'h6517112585930000659705a00613ede6, /* 1227 */
128'h159b67227c6030efe43a122505130000, /* 1228 */
128'h8dd9004979130029191b8b0589890014, /* 1229 */
128'h8dc5744270e288a10125e5b30034949b, /* 1230 */
128'h11418082612169e2790274a202b9b823, /* 1231 */
128'he406458185224605468147057100e022, /* 1232 */
128'h47058522f35ff0ef45818522f7dff0ef, /* 1233 */
128'hf0ef45816008f67ff0ef458146054685, /* 1234 */
128'he4061141808201414501640260a2d97f, /* 1235 */
128'h0405302302053c23460546814705e022, /* 1236 */
128'hef1ff0ef45818522f39ff0ef842a4581, /* 1237 */
128'h6008f23ff0ef46054685470545818522, /* 1238 */
128'he4261101d4dff06f0141458160a26402, /* 1239 */
128'h02f48263842e200007b7ec06e8226104, /* 1240 */
128'h0000659706100613e086869300005697, /* 1241 */
128'h6e2030ef03c505130000651702c58593, /* 1242 */
128'h8082610564a2644260e2fc8090411442, /* 1243 */
128'h842e200007b7ec06e8226104e4261101, /* 1244 */
128'h06800613dd4686930000569702f48263, /* 1245 */
128'hff85051300006517fe85859300006597, /* 1246 */
128'h644260e2e0a08c7d17fd678569e030ef, /* 1247 */
128'hec06e4266100e82211018082610564a2, /* 1248 */
128'h86930000569702f4026384ae200007b7, /* 1249 */
128'h6517fa2585930000659706f00613d9e6, /* 1250 */
128'h644260e2e424658030effb2505130000, /* 1251 */
128'he82200053903e04a11018082610564a2, /* 1252 */
128'h02f9026384ae842a200007b7ec06e426, /* 1253 */
128'h0000659707600613d686869300005697, /* 1254 */
128'h612030eff6c5051300006517f5c58593, /* 1255 */
128'h6105690264a2644260e2c84404993c23, /* 1256 */
128'he4cef486e8caeca67100f0a271598082, /* 1257 */
128'h020408a3ec66f062f45ef85afc56e0d2, /* 1258 */
128'h45814611d01ce03084b2892e0005d783, /* 1259 */
128'h458560080e049c636ca020ef00c90513, /* 1260 */
128'h04043a03200007b700043983bf5ff0ef, /* 1261 */
128'hc7090017f71344810049278316f99a63, /* 1262 */
128'h8cdd03243c234c1c4485e391448d8b89, /* 1263 */
128'he493160786638b85008a2783000a0963, /* 1264 */
128'hd71ff0ef852245814605468147050144, /* 1265 */
128'h5c17852200892583be1ff0ef85224581, /* 1266 */
128'h852200095583c4fff0efce2c0c130000, /* 1267 */
128'h852285a6c81ff0efe88a0a1300006a17, /* 1268 */
128'h46854705cf5ff0ef85224581cbdff0ef, /* 1269 */
128'h8593000f45b7d27ff0ef852245814605, /* 1270 */
128'hcd1ff0ef85224585e93ff0ef85222405, /* 1271 */
128'h25810015e593009899b785220d89b583, /* 1272 */
128'he48a8a9300006a9768198993eb7ff0ef, /* 1273 */
128'h6a0669a6694664e6740670a6efe9485c, /* 1274 */
128'h8082616545016ce27c027ba27b427ae2, /* 1275 */
128'hf0ef8522488cdb7ff0efe024852244cc, /* 1276 */
128'h00043883603cee079be38b85449cdf3f, /* 1277 */
128'h431147014781458163900107e6836541, /* 1278 */
128'h4803ec0689e36e89f005051300ff0e37, /* 1279 */
128'h0107e7b301e8183b070500371f1b0006, /* 1280 */
128'h0187d81bf2e50067036316fd06052781, /* 1281 */
128'h01c878330087981b010767330187971b, /* 1282 */
128'h00be873b8fd98fe9010767330087d79b, /* 1283 */
128'h47812585e31c97469381837517821702, /* 1284 */
128'h14900613b846869300005697b7654701, /* 1285 */
128'hd785051300006517d685859300006597, /* 1286 */
128'h0bb78b4ebd6100c4e493bd8541e030ef, /* 1287 */
128'hb685859300005597000b1d633b7d2000, /* 1288 */
128'h3903b7116f6000efd685051300006517, /* 1289 */
128'h855685d20f20061386e2017909630004, /* 1290 */
128'h24818cfd4c81485c070934833de030ef, /* 1291 */
128'h00f76f630c8937830209370312048e63, /* 1292 */
128'hf0ef85224581cc5cf9200793c7817c1c, /* 1293 */
128'hc3950044f793b27ff0ef85224581b6ff, /* 1294 */
128'h85ca00896913ff397913852201442903, /* 1295 */
128'h00efd0a505130000651785cad47ff0ef, /* 1296 */
128'h7913852201442903c3950084f7936800, /* 1297 */
128'h651785cad1fff0ef85ca00496913ff39, /* 1298 */
128'hcfb50014f793658000efd0a505130000, /* 1299 */
128'h00005697017c8c630384390300043c83, /* 1300 */
128'h332030ef855685d209c00613ad468693, /* 1301 */
128'hf693470d02043c2300492783cba97c1c, /* 1302 */
128'h468100c90793018c871308e69f630037, /* 1303 */
128'hc3900086161bff87051363104591480d, /* 1304 */
128'h2685c3988f518361ff87370301068763, /* 1305 */
128'he793485ccbb5603cfeb690e30791872a, /* 1306 */
128'hcc9d4c858889c85c9bf9485cc85c0027, /* 1307 */
128'h86930000569701748c63040439036004, /* 1308 */
128'h30232b4030ef855685d20ca00613a6e6, /* 1309 */
128'h8522ef8d8b8500892783000909630404, /* 1310 */
128'h8522484cc85c9bf54c85485cb4dff0ef, /* 1311 */
128'hbd95641020ef4505d80c8ee3c47ff0ef, /* 1312 */
128'h8522b77100f92623000cb783dbd98b85, /* 1313 */
128'h3c830109648397a667a1bf41b1dff0ef, /* 1314 */
128'h8566639c00878913fa978de394be0009, /* 1315 */
128'hb7dd87ca0ca139a020efe43e002c4621, /* 1316 */
128'hec26f02204800513717908b041635535, /* 1317 */
128'h842a1a4030ef892e84b2e44ef406e84a, /* 1318 */
128'h10ef9da505130000551785a2cc1d5551, /* 1319 */
128'hbd85051300006517862285aa89aa7850, /* 1320 */
128'h2423e01c200007b702098b634fe000ef, /* 1321 */
128'h4501c45c4789cb990024f793f4040124, /* 1322 */
128'h88858082614569a2694264e2740270a2, /* 1323 */
128'h18c030ef8522b7e5c45c4785d4fd4501, /* 1324 */
128'hf06f20000537458146098082bff9557d, /* 1325 */
128'h808225016108953e050e200007b7f73f, /* 1326 */
128'h0263200007b7e4066380e0221141711c, /* 1327 */
128'h659734c00613976686930000569702f4, /* 1328 */
128'h30efaca5051300006517aba585930000, /* 1329 */
128'h0141640260a2557de3914505703c1700, /* 1330 */
128'h10efe42eec064501842ae82211018082, /* 1331 */
128'h006f6105468560e26622644285a24d30, /* 1332 */
128'he84aec26f022f4062000051371797940, /* 1333 */
128'h05130000651784aa0aa030efe052e44e, /* 1334 */
128'h450144b010ef0001b5031b2030efb2e5, /* 1335 */
128'h00006517681c206010ef842a491010ef, /* 1336 */
128'h651706f445833f8000ef638cb1450513, /* 1337 */
128'h00006517546c3e8000efb12505130000, /* 1338 */
128'h3d2000ef91c115c20085d59bb1c50513, /* 1339 */
128'hd71bb12505130000651706c44583583c, /* 1340 */
128'hf7930ff777130187d61b0107d69b0087, /* 1341 */
128'h65175c0c3a6000ef26010ff6f6930ff7, /* 1342 */
128'h00006597545c398000efb02505130000, /* 1343 */
128'h6517a7a5859300006597c789a8c58593, /* 1344 */
128'h051300006517378000efaf2505130000, /* 1345 */
128'h10058593000065977448102030efafe5, /* 1346 */
128'h061300006617584c19c42783dc9fb0ef, /* 1347 */
128'h00006517db46061300006617e789a566, /* 1348 */
128'hf0ef84264581852633a000efadc50513, /* 1349 */
128'h00006997adca0a1300006a174481ed5f, /* 1350 */
128'h85a6e78901f4f79320000913adc98993, /* 1351 */
128'hf6132485854e0004458330c000ef8552, /* 1352 */
128'h6517fd249fe304052fa000ef819100f5, /* 1353 */
128'h64e2740270a22e8000ef08a505130000, /* 1354 */
128'h0103b7038082614545016a0269a26942, /* 1355 */
128'h1782278540f707b30003b6830083b783, /* 1356 */
128'h002300f3b8230017079300d7fe639381, /* 1357 */
128'h450180820007802345050103b78300a7, /* 1358 */
128'h9201020596130103b7830083b7038082, /* 1359 */
128'h00c6f5638e9dfff706930003b7038f99, /* 1360 */
128'h0103b70340a786bb87aa9d9dfff7059b, /* 1361 */
128'h001706938082852e0007002300b6e663, /* 1362 */
128'hbfe900d7002307850007c68300d3b823, /* 1363 */
128'h0693488540a0053be681000556634881, /* 1364 */
128'h86ba4e250ff6f81304100693c2190610, /* 1365 */
128'h67630ff3751302b6733b0005061b3859, /* 1366 */
128'h06850ff5751302b6563b0305051b046e, /* 1367 */
128'h0300051340e685bbfe718532fea68fa3, /* 1368 */
128'h00f6802302d007930008876302f5e963, /* 1369 */
128'h2581000680230015559b40e6853b0685, /* 1370 */
128'h00a8053b808200b61b63fff5081b86ba, /* 1371 */
128'h40c807bbb7d92585fea68fa30685bf5d, /* 1372 */
128'h26050006c8830007c30397ba93811782, /* 1373 */
128'hf0ca7119b7f106850117802300668023, /* 1374 */
128'hfc86e4d6e8d2eccef4a6f8a2597d011c, /* 1375 */
128'h0993f82af02ef42afc3e843684b2e0da, /* 1376 */
128'h77420209591303000a9306c00a130250, /* 1377 */
128'h76820017079bc52d8f1d0004c50377a2, /* 1378 */
128'h039304850135086304d7ff6393811782, /* 1379 */
128'h05450f630014c503bfe1e7bff0ef0201, /* 1380 */
128'h879bcb9d0004c7830355106347810489, /* 1381 */
128'hc503478100f6f36346a50ff7f793fd07, /* 1382 */
128'h02a6eb6306d50f630640069304890014, /* 1383 */
128'h08f509630630079304d50f6305800693, /* 1384 */
128'h6aa66a4669e6790674a6744670e6f55d, /* 1385 */
128'h048d0024c503808261090007051b6b06, /* 1386 */
128'h071300a76c6306e50e6307300713b74d, /* 1387 */
128'h46014685003800840b13f6e51ee30700, /* 1388 */
128'h10e30780071302e5006307500713a00d, /* 1389 */
128'h36134685003800840b13fa850613f6e5, /* 1390 */
128'h003800840b13f8b50693a81145c10016, /* 1391 */
128'h059be37ff0ef400845a946010016b693, /* 1392 */
128'h4503a809ddbff0ef0028020103930005, /* 1393 */
128'h845ad93ff0ef00840b13020103930004, /* 1394 */
128'h10ef852201247433600000840b13b5fd, /* 1395 */
128'h715db7f18522020103930005059b4db0, /* 1396 */
128'he436e4c6e0c2fc3ef83aec061034f436, /* 1397 */
128'hf436f032715d8082616160e2e8dff0ef, /* 1398 */
128'he0c2fc3ef83aec06100005931014862e, /* 1399 */
128'h710d8082616160e2e69ff0efe436e4c6, /* 1400 */
128'h0808100005931234862afe36fa32f62e, /* 1401 */
128'hf0efe436eec6eac2e6bee2baea22ee06, /* 1402 */
128'h645260f28522129020ef0808842ae3ff, /* 1403 */
128'h000303630087b303679c691c80826135, /* 1404 */
128'h0205979304b7ee63479d808245018302, /* 1405 */
128'h1101439c97ba83f94d07071300004717, /* 1406 */
128'h08c52483795c878297bae426e822ec06, /* 1407 */
128'h57b39381020497930c5010ef7540f55c, /* 1408 */
128'h808261054501e91c64a2644260e202f4, /* 1409 */
128'h95aa058e05e135f1bfd9617cbfe97d5c, /* 1410 */
128'he02211418082557d8082557db7e9659c, /* 1411 */
128'h679c681c00055e63ff5ff0ef842ae406, /* 1412 */
128'h014160a264028522000307630207b303, /* 1413 */
128'h8082557d80820141640260a245018302, /* 1414 */
128'h4587879300004797150200a7eb6347ad, /* 1415 */
128'h6d8505130000551780826108953e8175, /* 1416 */
128'h47a1715d83020007b303679c691c8082, /* 1417 */
128'he42e078517824785d23e47d502f11023, /* 1418 */
128'hcc3ed402e486100c200007930030e83e, /* 1419 */
128'h400407374d148082616160a6fd3ff0ef, /* 1420 */
128'h34032381308345018082450100e6fe63, /* 1421 */
128'hdc010113808224010113228134832301, /* 1422 */
128'h2291342385a2980101f1041322813823, /* 1423 */
128'hc703f579f95ff0ef1a05348322113c23, /* 1424 */
128'h47830dd4c70302f71c630a0447830a04, /* 1425 */
128'h10630c0447830c04c70302f716630dd4, /* 1426 */
128'h461100f71a630e0447830e04c70302f7, /* 1427 */
128'h0513d55156f010ef0d4485130d440593, /* 1428 */
128'hf4063e800513842af0227179b761fb60, /* 1429 */
128'hc40200011023858a460185226ea020ef, /* 1430 */
128'h20ef7d000513e509842af21ff0efc202, /* 1431 */
128'h4785717980826145740270a285226cc0, /* 1432 */
128'h842ac402c23ef406f022478500f11023, /* 1433 */
128'hf80787934ad4008007b745386914c195, /* 1434 */
128'h8f55400006b78f75600006b78ff58ff9, /* 1435 */
128'he119ec9ff0ef8522858a4601c43e8fd9, /* 1436 */
128'h47b5711d80826145740270a2c43c47b2, /* 1437 */
128'hfc4ee0ca07c55783c23e47d500f11023, /* 1438 */
128'he8a26a056989fdf949370107979bf852, /* 1439 */
128'h09134495c43e842e8aaaec86f456e4a6, /* 1440 */
128'h8556858a4601e00a0a13e00989930809, /* 1441 */
128'hf7b3c7891005f79345b2ed0de73ff0ef, /* 1442 */
128'h00005517c78d0125f7b3054793630135, /* 1443 */
128'h644660e6fba00513d4bff0ef53450513, /* 1444 */
128'h34fd808261257aa27a4279e2690664a6, /* 1445 */
128'h051300f057630014079b347dfe04c6e3, /* 1446 */
128'h5517fc8049e34501b7555d8020ef3e80, /* 1447 */
128'hbf7df9200513d09ff0ef50a505130000, /* 1448 */
128'hc42e00f1102347c17139e7a919c52783, /* 1449 */
128'hc23e842af426fc06f822858a460147d5, /* 1450 */
128'h4495cb918b891b842783c11dde3ff0ef, /* 1451 */
128'hf8ed34fdc901dcdff0ef8522858a4601, /* 1452 */
128'h4501bfd545018082612174a2744270e2, /* 1453 */
128'h892a4785e8a2ec86e0cae4a6711d8082, /* 1454 */
128'h02f1102302c9270347c906d7f66384b6, /* 1455 */
128'hcc3ee42e4755d432cf3108c927832601, /* 1456 */
128'hf0efc83eca26d23a854a100c47850030, /* 1457 */
128'h102347b10497f0634785e529842ad75f, /* 1458 */
128'hf0efd23ed402854a100c47f5460102f1, /* 1459 */
128'hc43ff0ef4645051300005517c11dd55f, /* 1460 */
128'h47c580826125690664a6644660e68522, /* 1461 */
128'h4401b7d50004841bb74d02f6063bbf61, /* 1462 */
128'he852ec4ef04af426f822fc067139b7c5, /* 1463 */
128'h10ef8ab684b28a2e4148842ace05e456, /* 1464 */
128'h8d9fa0ef852200b44583c11d892a4820, /* 1465 */
128'h551700b67a63014485b3681000054d63, /* 1466 */
128'h2583a0894481bd9ff0ef41a505130000, /* 1467 */
128'h0109378389a6f96decdff0ef854a08c9, /* 1468 */
128'h85d6865286a2844e0089f3630207e403, /* 1469 */
128'h89b308c96783fc851ae3f01ff0ef854a, /* 1470 */
128'h70e2fc0999e39aa2028784339a224089, /* 1471 */
128'h61216aa26a4269e274a2790285267442, /* 1472 */
128'h969bc23e47f500f11023479971398082, /* 1473 */
128'hf8228ed10106161b8edd030007b70086, /* 1474 */
128'h8526858a4601440dc43684aafc06f426, /* 1475 */
128'hd91ff0ef85263e800593e919c53ff0ef, /* 1476 */
128'hbfcdfc79347d8082612174a2744270e2, /* 1477 */
128'h9fb923213823bffc07b7db0101134d18, /* 1478 */
128'h2331342322913c232481302324113423, /* 1479 */
128'h980101f104131ce7f56349013ffc0737, /* 1480 */
128'hb7831e051863892ac09ff0ef84aa85a2, /* 1481 */
128'h1aa4b023766020ef20000513e7991a04, /* 1482 */
128'h10ef85a2200006131e0503631a04b503, /* 1483 */
128'h000047171cf76b6347210c0447831230, /* 1484 */
128'h8793400407b753b897ba078a00470713, /* 1485 */
128'h071367050d44278300e7fd63cc981ff7, /* 1486 */
128'h4783f8dc00d773630147d69307a68007, /* 1487 */
128'h0019f9938b8506f48f2309b449830a04, /* 1488 */
128'h08f480a30b344783c7890e244783e781, /* 1489 */
128'h09c44783c7898b890a04478300098a63, /* 1490 */
128'h0c848613091407130e24478306f48fa3, /* 1491 */
128'h07c6468109d405130a844783fcdc07c6, /* 1492 */
128'h959b0087979b00074583fff74783e0fc, /* 1493 */
128'h8c634685c39197aeffe745839fad0105, /* 1494 */
128'h87b30dd4478302f585b30e0445830009, /* 1495 */
128'h8f63fca714e30621070de21c07ce02b7, /* 1496 */
128'h0107979b468508d4470308e447830409, /* 1497 */
128'h0e04470397ba08c447039fb90087171b, /* 1498 */
128'hf8fc07ce02e787b30dd4478302f70733, /* 1499 */
128'h0107171b0187979b08a4470308b44783, /* 1500 */
128'h088447039fb90087171b089447039fb9, /* 1501 */
128'h0a044783f4fc07a6c319f4fc54d89fb9, /* 1502 */
128'h4685ce81e3918bfd09c44783c7898b85, /* 1503 */
128'h4785ed35e0bff0ef852645850af00613, /* 1504 */
128'hc7b98b850e0446830af447830af407a3, /* 1505 */
128'h00098663c79954dc08f4aa2300a6979b, /* 1506 */
128'h00a6969b0dd44783f8dc07a60d442783, /* 1507 */
128'h08f480230a74478308d4ac2302f686bb, /* 1508 */
128'h390323813483854a2401340324813083, /* 1509 */
128'hd71b50fc808225010113228139832301, /* 1510 */
128'h07bb278527058bfd8b7d0057d79b00a7, /* 1511 */
128'hd1691a04b503892abf4d08f4aa2302f7, /* 1512 */
128'h5929bf555951bf651a04b0235c8020ef, /* 1513 */
128'h34232281382322113c23dc010113bf45, /* 1514 */
128'h02b7e16302f588634789232130232291, /* 1515 */
128'h8526230134032381308354a9c5854681, /* 1516 */
128'h879b8082240101132281348322013903, /* 1517 */
128'h0b900613842e4685fef760e34705ffc5, /* 1518 */
128'hffe4059bf57184aad1fff0ef892a4585, /* 1519 */
128'h854a85a2980101f10413f1e9258199f5, /* 1520 */
128'hdf400493f7d50b944783e51998dff0ef, /* 1521 */
128'hf406e44ee84aec267179b74d84aab75d, /* 1522 */
128'h9be10079f6930ff5f99308154783f022, /* 1523 */
128'hcc7ff0ef84aa45850b3006138edd892e, /* 1524 */
128'h85ca00091c6300f51e63842a57b5c519, /* 1525 */
128'h05a315e010ef8526842a875ff0ef8526, /* 1526 */
128'h614569a2694264e2740270a285220135, /* 1527 */
128'h34232881382328113c23d60101138082, /* 1528 */
128'h34232741382327313c23292130232891, /* 1529 */
128'h34232581382325713c23276130232751, /* 1530 */
128'h0ac7e963478923b13c2325a130232591, /* 1531 */
128'h3ffc07b79f3dbff7879bbffc07b74d18, /* 1532 */
128'h05130000551784ae8b32892abfe78793, /* 1533 */
128'he7b90016779307e9460300e7eb6301e5, /* 1534 */
128'hf8400413f96ff0ef0405051300005517, /* 1535 */
128'h39032881348329013403298130838522, /* 1536 */
128'h3b0326813a8327013a03278139832801, /* 1537 */
128'h3d0324813c8325013c0325813b832601, /* 1538 */
128'h0989270380822a01011323813d832401, /* 1539 */
128'h81630045aa83db450185051300005517, /* 1540 */
128'h02ecf7bb0005ac83e79102eaf7bb060a, /* 1541 */
128'h5429f24ff0ef01e5051300005517cb89, /* 1542 */
128'h9c9be3994b8502eadabb02c92783bf41, /* 1543 */
128'h4e85478189d6856200c488138c0a009c, /* 1544 */
128'h0d6302e8f33b0017859b000828834e11, /* 1545 */
128'hb7c1ee4ff0ef01650513000055170003, /* 1546 */
128'h0065202302e8d33bb7f14b814a814c81, /* 1547 */
128'hcb898b850107c78397a6078e02088063, /* 1548 */
128'h013309bb0ffbfb9300dbebb300be96bb, /* 1549 */
128'h8a09000b8963fbc596e387ae05110821, /* 1550 */
128'h02f10a13f00600e3ff85051300005517, /* 1551 */
128'h19e3842af94ff0ef854a85d2fe0a7a13, /* 1552 */
128'h979b0106161b09ea478309fa4603ee05, /* 1553 */
128'h85ce01367a63963e09da47839e3d0087, /* 1554 */
128'hc783b5c1e56ff0effe85051300005517, /* 1555 */
128'h8b89c71989b60017f7130a7a46830084, /* 1556 */
128'h4611450547010016e993c3990fe6f993, /* 1557 */
128'h78130017581b4b189726070e0017059b, /* 1558 */
128'h979b0027571b00b517bb020804630018, /* 1559 */
128'h4189d99b4187d79b8b050189999b0187, /* 1560 */
128'hfcc592e3872e0ff9f99300f9e9b3c70d, /* 1561 */
128'h00005517ef898b850a6a478302d98263, /* 1562 */
128'hf9b3fff7c793b591370020eff9c50513, /* 1563 */
128'h00005517cb898b8509ba4783bfd100f9, /* 1564 */
128'he20b02e3b51d547ddbaff0effcc50513, /* 1565 */
128'h45850af006134685e3958b850afa4783, /* 1566 */
128'h47830afa07a34785e569a21ff0ef854a, /* 1567 */
128'h4d010880049308f92a2300a7979b0e0a, /* 1568 */
128'h458586260ff6f69301acd6bb08c00d93, /* 1569 */
128'h2d210ff4f4932485ed499f1ff0ef854a, /* 1570 */
128'hf693019ad6bb08f00d134c81ffb492e3, /* 1571 */
128'h2485e9359cbff0ef854a458586260ff6, /* 1572 */
128'h09b00d934d61ffa492e32ca10ff4f493, /* 1573 */
128'h0196d6bb45858656000c26834c818aa6, /* 1574 */
128'h2ca12a85e13999dff0ef854a0ff6f693, /* 1575 */
128'h0c110ff4f493248dffac90e30ffafa93, /* 1576 */
128'hf0ef854a458509c0061386defdb498e3, /* 1577 */
128'h9b630a7a4783d4fb0de34785ed19975f, /* 1578 */
128'h957ff0ef854a458509b0061346850137, /* 1579 */
128'hf0ef854a45850a70061386cebb3d842a, /* 1580 */
128'h842ae406e0221141b32ddd79842a945f, /* 1581 */
128'h0187b303679c681c00055e63810ff0ef, /* 1582 */
128'h45058302014160a26402852200030763, /* 1583 */
128'hf822fc06f426713980820141640260a2, /* 1584 */
128'h92635529478500f5866384aa4791f04a, /* 1585 */
128'h842e07c4d78300f110230370079304f5, /* 1586 */
128'hc43ec24a8526858a46010107979b4955, /* 1587 */
128'h4791c24a00f110234799ed19d52ff0ef, /* 1588 */
128'hf0ef8526858a4601c43e478900f41f63, /* 1589 */
128'h478580826121790274a2744270e2d34f, /* 1590 */
128'hf3634f5c6918ee09b7cdc402fef414e3, /* 1591 */
128'h059b00e7f46385be27814f1887ae00f5, /* 1592 */
128'h80828082c2cff06f02c50823dd0c0007, /* 1593 */
128'hfc86f8a2070d4b9c711910000737691c, /* 1594 */
128'hf862fc5ee0dae4d6e8d2eccef0caf4a6, /* 1595 */
128'h681cc509f11ff0ef842ac17c8fd9f466, /* 1596 */
128'h05130000551702042423eb8d6b9c679c, /* 1597 */
128'h8526744670e6f8500493bacff0efdde5, /* 1598 */
128'h7c427be26b066aa66a4669e674a67906, /* 1599 */
128'hf93ff0eff3e54481541c808261097ca2, /* 1600 */
128'h02042c2302f4082347851af42c23478d, /* 1601 */
128'h681c421010ef7d000513ba2ff0ef8522, /* 1602 */
128'h08842783f94584aa97826b9c679c8522, /* 1603 */
128'hd85c478508f422231a04282318042e23, /* 1604 */
128'hf1dff0ef852245814601b72ff0ef8522, /* 1605 */
128'h45d000ef8522f14984aacf2ff0ef8522, /* 1606 */
128'h00ff8737681c00f1102347a1000505a3, /* 1607 */
128'h47d50aa00713e3991aa007138ff94bdc, /* 1608 */
128'he911bf8ff0efc23ec43a8522858a4601, /* 1609 */
128'h800207b700f715630aa0079300c14703, /* 1610 */
128'h02900a934a55037009933e900913cc1c, /* 1611 */
128'h460140000cb780020c3700ff8bb74b05, /* 1612 */
128'hbb6ff0efc402c252013110238522858a, /* 1613 */
128'hf7b3c25a4bdc015110234c18681ce13d, /* 1614 */
128'h4601c43e0197e7b301871563c43e0177, /* 1615 */
128'h0007ca6347b2ed1db8eff0ef8522858a, /* 1616 */
128'hbf45331010ef3e80051306090863397d, /* 1617 */
128'hcc188001073700e68563800207374c14, /* 1618 */
128'h478506041e23d45c8b8541e7d79bc43c, /* 1619 */
128'h852202f51f63f9200793b55d18f40ca3, /* 1620 */
128'h443ced09c34ff0ef85224581c04ff0ef, /* 1621 */
128'h85224585bfd118f40c2347850007d663, /* 1622 */
128'hf0efc5a5051300005517d965c1cff0ef, /* 1623 */
128'h7161551cb58584aab595fa100493a10f, /* 1624 */
128'hfadafed6e352e74eeb4aef26f706f322, /* 1625 */
128'h8baae3b54401e6eeeaeaeee6f2e2f6de, /* 1626 */
128'h198bc783c7b1199bc7831ff010ef4501, /* 1627 */
128'h479d460104f110234789e7b5180b8ca3, /* 1628 */
128'h00e3842aabaff0efc482c2be855e008c, /* 1629 */
128'h008c46014495cf818b851b8ba7831205, /* 1630 */
128'hf4fd34fd100503e3842aaa0ff0ef855e, /* 1631 */
128'hd55d842ad99ff0ef855ea031020ba423, /* 1632 */
128'h7af66a1a69ba695a64fa741a70ba8522, /* 1633 */
128'h8082615d6db66d566cf67c167bb67b56, /* 1634 */
128'hf0ef855e0407c163180b8c23048ba783, /* 1635 */
128'h091390810205149316d010ef4501b16f, /* 1636 */
128'ha783f155842ab36ff0ef855e45853e80, /* 1637 */
128'h12a96ee3149010ef85260007cc63048b, /* 1638 */
128'hac23400007b7bfe91d7010ef06400513, /* 1639 */
128'h02fba6238b8541e7d79b048ba78300fb, /* 1640 */
128'h45111aa60f63450dbf0506fb9e234785, /* 1641 */
128'h061b40010637a029400406370ea61ee3, /* 1642 */
128'h000039978a9d0036d61b00cbac234006, /* 1643 */
128'h0f86460396ce964e068a8a3d61498993, /* 1644 */
128'hd61b02d606bb018ba88345051086a683, /* 1645 */
128'h04cba823180bae231a0ba8238a0500c7, /* 1646 */
128'h183b8abd0107d69b08dba22308dba423, /* 1647 */
128'ha683090ba8231408dc63090ba62300d5, /* 1648 */
128'h571b003f06b70107979b14068e6302cb, /* 1649 */
128'h070907854721938117828fd98ff50107, /* 1650 */
128'h0c0bb0230a0bbc23030787b300e797b3, /* 1651 */
128'h0e0bb0230c0bbc230c0bb8230c0bb423, /* 1652 */
128'h08fba6230107d463200007930afbb823, /* 1653 */
128'h08fba82300e7f46320000793090ba703, /* 1654 */
128'h979b471100e78e63577d04cba783c215, /* 1655 */
128'hc282c4be04e11023855e008c46010107, /* 1656 */
128'h495507cbd78304f11023479d902ff0ef, /* 1657 */
128'hf0efc4bec2ca855e008c0107979b4601, /* 1658 */
128'h57fd08fbaa234785e40516e3842a8e4f, /* 1659 */
128'he2051ae3842ac9aff0ef855e08fb80a3, /* 1660 */
128'hffbfe0ef855e00b545830f7000ef855e, /* 1661 */
128'h07b754075a63018ba703e0051fe3842a, /* 1662 */
128'h06f110230370079304fba02327891000, /* 1663 */
128'hd2ca855e0107979b108c460107cbd783, /* 1664 */
128'h0bf104934905d2caed05880ff0efd4be, /* 1665 */
128'hd48206f11023988102091a9303300793, /* 1666 */
128'hec56e826855e108c08104b210a854a11, /* 1667 */
128'h842afe0a16e33a7dc131850ff0efd05a, /* 1668 */
128'hd59bbd9940030637a7a940020637bb45, /* 1669 */
128'h6685b54d08bba82300b515bb89bd0165, /* 1670 */
128'h17828fd501e7569b8ff50027979b16f1, /* 1671 */
128'h00ff05374098b5558b1d938100f7571b, /* 1672 */
128'h8e698fd50087161b0187179b0187569b, /* 1673 */
128'h8fd58ef1f00706138fd167410087569b, /* 1674 */
128'h0187169b0187559b40d804fbaa232781, /* 1675 */
128'h8f718ecd0087571b8de90087159b8ecd, /* 1676 */
128'h212700638b3d0187d71b04ebac238f55, /* 1677 */
128'h971300ebac238001073720d702634689, /* 1678 */
128'h8fd920000737040ba7830007596302d7, /* 1679 */
128'h1ef71863800107b7018ba70304fba023, /* 1680 */
128'h4d05040ba903639c0407879300005797, /* 1681 */
128'h849300003497020d1a13044ba783f0be, /* 1682 */
128'hfc1383f979130ff1079300f9793342e4, /* 1683 */
128'h00f977b300e797bb478540980a05fe07, /* 1684 */
128'h840b0b1b4a81017d8b37160785632781, /* 1685 */
128'hf7b300f977b340dc0007ac8397d6109c, /* 1686 */
128'h00fc8d6345a1400007b7140781630197, /* 1687 */
128'h85b3100005b700fc88634591200007b7, /* 1688 */
128'h1c638daa971ff0ef855e0015b59340bc, /* 1689 */
128'h2000073700ec8d6347a1400007370e05, /* 1690 */
128'hb79340fc8cb3100007b700ec88634791, /* 1691 */
128'h8663409cdfdfe0ef855e02fbaa23001c, /* 1692 */
128'h0af1102347994d850ce79163470d01a7, /* 1693 */
128'h00fde7b317c12d81810007b7d33e47d5, /* 1694 */
128'he552e162855e110c040007930110d53e, /* 1695 */
128'h94638bbd010c4783e941e91fe0efc93e, /* 1696 */
128'h088ba58314079a631afba823409c09b7, /* 1697 */
128'h460118fbae2308bba2230017b79317ed, /* 1698 */
128'h0793fe07fd930ff10793947ff0ef855e, /* 1699 */
128'h979b4601475507cbd7830af110230370, /* 1700 */
128'he0efd53ee03ad33a8cee855e110c0107, /* 1701 */
128'hd502d33a0af1102347b56702e915e35f, /* 1702 */
128'he16ee43e855e110c0110040007134791, /* 1703 */
128'h67a20e050c63e0dfe0efe03ac93ae552, /* 1704 */
128'h1afba823017d85b74785f3ed37fd6702, /* 1705 */
128'h855e840585934601180bae23096ba223, /* 1706 */
128'h379704a1eafa94e347a10a918c9ff0ef, /* 1707 */
128'h051300004517e6f49fe32aa787930000, /* 1708 */
128'h80011737b61ddf400413cbdfe0ef7365, /* 1709 */
128'h971300ebac2380020737b519a007071b, /* 1710 */
128'h04934905bbc580030737de075ee30307, /* 1711 */
128'h09053ac54a159881190201000ab70ff1, /* 1712 */
128'hc33e47d508f110234799020a08633a7d, /* 1713 */
128'hf84af426c556855e010c040007931030, /* 1714 */
128'h8b8583a54cdcd0051ce3d61fe0efdc3e, /* 1715 */
128'hd79b0087961bf006869366c144dcfbe1, /* 1716 */
128'hd9e3040ba70302e796938fd18ff50087, /* 1717 */
128'h4581472db35d04fba02300876793da06, /* 1718 */
128'h11872583974e837902079713eaf768e3, /* 1719 */
128'hf006869300ff0537040d859366c1b545, /* 1720 */
128'h8f510187971b0187d61b0d91000da783, /* 1721 */
128'h8fd98ff58f510087d79b8e690087961b, /* 1722 */
128'h579b46a5008ca703fdb59ee3fefdae23, /* 1723 */
128'h800306b7018ba60300f6f8638bbd00c7, /* 1724 */
128'h97b6078a0fc686930000369704d61c63, /* 1725 */
128'h00cca68308fbae230087171b1487a783, /* 1726 */
128'h0126d71b8fd10186d61b8ff917fd67c1, /* 1727 */
128'h073b3e800613c305c38d03f777132781, /* 1728 */
128'h02d606bb02f757bb8a8d0106d69b02e6, /* 1729 */
128'h1afbaa231b0ba7830adba2230afba023, /* 1730 */
128'ha82308fba62320000793c79919cba783, /* 1731 */
128'h0005062300051523484000ef855e08fb, /* 1732 */
128'haaa78793ccccd6b7aaaab7b708cba703, /* 1733 */
128'h068600d036b327818ef98ff9ccc68693, /* 1734 */
128'h8ef90f068693f0f0f6b79fb500f037b3, /* 1735 */
128'hf0068693ff0106b79fb5068a00d036b3, /* 1736 */
128'h0207161376c19fb5068e00d036b38ef9, /* 1737 */
128'h0a8bb783d11c9fb9071200e037338f75, /* 1738 */
128'h074bd68307abd70302c7d7b3ed109201, /* 1739 */
128'h0513572585930000459784aa06fbc603, /* 1740 */
128'hc883070ba803a95fe0effef536230245, /* 1741 */
128'h569b0108571b0088579b06cbc603077b, /* 1742 */
128'h26810ff777130ff878130ff7f7930188, /* 1743 */
128'ha5ffe0ef04d485135505859300004597, /* 1744 */
128'h0624851354c5859300004597074ba603, /* 1745 */
128'ha3ffe0ef8a3d8abd0146561b0106569b, /* 1746 */
128'h07b7b8d102fba42347857e4010ef8526, /* 1747 */
128'h1a0bb683400407b704fba02327851000, /* 1748 */
128'hbb954ca5051300004517e691ecf76ce3, /* 1749 */
128'h0c46c78304fba0230017079b70000737, /* 1750 */
128'hf693ce910027f6931adba42303f7f693, /* 1751 */
128'h040ba70304eba0230217071bc68900c7, /* 1752 */
128'h040ba783c7998b8504eba02301076713, /* 1753 */
128'h044ba783040baa0304fba02300c7e793, /* 1754 */
128'h0000349700fa7a33855e4601088ba583, /* 1755 */
128'h0b1300003b174a85db4ff0effac48493, /* 1756 */
128'h97bb409cff0c8c9300003c974c2dfbeb, /* 1757 */
128'h091300003917cbb5278100fa77b300fa, /* 1758 */
128'h00494703409c10000db720000d37f9e9, /* 1759 */
128'h0009270340dc04f718630017b79317ed, /* 1760 */
128'h0b70061300894683c3a18ff900fa77b3, /* 1761 */
128'h4681c131debfe0ef855e0fb6f6934585, /* 1762 */
128'h088ba783ddbfe0ef855e45850b700613, /* 1763 */
128'h035baa2308fba223180bae231a0ba823, /* 1764 */
128'h9fe304a1fb9911e30931973fe0ef855e, /* 1765 */
128'hbb6d925fe0ef39e5051300004517f764, /* 1766 */
128'h471100d789634721400006b700092783, /* 1767 */
128'h02ebaa230017b71341b787b301a78663, /* 1768 */
128'hf941808ff0ef855e408c933fe0ef855e, /* 1769 */
128'h1afba823409ce79d0046f79300892683, /* 1770 */
128'h08bba2230017b79317ed088ba583ef8d, /* 1771 */
128'he0ef855ecb0ff0ef855e460118fbae23, /* 1772 */
128'h45850b7006130ff6f693bb91fd319fdf, /* 1773 */
128'hfcfc65e34581b7c9f521d31fe0ef855e, /* 1774 */
128'h4641bf6d11872583974e837902079713, /* 1775 */
128'h04f11023478d6da000ef06cb851300ec, /* 1776 */
128'h855ec4be0107979b008c460107cbd783, /* 1777 */
128'ha783ec051b63842a96ffe0efc2be47d5, /* 1778 */
128'h47a506fb9e2304e157830007d663018b, /* 1779 */
128'h008c460107cbd783c2be479d04f11023, /* 1780 */
128'h1163842a93bfe0efc4be855e0107979b, /* 1781 */
128'hae23018ba50345e6475647c646b6ea05, /* 1782 */
128'h063706bba42306eba22306fba02304db, /* 1783 */
128'h02e345098a3d01a6d61bf2c51a634000, /* 1784 */
128'h40010637f0a609634505f0c543638ca6, /* 1785 */
128'he54ff06ffa100413f0eff06f2006061b, /* 1786 */
128'h0d238082557d8082557d80824501c56c, /* 1787 */
128'hef9d439cbf07879300005797808218b5, /* 1788 */
128'h2d2300005717842ae406e02247851141, /* 1789 */
128'h00055563aeefe0ef852212a000efbcf7, /* 1790 */
128'h00ef13e000ef02c00513fc5ff0ef8522, /* 1791 */
128'h80824501808201414501640260a20dc0, /* 1792 */
128'h02e790636394631cba87071300005717, /* 1793 */
128'he0efe40634c505130000451785aa1141, /* 1794 */
128'h0fc7a60380820141853e478160a2f60f, /* 1795 */
128'h110141488082853ebfd187b600a60463, /* 1796 */
128'h65a210354703c105fbdff0efe42eec06, /* 1797 */
128'h00f70c630ff007930815470302b70063, /* 1798 */
128'h8082610560e25535eb3fe06f610560e2, /* 1799 */
128'hec06e4261101bfcdf8400513bfe54501, /* 1800 */
128'hcf0ff0ef842acd09f7dff0ef84aee822, /* 1801 */
128'h610564a2644260e2e0800f840413e501, /* 1802 */
128'h43889927879300005797bfd555358082, /* 1803 */
128'h579780820f8505138082c3980015071b, /* 1804 */
128'h0000579711018082438897a787930000, /* 1805 */
128'h176384beec06e4266380e822adc78793, /* 1806 */
128'h19a447838082610564a2644260e20094, /* 1807 */
128'h00005797b7d56000a9cff0ef8522c781, /* 1808 */
128'h9207a82300005797e79ce39caac78793, /* 1809 */
128'he7886798a947879300005797e5088082, /* 1810 */
128'h00005497e4a6711d8082e308e518e11c, /* 1811 */
128'hf05af456f852fc4e6080e8a2a7c48493, /* 1812 */
128'h4a1789aae0caec86e06ae466e862ec5e, /* 1813 */
128'h4b1722aa8a9300004a9723aa0a130000, /* 1814 */
128'h0c1b232b8b9300004b97232b0b130000, /* 1815 */
128'h029415634d29816c8c9300004c970005, /* 1816 */
128'h7b027aa27a4279e2690664a660e66446, /* 1817 */
128'h38050513000045176d026ca26c426be2, /* 1818 */
128'h89524c1cc7914901541cddcfe06f6125, /* 1819 */
128'h638c855a0fc42603681c89560007c363, /* 1820 */
128'hdb2fe0ef855e85ca00090663dbefe0ef, /* 1821 */
128'h8863da4fe0ef856685e200978e63601c, /* 1822 */
128'h600032a010ef79e505130000351701a9, /* 1823 */
128'hc1414401e04ae426ec06e8221101b771, /* 1824 */
128'h651ccbad511ccbbd4d5ccfad44014d1c, /* 1825 */
128'h45051c00059384aa892ec7ad639cc7bd, /* 1826 */
128'h2c234799c57c57fdcd21842a200010ef, /* 1827 */
128'h282303253023e90410f502a347850ef5, /* 1828 */
128'h3c2391c78793fffff797e65ff0ef0405, /* 1829 */
128'h179718f430232be787930000179716f4, /* 1830 */
128'h0ea42e23681c18f434232ae787930000, /* 1831 */
128'h8522e99ff0ef10f400230247c7838522, /* 1832 */
128'h1bc0106f80826105690264a2644260e2, /* 1833 */
128'h86b365186294611c6b86869300004697, /* 1834 */
128'h8f3d0127d713e11897360017671302d7, /* 1835 */
128'h00f717bb40f007b300f7553b93ed836d, /* 1836 */
128'hf06f8f25051300005517808225018d5d, /* 1837 */
128'hf0ef842afefff0efe022e4061141fc3f, /* 1838 */
128'h01412501640260a28d410105151bfe9f, /* 1839 */
128'h0005041bfdbff0efe022e40611418082, /* 1840 */
128'h640260a28d4115029001fd1ff0ef1402, /* 1841 */
128'h8fa30785fff5c703058587aa80820141, /* 1842 */
128'h058500c7896387aa962a8082fb75fee7, /* 1843 */
128'h87aa8082fb65fee78fa30785fff5c703, /* 1844 */
128'hfff5c7030585eb09001786930007c703, /* 1845 */
128'h87aab7d587b68082fb75fee78fa30785, /* 1846 */
128'hfb7d001786930007c70387b68082e219, /* 1847 */
128'hfed70fa300178713fff5c6830585963e, /* 1848 */
128'h87ba8082000780a300c715638082e291, /* 1849 */
128'h40f707bbfff5c783000547030585b7cd, /* 1850 */
128'h853ef37d0505e3994187d79b0187979b, /* 1851 */
128'h47030585a839478100c59463962e8082, /* 1852 */
128'hd79b0187979b40f707bbfff5c7830005, /* 1853 */
128'h0ff5f5938082853eff790505e3994187, /* 1854 */
128'hbfcd0505c399808200b7936300054783, /* 1855 */
128'h00b79363000547830ff5f59380824501, /* 1856 */
128'he7010007c70387aabfcd0505dffd8082, /* 1857 */
128'he42ee8221101bfcd0785808240a78533, /* 1858 */
128'h0ff5f593952265a2fe5ff0efec06842a, /* 1859 */
128'h4501fe857be3157d00b7866300054783, /* 1860 */
128'h00b7856387aa95aa80826105644260e2, /* 1861 */
128'hb7fd0785808240a78533e7010007c703, /* 1862 */
128'h8082ea9940c785330007c68387aa862a, /* 1863 */
128'h0785fe081be3000748030705fed80fe3, /* 1864 */
128'h85330007c60387aa86aabfcd872eb7d5, /* 1865 */
128'h00074803070500c80a638082ea1140d7, /* 1866 */
128'h4703bff90785bfd5872e8082fe081be3, /* 1867 */
128'hc6830785fee68fe380824501eb190005, /* 1868 */
128'he8221101bfd587aeb7e50505fafd0007, /* 1869 */
128'h879300004797e519842a84aeec06e426, /* 1870 */
128'h942af9dff0ef85a68522cc1163806ee7, /* 1871 */
128'h44016c07b92300004797ef8100044783, /* 1872 */
128'h852285a68082610564a2644260e28522, /* 1873 */
128'h00050023c78100054783c519f9fff0ef, /* 1874 */
128'he4261101bfd96aa7b323000047970505, /* 1875 */
128'hf73ff0ef8526842ac891e822ec066104, /* 1876 */
128'h8526644260e2e008050500050023c501, /* 1877 */
128'h87aacf9900054783c11d8082610564a2, /* 1878 */
128'h80238082e3110017c703ce810007c683, /* 1879 */
128'h779380824501b7e5078900d780a300e7, /* 1880 */
128'h07a2808204c79063963e87aacb9d0075, /* 1881 */
128'h8833469d00c508b3872aff6d377d8fd5, /* 1882 */
128'h02e787335761003657930106ef6340e8, /* 1883 */
128'hbfd10ff5f6934725bfc1963a97aa078e, /* 1884 */
128'hbf6dfeb78fa30785bfe1fef73c230721, /* 1885 */
128'h963e87aacb9d8b9d00a5e7b300b50a63, /* 1886 */
128'hbc2307a1ff8738030721808202c79e63, /* 1887 */
128'h57e100365713ff06e8e340f88833ff07, /* 1888 */
128'hbfc100e507b3963e95ba070e02f707b3, /* 1889 */
128'hc7030585bfe1469d00c508b387aa872e, /* 1890 */
128'h842af0227179bf65fee78fa30785fff5, /* 1891 */
128'hdcdff0efe02ee84af406e432ec26852e, /* 1892 */
128'h091300c564636582892ace1184aa6622, /* 1893 */
128'h00040023f79ff0ef944a864a8522fff6, /* 1894 */
128'h11418082614564e269428526740270a2, /* 1895 */
128'h8522f57ff0ef00a5e963842ae406e022, /* 1896 */
128'h073300c506b395b280820141640260a2, /* 1897 */
128'h16fd0005c78315fdd7e500e587b340b6, /* 1898 */
128'h853e478100c51563962ab7fd00f68023, /* 1899 */
128'h0505fbed9f990005c703000547838082, /* 1900 */
128'h00054783808200c51363962ab7dd0585, /* 1901 */
128'h852e842af0227179bfc50505feb78de3, /* 1902 */
128'h049bd1fff0ef89aee84af406e44eec26, /* 1903 */
128'h5b630005091bd13ff0ef8522c8890005, /* 1904 */
128'h69a2694264e2740270a2852244010099, /* 1905 */
128'hf8bff0ef397d852285ce862680826145, /* 1906 */
128'h00c514630ff5f593962abfe90405d175, /* 1907 */
128'hfeb70be3001507930005470380824501, /* 1908 */
128'h260100c7ef630ff5f59347c1b7ed853e, /* 1909 */
128'h1ce30007c7038082853e4781e60187aa, /* 1910 */
128'h47a1c31d00757713b7f5367d0785feb7, /* 1911 */
128'h1ce30007c80387aa0007069b40e7873b, /* 1912 */
128'h953e938102071793faf5078536fdfcb8, /* 1913 */
128'h8fd90107179300b7e733008597938e1d, /* 1914 */
128'heb1187aa27018edd0036571302079693, /* 1915 */
128'h367d0785f8b71fe30007c703d24d8a1d, /* 1916 */
128'hc70300d80a63008785130007b803bfcd, /* 1917 */
128'h87aabfa5fef51be30785f8b712e30007, /* 1918 */
128'h0300079300054703e7a9419cb7f1377d, /* 1919 */
128'h0f878793000027970015470308f71163, /* 1920 */
128'h0207071bc6898a850006c68300e786b3, /* 1921 */
128'h0025470304d71b63078006930ff77713, /* 1922 */
128'hc19c47c1c3b10447f7930007c78397ba, /* 1923 */
128'h030007930005470302f71c6347c14198, /* 1924 */
128'h0a870713000027170015478302f71663, /* 1925 */
128'hf7930207879bc7098b0500074703973e, /* 1926 */
128'h47a18082050900e79363078007130ff7, /* 1927 */
128'hec06006c842ee8221101bf6d47a9bf7d, /* 1928 */
128'h00002817468100c16583f63ff0efc632, /* 1929 */
128'h00f806330007079b0005470306480813, /* 1930 */
128'h60e2ec05000898630446789300064603, /* 1931 */
128'h00088b63004678938082610585366442, /* 1932 */
128'h96be050502d586b3feb7f4e3fd07879b, /* 1933 */
128'h879b0ff7f793fe07079bc6098a09b7d1, /* 1934 */
128'hfc06f426f8227139b7e1e008b7cdfc97, /* 1935 */
128'hb0dff0ef84b2842ae42e00063023f04a, /* 1936 */
128'h6121790274a2744270e25529e90165a2, /* 1937 */
128'h67e2f5dff0ef8522082c892a862e8082, /* 1938 */
128'h9be307858f81cb010007c703fe8782e3, /* 1939 */
128'h4683b7e94501e088fcf718e347a9fd27, /* 1940 */
128'h1141f2dff06f00e6846302d007130005, /* 1941 */
128'h014140a0053360a2f23ff0efe4060505, /* 1942 */
128'h601cf0dff0ef842ee406e02211418082, /* 1943 */
128'h00e6ea6302d704630007c70304b00693, /* 1944 */
128'h80820141640260a202d70e6304700693, /* 1945 */
128'hfed716e306b0069302d7076304d00693, /* 1946 */
128'hc683fce69fe3052a069007130017c683, /* 1947 */
128'hb7e9e01c078d00e69863042007130027, /* 1948 */
128'h842ee8221101bfd50789bff1052a052a, /* 1949 */
128'h468100c16583e0fff0efc632ec06006c, /* 1950 */
128'h0007079b00054703f108081300002817, /* 1951 */
128'h00089863044678930006460300f80633, /* 1952 */
128'h00467893808261058536644260e2ec05, /* 1953 */
128'h02d586b3feb7f4e3fd07879b00088b63, /* 1954 */
128'hf793fe07079bc6098a09b7d196be0505, /* 1955 */
128'he0221141b7e1e008b7cdfc97879b0ff7, /* 1956 */
128'hc70304b00693601cf87ff0ef842ee406, /* 1957 */
128'h0e630470069300e6ea6302d704630007, /* 1958 */
128'h076304d0069380820141640260a202d7, /* 1959 */
128'h07130017c683fed716e306b0069302d7, /* 1960 */
128'h042007130027c683fce69fe3052a0690, /* 1961 */
128'hbff1052a052ab7e9e01c078d00e69863, /* 1962 */
128'hf0efe589842ae406e0221141bfd50789, /* 1963 */
128'h879300002797fff5c70300a405b395bf, /* 1964 */
128'he7198b1100074703973efff58513e367, /* 1965 */
128'hfea47ae3157d80820141557d640260a2, /* 1966 */
128'h6402f77d8b1100074703973e00054703, /* 1967 */
128'h4581d7dff06f014105054581462960a2, /* 1968 */
128'h00a10723812100a107a31141fa5ff06f, /* 1969 */
128'h2c878793000047978082014100e15503, /* 1970 */
128'haa5ff06f95be9201160291811582639c, /* 1971 */
128'h8082853ee3190005470345a946254781, /* 1972 */
128'h02f587bb00d667630ff6f693fd07069b, /* 1973 */
128'he406e0221141bff90505fd07879b9fb9, /* 1974 */
128'h55bb45a900b7f86347a500a04563842e, /* 1975 */
128'h640202a4753b4529fe7ff0ef357d02b4, /* 1976 */
128'h081007935000006f03050513014160a2, /* 1977 */
128'h37230000471724f737230000471707e2, /* 1978 */
128'h2404041300004417e8221101808224f7, /* 1979 */
128'ha15ff0efec06600885aa84ae862ee426, /* 1980 */
128'h8082610564a26442e00c95a660e2600c, /* 1981 */
128'h00004497e42621678793000047971101, /* 1982 */
128'h0513000035176380e822609020448493, /* 1983 */
128'h85a26088b87fd0ef85a29c11ec067be5, /* 1984 */
128'h051300003517862286aa608ce63fc0ef, /* 1985 */
128'hd0ef7c25051300003517b6dfd0ef7b65, /* 1986 */
128'h5e6385df90efef65051300000517b61f, /* 1987 */
128'h0000351740a005b364a260e264420005, /* 1988 */
128'h64a260e26442b39fd06f61057b450513, /* 1989 */
128'ha0ef8432e406e02211416680006f6105, /* 1990 */
128'h80820141640260a2557d0085036387ef, /* 1991 */
128'h89aae64e01258413f222716980824501, /* 1992 */
128'h0505f7eff0ef892eea4aee26f6068522, /* 1993 */
128'hf0ef95260505f72ff0ef852600a404b3, /* 1994 */
128'h479704e7ee631ff00793fff5071be93f, /* 1995 */
128'h351784aaf50ff0ef852212a7a5230000, /* 1996 */
128'h0ff007939526f42ff0ef52a505130000, /* 1997 */
128'h00003517842af32ff0ef852204a7f263, /* 1998 */
128'h0000351700a405b3f24ff0ef50c50513, /* 1999 */
128'h695264f2741270b2a8bfd0ef72450513, /* 2000 */
128'h272300004717200007938082615569b2, /* 2001 */
128'h863ff0ef850a458110000613b7550cf7, /* 2002 */
128'h4703deaff0ef850a4c85859300003597, /* 2003 */
128'h85930000359700f7096302f007930129, /* 2004 */
128'hdf2ff0ef850a85a2dfaff0ef850a6f65, /* 2005 */
128'h00003517858a43900887879300004797, /* 2006 */
128'h451107e208100793a1bfd0ef6dc50513, /* 2007 */
128'h06f738230000471706f7382300004717, /* 2008 */
128'hf0ef4501e4a7962300004797d85ff0ef, /* 2009 */
128'h000045974611e4a7902300004797d77f, /* 2010 */
128'h000047174785eb1ff0ef854ee3458593, /* 2011 */
128'he04ae426ec06e8221101b79102f71823, /* 2012 */
128'hf0ef84ae450d892a08c7df638432478d, /* 2013 */
128'h0000451708a7956325010004d783d37f, /* 2014 */
128'h9a6325010024d783d21ff0ef00055503, /* 2015 */
128'h4511dabff0ef00448513ffc4059b06a7, /* 2016 */
128'h00004517dca7962300004797d05ff0ef, /* 2017 */
128'h9c23000047974611cf1ff0effd055503, /* 2018 */
128'he2bff0ef854adae5859300004597daa7, /* 2019 */
128'h4515fa65d58300004597256000ef4535, /* 2020 */
128'h00004797240000ef02000513d1bff0ef, /* 2021 */
128'h11230000471727850007d783f9078793, /* 2022 */
128'hcf63278d439cf767879300004797f8f7, /* 2023 */
128'h6442905fd0ef5e650513000035170087, /* 2024 */
128'h644260e2d49ff06f6105690264a260e2, /* 2025 */
128'hc783f022f406717980826105690264a2, /* 2026 */
128'h00f10f230115c78300f10fa347090105, /* 2027 */
128'h740202e78a63470d00e78e6301e15783, /* 2028 */
128'h8b3fd06f61455c6505130000351770a2, /* 2029 */
128'h8a3fd0efe42e59e5051300003517842a, /* 2030 */
128'h7402d8bff06f614570a265a274028522, /* 2031 */
128'hdc010113ebfff06f614505c170a24190, /* 2032 */
128'h84ae842a232130232291342322813823, /* 2033 */
128'hf0ef22113c2300282180061345818932, /* 2034 */
128'hf0efe802c44a08282040061385a6e60f, /* 2035 */
128'h340323813083f63ff0ef8522002cea2f, /* 2036 */
128'h80822401011322013903228134832301, /* 2037 */
128'h000045974611cb81e8c7d78300004797, /* 2038 */
128'h00efe40611418082cf3ff06fc7458593, /* 2039 */
128'h1001a70300e57763878e1041e7035040, /* 2040 */
128'h60a21007e78310a7a22310e1a0232705, /* 2041 */
128'h80824501808201418d5d910117821502, /* 2042 */
128'h842afc1ff0ef84aae426e822ec061101, /* 2043 */
128'h9101150202f407b33e800793440000ef, /* 2044 */
128'h8082610564a28d0502a7d533644260e2, /* 2045 */
128'h414000ef842af95ff0efe022e4061141, /* 2046 */
128'h640260a202f407b324078793000f47b7, /* 2047 */
128'hec061101808202a7d533014191011502, /* 2048 */
128'h00ef892af63ff0ef84aae04ae426e822, /* 2049 */
128'h543324040413000f443702a485333e20, /* 2050 */
128'h60e2fe856ee3f45ff0ef0405944a0285, /* 2051 */
128'h94b7e426110180826105690264a26442, /* 2052 */
128'h892268048493842ae04aec06e8220098, /* 2053 */
128'hfa1ff0ef41240433854a89260084f363, /* 2054 */
128'h002380826105690264a2644260e2f47d, /* 2055 */
128'hc503100007b7808200054503808200b5, /* 2056 */
128'h01474783100007378082020575130147, /* 2057 */
128'h100007b7808200a70023dfe50207f793, /* 2058 */
128'h8023476d00e78623f800071300078223, /* 2059 */
128'hfc70071300e78623470d0007822300e7, /* 2060 */
128'h1141808200e788230200071300e78423, /* 2061 */
128'h640260a2e50900044503842ae406e022, /* 2062 */
128'h00002797b7f50405fa5ff0ef80820141, /* 2063 */
128'h470397aa973e811100f57713d5c78793, /* 2064 */
128'h808200f5802300e580a30007c7830007, /* 2065 */
128'hfd1ff0efec068121842a002ce8221101, /* 2066 */
128'hf5dff0ef00914503f65ff0ef00814503, /* 2067 */
128'hf0ef00814503fb7ff0ef0ff47513002c, /* 2068 */
128'h6105644260e2f43ff0ef00914503f4bf, /* 2069 */
128'h4461892af406e84aec26f02271798082, /* 2070 */
128'hf81ff0ef0ff57513002c0089553b54e1, /* 2071 */
128'hf0ef00914503f13ff0ef346100814503, /* 2072 */
128'h6145694264e2740270a2fe9410e3f0bf, /* 2073 */
128'h0413892af406e84aec26f02271798082, /* 2074 */
128'hf0ef0ff57513002c0089553354e10380, /* 2075 */
128'h00914503ed1ff0ef346100814503f3ff, /* 2076 */
128'h694264e2740270a2fe9410e3ec9ff0ef, /* 2077 */
128'h4503f13ff0efec06002c110180826145, /* 2078 */
128'h60e2e9fff0ef00914503ea7ff0ef0081, /* 2079 */
128'h7139439ce34787930000479780826105, /* 2080 */
128'h84b2842e892aec4efc06f04af426f822, /* 2081 */
128'hf3afb0efbdc505130000451702b78563, /* 2082 */
128'h744270e2e0a7a42300004797c10d2501, /* 2083 */
128'h0000471757fd8082612169e2790274a2, /* 2084 */
128'h05130000451785ca86260074def72623, /* 2085 */
128'ha92300004797c50d2501814fb0efba65, /* 2086 */
128'h05130000351785a6049675634632dca7, /* 2087 */
128'hdaf72a23000047174785d0cfd0ef23e5, /* 2088 */
128'h0009099b00c4591be05ff0ef4521b775, /* 2089 */
128'h4503993e003979132387879300003797, /* 2090 */
128'h9c25bf5d320010ef854ede7ff0ef0009, /* 2091 */
128'h85aae0221141bf95d687ac2300004797, /* 2092 */
128'hcb2fd0efe40620e5051300003517842a, /* 2093 */
128'h64028322f14025730ff0000f0000100f, /* 2094 */
128'h114183020141bbe585930000259760a2, /* 2095 */
128'h051300004517ef658593000035974605, /* 2096 */
128'h3517c9112501d79fa0efe022e406d365, /* 2097 */
128'hc62fd06f014160a264021f2505130000, /* 2098 */
128'h35974605c56fd0ef2005051300003517, /* 2099 */
128'ha0efaba5051300004517212585930000, /* 2100 */
128'hb7e120a5051300003517c5112501d9bf, /* 2101 */
128'h00000517c26fd0ef0885051300003517, /* 2102 */
128'h00004797cc07a42300004797e9850513, /* 2103 */
128'h479700054863842a912f90efca07ae23, /* 2104 */
128'h6402408005b3cf81439ccae787930000, /* 2105 */
128'hbe2fd06f014105e505130000351760a2, /* 2106 */
128'hc5112501b9afb0efa505051300004517, /* 2107 */
128'h000035974605bfb91b85051300003517, /* 2108 */
128'h3517c5112501cb9fa0ef4501e2c58593, /* 2109 */
128'h0023ee1ff0ef8522b7811b2505130000, /* 2110 */
128'ha001d69ff0efe4062501114190020000, /* 2111 */
128'h471780824501808224050513000f4537, /* 2112 */
128'h869300756513157d631cc22707130000, /* 2113 */
128'h8082953e055e10d00513e30895360017, /* 2114 */
128'hf0efe4328532ec06e822110102b50633, /* 2115 */
128'h8522944ff0ef45816622c509842afd1f, /* 2116 */
128'h000035171141808280826105644260e2, /* 2117 */
128'hc0ef20000537b28fd0efe40614c50513, /* 2118 */
128'h45018082450180820141450160a2ee5f, /* 2119 */
128'h1141808202f5553347a9b00025738082, /* 2120 */
128'h138505130000351785aa862e86b28736, /* 2121 */
128'h1141a001cbbff0ef4505aecfd0efe406, /* 2122 */
128'h408007b3f57ff0efe406952e842ae022, /* 2123 */
128'h80824505808201418d7d640260a29522, /* 2124 */
128'hf406ec26f02271798082450580824505, /* 2125 */
128'h64e2740270a20096186300c684bb842e, /* 2126 */
128'he37fc0efe432852285b2808261454501, /* 2127 */
128'h450980824509bff92605200404136622, /* 2128 */
128'h80824501808280828082808245098082, /* 2129 */
128'he426e822ec061101bbbff06f80824501, /* 2130 */
128'h986300d5043300d584b3003796934781, /* 2131 */
128'h380380826105450164a2644260e200c7, /* 2132 */
128'h000035176090600c02e8036360980004, /* 2133 */
128'h0000351785a28626a2afd0ef0ac50513, /* 2134 */
128'h711dbf5d0785a001a1afd0ef0c450513, /* 2135 */
128'hfc4ee8a20c45051300003517892ae0ca, /* 2136 */
128'he466e4a6ec86e862ec5ef05af456f852, /* 2137 */
128'h0b0a0a1300003a179eafd0ef44018b2e, /* 2138 */
128'h00003c17fff949930b8b8b9300003b97, /* 2139 */
128'h00040c9b9c6fd0ef85524ac10bcc0c13, /* 2140 */
128'h03649863448187ca9bafd0ef855e85e6, /* 2141 */
128'h87ca9a4fd0ef856285e69acfd0ef8552, /* 2142 */
128'h00003517fd5417e3040502b49b634581, /* 2143 */
128'h008486b3a889450198afd0ef0e450513, /* 2144 */
128'he39840e9873300349713c689873e8a85, /* 2145 */
128'h8a856390008586b3bf5d07a104856398, /* 2146 */
128'h02e60d6340e9873300359713c689873e, /* 2147 */
128'h3517944fd0ef0465051300003517058e, /* 2148 */
128'h644660e6557d938fd0ef072505130000, /* 2149 */
128'h6c426be27b027aa27a4279e2690664a6, /* 2150 */
128'he0d27159bfa507a10585808261256ca2, /* 2151 */
128'hf85ae4ceeca6020005138aaa6a05fc56, /* 2152 */
128'he46ee86aec66e8caf0a2f486f062f45e, /* 2153 */
128'h9c4a0a134981b3fff0ef44818bb28b2e, /* 2154 */
128'h00fa8db3003497933a8c0c1300003c17, /* 2155 */
128'h040505130000351703749b6300fb0cb3, /* 2156 */
128'h7ba26a0669a6694670a674068befd0ef, /* 2157 */
128'h7b4264e685da86266da26d426ce27c02, /* 2158 */
128'h842abddfe0efe33ff06f61657ae28556, /* 2159 */
128'hbcbfe0ef892abd1fe0ef8d2abd7fe0ef, /* 2160 */
128'h00a96533010d1d1b0105151b0344f7b3, /* 2161 */
128'h00acb0238d4191011402150201a46433, /* 2162 */
128'hf7930985aadff0ef4521ef8100adb023, /* 2163 */
128'hb7ad0485a9dff0ef0007c50397e20039, /* 2164 */
128'hec4ef04af426f822fc06e032e42e7139, /* 2165 */
128'he0ef892ab6ffe0ef842ab75fe0ef89aa, /* 2166 */
128'h0109179b0105151bb63fe0ef84aab69f, /* 2167 */
128'h8d5d9101178265a2660215028fc18d45, /* 2168 */
128'h00c79c63974e00e58833003797134781, /* 2169 */
128'h6121863e69e2854e790274a270e27442, /* 2170 */
128'h00083703e3148ea907856314d79ff06f, /* 2171 */
128'hfc06e032e42e7139b7f100e830238f29, /* 2172 */
128'h842aafdfe0ef89aaec4ef04af426f822, /* 2173 */
128'haebfe0ef84aaaf1fe0ef892aaf7fe0ef, /* 2174 */
128'h660215028fc18d450109179b0105151b, /* 2175 */
128'h88330037971347818d5d9101178265a2, /* 2176 */
128'h790274a270e2744200c79c63974e00e5, /* 2177 */
128'h07856314d01ff06f6121863e69e2854e, /* 2178 */
128'hb7f100e830238f0900083703e3148e89, /* 2179 */
128'hec4ef04af426f822fc06e032e42e7139, /* 2180 */
128'he0ef892aa7ffe0ef842aa85fe0ef89aa, /* 2181 */
128'h0109179b0105151ba73fe0ef84aaa79f, /* 2182 */
128'h8d5d9101178265a2660215028fc18d45, /* 2183 */
128'h00c79c63974e00e58833003797134781, /* 2184 */
128'h6121863e69e2854e790274a270e27442, /* 2185 */
128'h3703e31402a686b307856314c89ff06f, /* 2186 */
128'he42e7139b7e100e8302302a707330008, /* 2187 */
128'he0ef89aaec4ef04af426f822fc06e032, /* 2188 */
128'h84aa9fdfe0ef892aa03fe0ef842aa09f, /* 2189 */
128'h8fc18d450109179b0105151b9f7fe0ef, /* 2190 */
128'h971347818d5d9101178265a266021502, /* 2191 */
128'h70e2744200c79c63974e00e588330037, /* 2192 */
128'hc0dff06f6121863e69e2854e790274a2, /* 2193 */
128'h3703e31402a6d6b3078563144505e111, /* 2194 */
128'he42e7139b7d100e8302302a757330008, /* 2195 */
128'he0ef89aaec4ef04af426f822fc06e032, /* 2196 */
128'h84aa97dfe0ef892a983fe0ef842a989f, /* 2197 */
128'h8fc18d450109179b0105151b977fe0ef, /* 2198 */
128'h971347818d5d9101178265a266021502, /* 2199 */
128'h70e2744200c79c63974e00e588330037, /* 2200 */
128'hb8dff06f6121863e69e2854e790274a2, /* 2201 */
128'h30238f4900083703e3148ec907856314, /* 2202 */
128'hf426f822fc06e032e42e7139b7f100e8, /* 2203 */
128'h90bfe0ef842a911fe0ef89aaec4ef04a, /* 2204 */
128'h0105151b8fffe0ef84aa905fe0ef892a, /* 2205 */
128'h178265a2660215028fc18d450109179b, /* 2206 */
128'h974e00e588330037971347818d5d9101, /* 2207 */
128'h69e2854e790274a270e2744200c79c63, /* 2208 */
128'he3148ee907856314b15ff06f6121863e, /* 2209 */
128'he42e7139b7f100e830238f6900083703, /* 2210 */
128'he0ef89aaec4ef04af426f822fc06e032, /* 2211 */
128'h84aa88dfe0ef892a893fe0ef842a899f, /* 2212 */
128'h8fc18cc90109179b0105151b887fe0ef, /* 2213 */
128'h169347018fc59081178265a266021482, /* 2214 */
128'h70e2744200c71c6396ae00d988330037, /* 2215 */
128'ha9dff06f6121863a69e2854e790274a2, /* 2216 */
128'h7159bfc9070500a83023e28800f70533, /* 2217 */
128'he4cef0a2ba45051300003517892ae8ca, /* 2218 */
128'hec66eca6f486f062f45ef85afc56e0d2, /* 2219 */
128'h0a1300003a17cc9fc0ef44018b3289ae, /* 2220 */
128'h0c1300003c17b96b8b9300003b97b8ea, /* 2221 */
128'hfff44493ca7fc0ef855204000a93b9ec, /* 2222 */
128'h460140900cb3c99fc0ef8885855e85a2, /* 2223 */
128'h0566186397ce00f905b30036179314fd, /* 2224 */
128'hc73fc0ef856285a2c7bfc0efe4328552, /* 2225 */
128'h2405e12984aaa03ff0ef854a85ce6622, /* 2226 */
128'hc53fc0efbac5051300003517fb541be3, /* 2227 */
128'h7ae26a0669a664e669468526740670a6, /* 2228 */
128'h00167693808261656ce27c027ba27b42, /* 2229 */
128'h54fdbf590605e198e3988726c2918766, /* 2230 */
128'had0505130000351784aaeca67159bfc1, /* 2231 */
128'hf062f45ef85afc56e0d2e4cee8caf0a2, /* 2232 */
128'hbf3fc0ef44018ab2892ee86af486ec66, /* 2233 */
128'hdb8b0b1300003b17ab89899300003997, /* 2234 */
128'hab0c0c1300003c17db8b8b9300003b97, /* 2235 */
128'hc0ef854e04000a13ab8c8c9300003c97, /* 2236 */
128'h856285a2000bbd03cba500147793bc1f, /* 2237 */
128'h85b300361793fffd45134601baffc0ef, /* 2238 */
128'hb93fc0efe432854e05561c6397ca00f4, /* 2239 */
128'hf0ef852685ca6622b8bfc0ef856685a2, /* 2240 */
128'h00003517fb441ae32405e5298d2a91bf, /* 2241 */
128'h64e6856a740670a6b6bfc0efac450513, /* 2242 */
128'h6ce27c027ba27b427ae26a0669a66946, /* 2243 */
128'h00167693bf49000b3d03808261656d42, /* 2244 */
128'h5d7db7790605e198e398872ac291876a, /* 2245 */
128'h9e05051300003517842ae8a2711db7e1, /* 2246 */
128'hec86e862ec5ef05af456f852e0cae4a6, /* 2247 */
128'h00003917b07fc0ef4c018ab284aefc4e, /* 2248 */
128'h00003b979d4b0b1300003b179cc90913, /* 2249 */
128'h099bae5fc0ef854a10000a139dcb8b93, /* 2250 */
128'h1793008c1713ad9fc0ef855a85ce000c, /* 2251 */
128'h17138fd9018c17130187e7b38fd9010c, /* 2252 */
128'h8fd9030c17138fd9028c17138fd9020c, /* 2253 */
128'h00e406b30036171346018fd9038c1713, /* 2254 */
128'h85cea95fc0efe432854a055617639726, /* 2255 */
128'h81dff0ef852285a66622a8dfc0ef855e, /* 2256 */
128'h051300003517f94c19e30c05e91d89aa, /* 2257 */
128'h690664a6854e644660e6a6dfc0ef9c65, /* 2258 */
128'h808261256c426be27b027aa27a4279e2, /* 2259 */
128'hf4a67119bff159fdb74d0605e29ce31c, /* 2260 */
128'heccef0caf8a28f6505130000351784aa, /* 2261 */
128'hfc86f06af466f862fc5ee0dae4d6e8d2, /* 2262 */
128'h00003a17a17fc0ef44018b32892eec6e, /* 2263 */
128'h07f00b938e4c8c9300003c978dca0a13, /* 2264 */
128'h0a938e2d0d1300003d1703f00c134985, /* 2265 */
128'h9e3fc0ef856685a29ebfc0ef85520800, /* 2266 */
128'h17934601008995b300e99733408b873b, /* 2267 */
128'he432855205661a6397ca00f486b30036, /* 2268 */
128'h85ca66229b7fc0ef856a85a29bffc0ef, /* 2269 */
128'hfb541be32405e1398daaf46ff0ef8526, /* 2270 */
128'h744670e6997fc0ef8f05051300003517, /* 2271 */
128'h7be26b066aa66a4669e6790674a6856e, /* 2272 */
128'h008c6663808261096de27d027ca27c42, /* 2273 */
128'h5dfdbfe5e298e398bf610605e28ce38c, /* 2274 */
128'h810505130000351784aaf4a67119b7f1, /* 2275 */
128'hf862fc5ee0dae4d6e8d2eccef0caf8a2, /* 2276 */
128'hc0ef44018b32892eec6efc86f06af466, /* 2277 */
128'h8c9300002c977f6a0a1300002a17931f, /* 2278 */
128'h00002d1703f00c13498507f00b937fec, /* 2279 */
128'h85a2905fc0ef855208000a937fcd0d13, /* 2280 */
128'h96b300f997b3408b87bb8fdfc0ef8566, /* 2281 */
128'h003617134601fff6c693fff7c7930089, /* 2282 */
128'hc0efe432855205661a63974a00e485b3, /* 2283 */
128'h852685ca66228c9fc0ef856a85a28d1f, /* 2284 */
128'h3517fb5417e32405e1398daae58ff0ef, /* 2285 */
128'h856e744670e68a9fc0ef802505130000, /* 2286 */
128'h7c427be26b066aa66a4669e6790674a6, /* 2287 */
128'he314008c6663808261096de27d027ca2, /* 2288 */
128'hb7f15dfdbfe5e19ce31cbf610605e194, /* 2289 */
128'hf8a2722505130000251784aaf4a67119, /* 2290 */
128'hf466f862fc5ee0dae4d6e8d2eccef0ca, /* 2291 */
128'h843fc0ef44018a32892eec6efc86f06a, /* 2292 */
128'h710c0c1300002c177089899300002997, /* 2293 */
128'h2c9703f00b9308100b134d0507f00a93, /* 2294 */
128'h856285a2817fc0ef854e70ac8c930000, /* 2295 */
128'h00fd17b3408b07bb408a873b80ffc0ef, /* 2296 */
128'h16b300fd17b30024079b8f5d00ed1733, /* 2297 */
128'h16934601fff7c313fff748938fd5008d, /* 2298 */
128'he432854e05461c6396ca00d485330036, /* 2299 */
128'h85ca6622fc6fc0ef856685a2fcefc0ef, /* 2300 */
128'h080007932405ed298daad56ff0ef8526, /* 2301 */
128'hfa2fc0ef6fc5051300002517f8f41be3, /* 2302 */
128'h6aa66a4669e6790674a6856e744670e6, /* 2303 */
128'h808261096de27d027ca27c427be26b06, /* 2304 */
128'h85be00081363859a008bea6300167813, /* 2305 */
128'h85bafe081be385c6b7610605e10ce28c, /* 2306 */
128'h00002517892af0ca7119bf755dfdbfc5, /* 2307 */
128'hec6ef06af466fc5ee8d2ecce60c50513, /* 2308 */
128'he03289aef862e0dae4d6f4a6f8a2fc86, /* 2309 */
128'h2c975f2a0a1300002a17f2cfc0ef4b81, /* 2310 */
128'h4da1602d0d1300002d175fac8c930000, /* 2311 */
128'hc0ef85524401003b949b01779c334785, /* 2312 */
128'h4a93ef4fc0ef856685da00848b3bf00f, /* 2313 */
128'h974e00e908330036171367824601fffc, /* 2314 */
128'h856a85daed6fc0efe432855206f61063, /* 2315 */
128'h8b2ac5eff0ef854a85ce6622ecefc0ef, /* 2316 */
128'h040007932b85fbb41be38c562405e931, /* 2317 */
128'hea2fc0ef5fc5051300002517fafb90e3, /* 2318 */
128'h6aa66a4669e6790674a6855a744670e6, /* 2319 */
128'h808261096de27d027ca27c427be26b06, /* 2320 */
128'h00b83023e30c85d6e11185e200167513, /* 2321 */
128'hf4cef8cafca67175b7e95b7db7490605, /* 2322 */
128'he8daecd6f0d2698502000513892e84aa, /* 2323 */
128'he032f46ef86ae122e506fc66e0e2e4de, /* 2324 */
128'h138c0c1300003c174a01892ff0ef4a81, /* 2325 */
128'h8bca8b268f4c8c9300003c979c498993, /* 2326 */
128'h04fd956396da003d969367824d214d81, /* 2327 */
128'h0863ed45842aba2ff0ef852685ca866e, /* 2328 */
128'h8522df4fc0ef5765051300002517020a, /* 2329 */
128'h6b466ae67a0679a6794674e6640a60aa, /* 2330 */
128'h4a05808261497da27d427ce26c066ba6, /* 2331 */
128'he0ef842a90efe0efec36b7758ba68b4a, /* 2332 */
128'h67a28fcfe0efe42a902fe0efe82a908f, /* 2333 */
128'h15028c510106161b8d5d0105151b6642, /* 2334 */
128'h08a7bc23000037978d4166e291011402, /* 2335 */
128'h00fb86330006c683018786b34781e288, /* 2336 */
128'hf7b3ffa795e300d600230ff6f6930785, /* 2337 */
128'h001a879bfbdfe0ef4521ef910ba1033d, /* 2338 */
128'hfa9fe0ef0007c50397e68b8d00078a9b, /* 2339 */
128'hf0d2f4cef8ca7175bfa1547dbf0d0d85, /* 2340 */
128'he8daecd6fca66a050200051389ae892a, /* 2341 */
128'h8cb2f46ee122e506f86afc66e0e2e4de, /* 2342 */
128'h02048493000034974a81f73fe0ef4b01, /* 2343 */
128'h8c4e8bca7d4d0d1300002d179c4a0a13, /* 2344 */
128'h059d956397de00fc06b3003d97934d81, /* 2345 */
128'h8863e579842aa82ff0ef854a85ce866e, /* 2346 */
128'h8522cd4fc0ef4565051300002517020a, /* 2347 */
128'h6b466ae67a0679a6794674e6640a60aa, /* 2348 */
128'h4a85808261497da27d427ce26c066ba6, /* 2349 */
128'h842afedfd0efe836ec3eb7758c4a8bce, /* 2350 */
128'hfdbfd0efe02afe1fd0efe42afe7fd0ef, /* 2351 */
128'h8c518d590106161b0105151b67026622, /* 2352 */
128'hf8a7b023000037978d41910114021502, /* 2353 */
128'h902393c117c20004d783e38866c267e2, /* 2354 */
128'hd78300f6912393c117c20024d78300f6, /* 2355 */
128'h17c20064d78300f6922393c117c20044, /* 2356 */
128'he0ef4521ef91034df7b300f6932393c1, /* 2357 */
128'hc50397ea8b8d00078b1b001b079be87f, /* 2358 */
128'h6505b789547dbf290d85e73fe0ef0007, /* 2359 */
128'hfca6e122fff586138932f8ca71758082, /* 2360 */
128'h378505130000251785aa962a84ae842a, /* 2361 */
128'hf86afc66e0e2e4dee8daecd6f0d2f4ce, /* 2362 */
128'hd9930044d793bd8fc0efec36e506f46e, /* 2363 */
128'h44854a81e43e99a20034d793e83e0014, /* 2364 */
128'h360b8b9300002b97360b0b1300002b17, /* 2365 */
128'h360c8c9300002c97360c0c1300002c17, /* 2366 */
128'h368d8d9300002d97368d0d1300002d17, /* 2367 */
128'h0000251702997863e78a0a1300003a17, /* 2368 */
128'h74e68556640a60aab7afc0ef35c50513, /* 2369 */
128'h7ce26c066ba66b466ae67a0679a67946, /* 2370 */
128'hb52fc0ef855a85a6808261497da27d42, /* 2371 */
128'hc0ef8562b46fc0ef855e85ca00090663, /* 2372 */
128'hf0ef852265a2b38fc0ef856a85e6b40f, /* 2373 */
128'h6762010a2783b28fc0ef856eed15920f, /* 2374 */
128'h051300002517c58d000a358302f74963, /* 2375 */
128'h852285ce6642008a3783b0cfc0ef2de5, /* 2376 */
128'h4a89af4fc0ef2ce50513000025179782, /* 2377 */
128'h0485ae4fc0ef0865051300002517b7e9, /* 2378 */
128'hf022f4062bc50513000025177179bfa1, /* 2379 */
128'h251704000593c19fe0efe44ee84aec26, /* 2380 */
128'h051300002517ab8fc0ef2ba505130000, /* 2381 */
128'hc0ef2fa5051300002517aacfc0ef2d65, /* 2382 */
128'ha92fc0ef44850365051300002517aa0f, /* 2383 */
128'h46054685008495b3497901f499934441, /* 2384 */
128'h70a2ff2417e3e6dff0ef240501358533, /* 2385 */
128'h460580828082614569a2694264e27402, /* 2386 */
128'h45a901f61e1346814881470100c5131b, /* 2387 */
128'h0007802397aa000780234000081387f2, /* 2388 */
128'h97aa387d0007802397aa0007802397aa, /* 2389 */
128'h8e15c020267302b71d632705fe0813e3, /* 2390 */
128'h02a68733411686b33e800513c00026f3, /* 2391 */
128'h02a767b302b345bb02c7473340000593, /* 2392 */
128'h9f2fc06f294505130000251702a74733, /* 2393 */
128'h1141bf51c00028f3c02026f3fac710e3, /* 2394 */
128'h4509f75ff0ef4505f7bff0ef4501e406, /* 2395 */
128'hf63ff0ef4521f69ff0ef4511f6fff0ef, /* 2396 */
128'h400007b791011502bff1f5dff0ef4541, /* 2397 */
128'h07b7808225016388400007b78082e388, /* 2398 */
128'h400007b7808225016b880007b8234000, /* 2399 */
128'h0106161b8d5d0085979b808225017b88, /* 2400 */
128'h4000073747812581f7888d51400007b7, /* 2401 */
128'h8b097a98400006b73e80079300b7ef63, /* 2402 */
128'he60380827388400007b7ffe537fdc319, /* 2403 */
128'he406e0221141bfe1f710069127850006, /* 2404 */
128'h250135fd0045551b00b7d863842a4785, /* 2405 */
128'h943e20a7879300002797883dfebff0ef, /* 2406 */
128'h07b7a1ffe06f014160a2640200044503, /* 2407 */
128'h11010085151b67050185579b9d3d00b0, /* 2408 */
128'h842ec62ae8228fd90585651330070713, /* 2409 */
128'hf5bff0efec06c43e454d458946010034, /* 2410 */
128'h079385a2f4fff0ef454d460100344589, /* 2411 */
128'h058537e100d5802300f556b357610380, /* 2412 */
128'he0a2715d80826105644260e2fee79ae3, /* 2413 */
128'h8a2e84aae486ec56f052f44ef84afc26, /* 2414 */
128'h0144053b40000ab7ff86099b44018932, /* 2415 */
128'h16024089063bf79ff0ef002c03346663, /* 2416 */
128'h74e2640660a6ecbfd0ef92018526002c, /* 2417 */
128'hf0ef85a6808261616ae27a0279a27942, /* 2418 */
128'hb02304a19381178200c4579b2421f51f, /* 2419 */
128'he406ca250513000025171141bf6d00fa, /* 2420 */
128'hd3bf70eff88505130000051783efc0ef, /* 2421 */
128'h05130000251740a005b360a200055c63, /* 2422 */
128'hb4ffe06f014160a281afc06f0141c965, /* 2423 */
128'hfc067139957fe06f1a85051300002517, /* 2424 */
128'he0efe05ae456e852ec4ef04af426f822, /* 2425 */
128'h4401935fe0ef0e6505130000251790ff, /* 2426 */
128'h07b344950e49091300002917080009b7, /* 2427 */
128'hb0ef0405854a0004059b6390078e0134, /* 2428 */
128'h00002b174901da6f80effe9416e3fc1f, /* 2429 */
128'h0c0a8a9300002a97400004b7284b0b13, /* 2430 */
128'hc783016907b349910d0a0a1300002a17, /* 2431 */
128'h240125816080608ce09c090585560007, /* 2432 */
128'h25818552688c0004b823f7dfb0ef8622, /* 2433 */
128'h0054579b0ff47413fd391be3f6ffb0ef, /* 2434 */
128'h078a65a707130000071702f764634719, /* 2435 */
128'h0905051300002517878297ba439c97ba, /* 2436 */
128'h00002517a001aa9fe0ef8522f3ffb0ef, /* 2437 */
128'hb7f5edbff0ef8522f2bfb0ef08c50513, /* 2438 */
128'hc37ff0eff17fb0ef0885051300002517, /* 2439 */
128'h80eff05fb0ef0865051300002517bfe9, /* 2440 */
128'hef3fb0ef0845051300002517b7e1e14f, /* 2441 */
128'h00000000000000000000bf5dd0fff0ef, /* 2442 */
128'h00000000000000000000000000000000, /* 2443 */
128'h00000000000000000000000000000000, /* 2444 */
128'h00000000000000000000000000000000, /* 2445 */
128'h00000000000000000000000000000000, /* 2446 */
128'h00000000000000000000000000000000, /* 2447 */
128'h08082828282828080808080808080808, /* 2448 */
128'h08080808080808080808080808080808, /* 2449 */
128'h101010101010101010101010101010a0, /* 2450 */
128'h10101010101004040404040404040404, /* 2451 */
128'h01010101010101010141414141414110, /* 2452 */
128'h10101010100101010101010101010101, /* 2453 */
128'h02020202020202020242424242424210, /* 2454 */
128'h08101010100202020202020202020202, /* 2455 */
128'h00000000000000000000000000000000, /* 2456 */
128'h00000000000000000000000000000000, /* 2457 */
128'h101010101010101010101010101010a0, /* 2458 */
128'h10101010101010101010101010101010, /* 2459 */
128'h01010101010101010101010101010101, /* 2460 */
128'h02010101010101011001010101010101, /* 2461 */
128'h02020202020202020202020202020202, /* 2462 */
128'h02020202020202021002020202020202, /* 2463 */
128'hc1bdceee242070dbe8c7b756d76aa478, /* 2464 */
128'hfd469501a83046134787c62af57c0faf, /* 2465 */
128'h895cd7beffff5bb18b44f7af698098d8, /* 2466 */
128'h49b40821a679438efd9871936b901122, /* 2467 */
128'he9b6c7aa265e5a51c040b340f61e2562, /* 2468 */
128'he7d3fbc8d8a1e68102441453d62f105d, /* 2469 */
128'h455a14edf4d50d87c33707d621e1cde6, /* 2470 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /* 2471 */
128'hfde5380c6d9d61228771f681fffa3942, /* 2472 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /* 2473 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /* 2474 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /* 2475 */
128'hfc93a039ab9423a7432aff97f4292244, /* 2476 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /* 2477 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /* 2478 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /* 2479 */
128'h0c07020d08030e09040f0a05000b0601, /* 2480 */
128'h020f0c090603000d0a0704010e0b0805, /* 2481 */
128'h09020b040d060f08010a030c050e0700, /* 2482 */
128'h6c5f7465735f64735f63736972776f6c, /* 2483 */
128'h6e67696c615f64730000000000006465, /* 2484 */
128'h645f6b6c635f64730000000000000000, /* 2485 */
128'h69747465735f64730000000000007669, /* 2486 */
128'h735f646d635f6473000000000000676e, /* 2487 */
128'h74657365725f64730000000074726174, /* 2488 */
128'h6e636b6c625f64730000000000000000, /* 2489 */
128'h69736b6c625f64730000000000000074, /* 2490 */
128'h6f656d69745f6473000000000000657a, /* 2491 */
128'h655f7172695f64730000000000007475, /* 2492 */
128'h5f63736972776f6c000000000000006e, /* 2493 */
128'h00000000646d635f74726174735f6473, /* 2494 */
128'h746e695f746961775f63736972776f6c, /* 2495 */
128'h000000000067616c665f747075727265, /* 2496 */
128'h00007172695f64735f63736972776f6c, /* 2497 */
128'h695f646d635f64735f63736972776f6c, /* 2498 */
128'h5f63736972776f6c0000000000007172, /* 2499 */
128'h007172695f646e655f617461645f6473, /* 2500 */
128'h0000000087fe9c880000000087feaf50, /* 2501 */
128'h004c4b40004c4b400030000020000000, /* 2502 */
128'h6d6d5f6472616f62000000020000ffff, /* 2503 */
128'h0000000087fe4e920064637465675f63, /* 2504 */
128'h0000000087fe4cfe0000000087fe4aa0, /* 2505 */
128'h00000000000000000000000000000000, /* 2506 */
128'hffffbb74ffffbb70ffffbb70ffffbb4a, /* 2507 */
128'hffffbb78ffffbb78ffffbb78ffffbb78, /* 2508 */
128'h0000000087feb2780000000087feb268, /* 2509 */
128'h0000000087feb2a00000000087feb288, /* 2510 */
128'h0000000087feb2d00000000087feb2b8, /* 2511 */
128'h0000000087feb3000000000087feb2e8, /* 2512 */
128'h0000000087feb3300000000087feb318, /* 2513 */
128'h0000000087feb3600000000087feb348, /* 2514 */
128'h40040300400402004004010040040000, /* 2515 */
128'h40050000400405004004040140040400, /* 2516 */
128'h30000000000000030000000040050100, /* 2517 */
128'h60000000000000053000000000000001, /* 2518 */
128'h70000000000000027000000000000004, /* 2519 */
128'h00000001400000007000000000000000, /* 2520 */
128'h00000005000000012000000000000006, /* 2521 */
128'h20000000000000020000000040000000, /* 2522 */
128'h00000000100000000000000100000000, /* 2523 */
128'h1e19140f0d0c0a000000000000000000, /* 2524 */
128'h000186a00000271050463c37322d2823, /* 2525 */
128'h017d7840017d784000989680000f4240, /* 2526 */
128'h031975000319750002faf080018cba80, /* 2527 */
128'h02faf08005f5e10002faf080017d7840, /* 2528 */
128'h00000020000000000bebc2000c65d400, /* 2529 */
128'h00000200000001000000008000000040, /* 2530 */
128'h00002000000010000000080000000400, /* 2531 */
128'h0000c000000080000000600000004000, /* 2532 */
128'h37363534333231300002000000010000, /* 2533 */
128'h2043534952776f4c4645444342413938, /* 2534 */
128'h746f6f622d7520646573696d696e696d, /* 2535 */
128'h00000000647261432d445320726f6620, /* 2536 */
128'hfffff9cafffff9e0fffff9ccfffff9b8, /* 2537 */
128'h00000000fffffa04fffff9cafffff9f2, /* 2538 */
128'he00600003800000039080000edfe0dd0, /* 2539 */
128'h00000000100000001100000028000000, /* 2540 */
128'h0000000000000000a806000059010000, /* 2541 */
128'h00000000010000000000000000000000, /* 2542 */
128'h02000000000000000400000003000000, /* 2543 */
128'h020000000f0000000400000003000000, /* 2544 */
128'h2c6874651b0000001400000003000000, /* 2545 */
128'h007665642d657261622d656e61697261, /* 2546 */
128'h2c687465260000001000000003000000, /* 2547 */
128'h0100000000657261622d656e61697261, /* 2548 */
128'h1a0000000300000000006e65736f6863, /* 2549 */
128'h303140747261752f636f732f2c000000, /* 2550 */
128'h0000003030323531313a303030303030, /* 2551 */
128'h00000000737570630100000002000000, /* 2552 */
128'h01000000000000000400000003000000, /* 2553 */
128'h000000000f0000000400000003000000, /* 2554 */
128'h40787d01380000000400000003000000, /* 2555 */
128'h03000000000000304075706301000000, /* 2556 */
128'h0300000080f0fa024b00000004000000, /* 2557 */
128'h03000000007570635b00000004000000, /* 2558 */
128'h03000000000000006700000004000000, /* 2559 */
128'h0000000079616b6f6b00000005000000, /* 2560 */
128'h7a6874651b0000001300000003000000, /* 2561 */
128'h0000766373697200656e61697261202c, /* 2562 */
128'h34367672720000000b00000003000000, /* 2563 */
128'h0b000000030000000000636466616d69, /* 2564 */
128'h0000393376732c76637369727c000000, /* 2565 */
128'h01000000850000000000000003000000, /* 2566 */
128'h6f72746e6f632d747075727265746e69, /* 2567 */
128'h04000000030000000000000072656c6c, /* 2568 */
128'h0000000003000000010000008f000000, /* 2569 */
128'h1b0000000f00000003000000a0000000, /* 2570 */
128'h000063746e692d7570632c7663736972, /* 2571 */
128'h01000000b50000000400000003000000, /* 2572 */
128'h01000000bb0000000400000003000000, /* 2573 */
128'h01000000020000000200000002000000, /* 2574 */
128'h0030303030303030384079726f6d656d, /* 2575 */
128'h6f6d656d5b0000000700000003000000, /* 2576 */
128'h67000000100000000300000000007972, /* 2577 */
128'h00000008000000000000008000000000, /* 2578 */
128'h0300000000636f730100000002000000, /* 2579 */
128'h03000000020000000000000004000000, /* 2580 */
128'h03000000020000000f00000004000000, /* 2581 */
128'h616972612c6874651b0000001f000000, /* 2582 */
128'h706d697300636f732d657261622d656e, /* 2583 */
128'h000000000300000000007375622d656c, /* 2584 */
128'h303240746e696c6301000000c3000000, /* 2585 */
128'h0d000000030000000000003030303030, /* 2586 */
128'h30746e696c632c76637369721b000000, /* 2587 */
128'hca000000100000000300000000000000, /* 2588 */
128'h07000000010000000300000001000000, /* 2589 */
128'h00000000670000001000000003000000, /* 2590 */
128'h0300000000000c000000000000000002, /* 2591 */
128'h006c6f72746e6f63de00000008000000, /* 2592 */
128'h7075727265746e690100000002000000, /* 2593 */
128'h3030634072656c6c6f72746e6f632d74, /* 2594 */
128'h04000000030000000000000030303030, /* 2595 */
128'h04000000030000000000000000000000, /* 2596 */
128'h0c00000003000000010000008f000000, /* 2597 */
128'h003063696c702c76637369721b000000, /* 2598 */
128'h03000000a00000000000000003000000, /* 2599 */
128'h0b00000001000000ca00000010000000, /* 2600 */
128'h10000000030000000900000001000000, /* 2601 */
128'h000000000000000c0000000067000000, /* 2602 */
128'he8000000040000000300000000000004, /* 2603 */
128'hfb000000040000000300000007000000, /* 2604 */
128'hb5000000040000000300000003000000, /* 2605 */
128'hbb000000040000000300000002000000, /* 2606 */
128'h75626564010000000200000002000000, /* 2607 */
128'h0000304072656c6c6f72746e6f632d67, /* 2608 */
128'h637369721b0000001000000003000000, /* 2609 */
128'h03000000003331302d67756265642c76, /* 2610 */
128'hffff000001000000ca00000008000000, /* 2611 */
128'h00000000670000001000000003000000, /* 2612 */
128'h03000000001000000000000000000000, /* 2613 */
128'h006c6f72746e6f63de00000008000000, /* 2614 */
128'h30303140747261750100000002000000, /* 2615 */
128'h08000000030000000000003030303030, /* 2616 */
128'h03000000003035373631736e1b000000, /* 2617 */
128'h00000010000000006700000010000000, /* 2618 */
128'h04000000030000000010000000000000, /* 2619 */
128'h040000000300000080f0fa024b000000, /* 2620 */
128'h040000000300000000c2010006010000, /* 2621 */
128'h04000000030000000200000014010000, /* 2622 */
128'h04000000030000000100000025010000, /* 2623 */
128'h04000000030000000200000030010000, /* 2624 */
128'h0100000002000000040000003a010000, /* 2625 */
128'h3030303240636d6d2d63736972776f6c, /* 2626 */
128'h10000000030000000000000030303030, /* 2627 */
128'h00000000000000200000000067000000, /* 2628 */
128'h14010000040000000300000000000100, /* 2629 */
128'h25010000040000000300000002000000, /* 2630 */
128'h1b0000000c0000000300000002000000, /* 2631 */
128'h0200000000636d6d2d63736972776f6c, /* 2632 */
128'h406874652d63736972776f6c01000000, /* 2633 */
128'h03000000000000003030303030303033, /* 2634 */
128'h2d63736972776f6c1b0000000c000000, /* 2635 */
128'h5b000000080000000300000000687465, /* 2636 */
128'h0400000003000000006b726f7774656e, /* 2637 */
128'h04000000030000000200000014010000, /* 2638 */
128'h06000000030000000300000025010000, /* 2639 */
128'h0300000000007fe3023e180047010000, /* 2640 */
128'h00000030000000006700000010000000, /* 2641 */
128'h01000000020000000080000000000000, /* 2642 */
128'h303440646e7277682d63736972776f6c, /* 2643 */
128'h0e000000030000000000303030303030, /* 2644 */
128'h6e7277682d63736972776f6c1b000000, /* 2645 */
128'h67000000100000000300000000000064, /* 2646 */
128'h00100000000000000000004000000000, /* 2647 */
128'h09000000020000000200000002000000, /* 2648 */
128'h2300736c6c65632d7373657264646123, /* 2649 */
128'h61706d6f6300736c6c65632d657a6973, /* 2650 */
128'h6f647473006c65646f6d00656c626974, /* 2651 */
128'h65736162656d697400687461702d7475, /* 2652 */
128'h6b636f6c630079636e6575716572662d, /* 2653 */
128'h63697665640079636e6575716572662d, /* 2654 */
128'h75746174730067657200657079745f65, /* 2655 */
128'h2d756d6d006173692c76637369720073, /* 2656 */
128'h230074696c70732d626c740065707974, /* 2657 */
128'h00736c6c65632d747075727265746e69, /* 2658 */
128'h6f72746e6f632d747075727265746e69, /* 2659 */
128'h646e6168702c78756e696c0072656c6c, /* 2660 */
128'h727265746e69007365676e617200656c, /* 2661 */
128'h6572006465646e657478652d73747075, /* 2662 */
128'h616d2c76637369720073656d616e2d67, /* 2663 */
128'h766373697200797469726f6972702d78, /* 2664 */
128'h70732d746e6572727563007665646e2c, /* 2665 */
128'h61702d747075727265746e6900646565, /* 2666 */
128'h0073747075727265746e6900746e6572, /* 2667 */
128'h6f692d6765720074666968732d676572, /* 2668 */
128'h63616d2d6c61636f6c0068746469772d, /* 2669 */
128'h0000000000000000737365726464612d, /* 2670 */
128'h0000000000203a642520656369766544, /* 2671 */
128'h00203a6425206563697665642073250a, /* 2672 */
128'h00000000203a6425206563697665440a, /* 2673 */
128'h000a656369766564206e776f6e6b6e75, /* 2674 */
128'h00000a2973252c73252870756b6f6f6c, /* 2675 */
128'h7265206c616e7265746e692070636864, /* 2676 */
128'h00000000000000000a7025202c726f72, /* 2677 */
128'h5145525f5043484420676e69646e6553, /* 2678 */
128'h4b434120504348440000000a54534555, /* 2679 */
128'h696c432050434844000000000000000a, /* 2680 */
128'h203a7373657264644120504920746e65, /* 2681 */
128'h0000000a64252e64252e64252e642520, /* 2682 */
128'h73657264644120504920726576726553, /* 2683 */
128'h0a64252e64252e64252e642520203a73, /* 2684 */
128'h6120726574756f520000000000000000, /* 2685 */
128'h252e64252e642520203a737365726464, /* 2686 */
128'h6b73616d2074654e0000000a64252e64, /* 2687 */
128'h64252e642520203a7373657264646120, /* 2688 */
128'h697420657361654c000a64252e64252e, /* 2689 */
128'h7364253a6d64253a686425203d20656d, /* 2690 */
128'h3d206e69616d6f44000000000000000a, /* 2691 */
128'h4820746e65696c4300000a2273252220, /* 2692 */
128'h000a22732522203d20656d616e74736f, /* 2693 */
128'h000000000a44455050494b53204b4341, /* 2694 */
128'h000000000000000a4b414e2050434844, /* 2695 */
128'h73657264646120646574736575716552, /* 2696 */
128'h0000000000000a646573756665722073, /* 2697 */
128'h000000000000000a732520726f727245, /* 2698 */
128'h6e6f6974706f2064656c646e61686e75, /* 2699 */
128'h656c646e61686e55000000000a642520, /* 2700 */
128'h64252065646f63706f20504348442064, /* 2701 */
128'h20676e69646e6553000000000000000a, /* 2702 */
128'h000a595245564f435349445f50434844, /* 2703 */
128'h00000000000a29732528726f72726570, /* 2704 */
128'h3a2043414d2073250000000030687465, /* 2705 */
128'h3a583230253a583230253a5832302520, /* 2706 */
128'h000a583230253a583230253a58323025, /* 2707 */
128'h484420646e65732074276e646c756f43, /* 2708 */
128'h206e6f20595245564f43534944205043, /* 2709 */
128'h00000a7325203a732520656369766564, /* 2710 */
128'h5043484420726f6620676e6974696157, /* 2711 */
128'h2020202020202020000a524546464f5f, /* 2712 */
128'h00000000000063250000000000000020, /* 2713 */
128'h0000005832302520000000000000002e, /* 2714 */
128'h00000000732573250000000000000a0a, /* 2715 */
128'h00000000007325203a646c697542202c, /* 2716 */
128'h73257a4820756c250000000000007325, /* 2717 */
128'h0000000000756c250000000000000000, /* 2718 */
128'h0073257a4863252000000000646c252e, /* 2719 */
128'h00000000007325736574794220756c25, /* 2720 */
128'h00003a786c3830250073254269632520, /* 2721 */
128'h000a73252020202000786c6c2a302520, /* 2722 */
128'h000000203a5d64255b6e6f6974636553, /* 2723 */
128'h727265207974696e6173207264646170, /* 2724 */
128'h2c7825286e666c6500000a702520726f, /* 2725 */
128'h000000000a3b29782578302c78257830, /* 2726 */
128'h782578302c302c7825287465736d656d, /* 2727 */
128'h464f5f4f4c43414d00000000000a3b29, /* 2728 */
128'h464f5f494843414d0000000054455346, /* 2729 */
128'h46464f5f524c50540000000054455346, /* 2730 */
128'h46464f5f534346540000000000544553, /* 2731 */
128'h4c5254434f49444d0000000000544553, /* 2732 */
128'h46464f5f534346520054455346464f5f, /* 2733 */
128'h5346464f5f5253520000000000544553, /* 2734 */
128'h46464f5f444142520000000000005445, /* 2735 */
128'h46464f5f524c50520000000000544553, /* 2736 */
128'h000000003f3f3f3f0000000000544553, /* 2737 */
128'h000064252b54455346464f5f524c5052, /* 2738 */
128'h6f746f72502050490000000000000047, /* 2739 */
128'h00000000000000000a50495049203d20, /* 2740 */
128'h6f746f72502050490000000000000054, /* 2741 */
128'h6f746f7250205049000a504745203d20, /* 2742 */
128'h6165682074736574000a505550203d20, /* 2743 */
128'h6e6f6320747365740000000a3a726564, /* 2744 */
128'h6f746f7250205049000a3a73746e6574, /* 2745 */
128'h6f746f7250205049000a504449203d20, /* 2746 */
128'h6f746f725020504900000a5054203d20, /* 2747 */
128'h00000000000000000a50434344203d20, /* 2748 */
128'h6f746f72502050490000000000000036, /* 2749 */
128'h00000000000000000a50565352203d20, /* 2750 */
128'h000a455247203d206f746f7250205049, /* 2751 */
128'h000a505345203d206f746f7250205049, /* 2752 */
128'h00000a4841203d206f746f7250205049, /* 2753 */
128'h000a50544d203d206f746f7250205049, /* 2754 */
128'h5054454542203d206f746f7250205049, /* 2755 */
128'h6f746f72502050490000000000000a48, /* 2756 */
128'h000000000000000a5041434e45203d20, /* 2757 */
128'h6f746f7250205049000000000000004d, /* 2758 */
128'h00000000000000000a504d4f43203d20, /* 2759 */
128'h0a50544353203d206f746f7250205049, /* 2760 */
128'h6f746f72502050490000000000000000, /* 2761 */
128'h00000000000a4554494c504455203d20, /* 2762 */
128'h0a534c504d203d206f746f7250205049, /* 2763 */
128'h6f746f72502050490000000000000000, /* 2764 */
128'h6f746f7270205049000a574152203d20, /* 2765 */
128'h2820646574726f707075736e75203d20, /* 2766 */
128'h79745f6f746f7270000000000a297825, /* 2767 */
128'h0000000000000a78257830203d206570, /* 2768 */
128'h727265746e692064656c646e61686e75, /* 2769 */
128'h414d2070757465530000000a21747075, /* 2770 */
128'h4d454f2049505351000a726464612043, /* 2771 */
128'h0000000000000a7825203d205d64255b, /* 2772 */
128'h00000a786c253a786c25203d2043414d, /* 2773 */
128'h3025203d20737365726464612043414d, /* 2774 */
128'h3230253a783230253a783230253a7832, /* 2775 */
128'h0000000a2e783230253a783230253a78, /* 2776 */
128'h00007f7c5d5b3f3e3d3c3b3a2c2b2a22, /* 2777 */
128'h007f7c5d5b3f3e3d3c3b3a2e2c2b2a22, /* 2778 */
128'h66656463626139383736353433323130, /* 2779 */
128'h72776f6c2f6372730000000000000000, /* 2780 */
128'h00000000000000632e636d6d5f637369, /* 2781 */
128'h61625f6473203d3d20657361625f6473, /* 2782 */
128'h5f63736972776f6c00726464615f6573, /* 2783 */
128'h000a74756f656d6974207325203a6473, /* 2784 */
128'h616d202c6465766f6d65722064726143, /* 2785 */
128'h6425206f74206465676e616863206b73, /* 2786 */
128'h736e692064726143000000000000000a, /* 2787 */
128'h6e616863206b73616d202c6465747265, /* 2788 */
128'h0000000000000a6425206f7420646567, /* 2789 */
128'h25207461206465746165726320636d6d, /* 2790 */
128'h0000000a7825203d2074736f68202c78, /* 2791 */
128'h0000000000006f4e0000000000736559, /* 2792 */
128'h002020203a434d4d0000000052444420, /* 2793 */
128'h00000000000a7325203a656369766544, /* 2794 */
128'h3a4449207265727574636166756e614d, /* 2795 */
128'h0a7825203a4d454f000000000a782520, /* 2796 */
128'h6325203a656d614e0000000000000000, /* 2797 */
128'h0000000000000a206325632563256325, /* 2798 */
128'h00000a6425203a646565705320737542, /* 2799 */
128'h25203a79746963617061432068676948, /* 2800 */
128'h79746963617061430000000000000a73, /* 2801 */
128'h7464695720737542000000000000203a, /* 2802 */
128'h000000000a73257469622d6425203a68, /* 2803 */
128'h0000007825782520000000203a78250a, /* 2804 */
128'h00000000000064735f63736972776f6c, /* 2805 */
128'h0000000065646f6d206e776f6e6b6e55, /* 2806 */
128'h7830203a726f72724520737574617453, /* 2807 */
128'h2074756f656d69540000000a58383025, /* 2808 */
128'h616572206472616320676e6974696177, /* 2809 */
128'h6c69616620636d6d00000000000a7964, /* 2810 */
128'h6d6320706f747320646e6573206f7420, /* 2811 */
128'h6f6c62203a434d4d0000000000000a64, /* 2812 */
128'h20786c257830207265626d756e206b63, /* 2813 */
128'h6c2578302878616d2073646565637865, /* 2814 */
128'h203d3e20434d4d6500000000000a2978, /* 2815 */
128'h726f6620646572697571657220342e34, /* 2816 */
128'h642072657375206465636e61686e6520, /* 2817 */
128'h000000000000000a6165726120617461, /* 2818 */
128'h757320746f6e2073656f642064726143, /* 2819 */
128'h696e6f697469747261702074726f7070, /* 2820 */
128'h656f64206472614300000000000a676e, /* 2821 */
128'h20434820656e6966656420746f6e2073, /* 2822 */
128'h00000a657a69732070756f7267205057, /* 2823 */
128'h636e61686e6520617461642072657355, /* 2824 */
128'h5720434820746f6e2061657261206465, /* 2825 */
128'h696c6120657a69732070756f72672050, /* 2826 */
128'h72617020692550470000000a64656e67, /* 2827 */
128'h505720434820746f6e206e6f69746974, /* 2828 */
128'h67696c6120657a69732070756f726720, /* 2829 */
128'h656f642064726143000000000a64656e, /* 2830 */
128'h6e652074726f7070757320746f6e2073, /* 2831 */
128'h657475626972747461206465636e6168, /* 2832 */
128'h6e65206c61746f54000000000000000a, /* 2833 */
128'h6563786520657a6973206465636e6168, /* 2834 */
128'h20752528206d756d6978616d20736465, /* 2835 */
128'h656f64206472614300000a297525203e, /* 2836 */
128'h6f682074726f7070757320746f6e2073, /* 2837 */
128'h61702064656c6c6f72746e6f63207473, /* 2838 */
128'h6572206574697277206e6f6974697472, /* 2839 */
128'h6e6974746573207974696c696261696c, /* 2840 */
128'h726c61206472614300000000000a7367, /* 2841 */
128'h64656e6f697469747261702079646165, /* 2842 */
128'h206f6e203a434d4d000000000000000a, /* 2843 */
128'h0000000a746e65736572702064726163, /* 2844 */
128'h73657220746f6e206469642064726143, /* 2845 */
128'h20656761746c6f76206f7420646e6f70, /* 2846 */
128'h00000000000000000a217463656c6573, /* 2847 */
128'h7463656c6573206f7420656c62616e75, /* 2848 */
128'h00000000000000000a65646f6d206120, /* 2849 */
128'h646e756f66206473635f747865206f4e, /* 2850 */
128'h78363025206e614d0000000000000a21, /* 2851 */
128'h000000783430257834302520726e5320, /* 2852 */
128'h00000000632563256325632563256325, /* 2853 */
128'h6167656c20434d4d00000064252e6425, /* 2854 */
128'h636167654c2044530000000000007963, /* 2855 */
128'h6867694820434d4d0000000000000079, /* 2856 */
128'h0000297a484d36322820646565705320, /* 2857 */
128'h35282064656570532068676948204453, /* 2858 */
128'h6867694820434d4d000000297a484d30, /* 2859 */
128'h0000297a484d32352820646565705320, /* 2860 */
128'h7a484d32352820323552444420434d4d, /* 2861 */
128'h31524453205348550000000000000029, /* 2862 */
128'h00000000000000297a484d3532282032, /* 2863 */
128'h7a484d30352820353252445320534855, /* 2864 */
128'h35524453205348550000000000000029, /* 2865 */
128'h000000000000297a484d303031282030, /* 2866 */
128'h7a484d30352820303552444420534855, /* 2867 */
128'h31524453205348550000000000000029, /* 2868 */
128'h0000000000297a484d38303228203430, /* 2869 */
128'h0000297a484d30303228203030325348, /* 2870 */
128'h6f6e2064252065636976654420434d4d, /* 2871 */
128'h00000000000000000a646e756f662074, /* 2872 */
128'h000000000000445300000000434d4d65, /* 2873 */
128'h000000297325282000006425203a7325, /* 2874 */
128'h6e656c20656c69460000000000636d6d, /* 2875 */
128'h000000000000000a6425203d20687467, /* 2876 */
128'h0a7325203d202964252c70252835646d, /* 2877 */
128'h666c652064616f6c0000000000000000, /* 2878 */
128'h000a79726f6d656d20524444206f7420, /* 2879 */
128'h2064656c696166206461657220666c65, /* 2880 */
128'h000000646c252065646f632068746977, /* 2881 */
128'h6f6f7420687461702074736575716552, /* 2882 */
128'h00000000000a646c25202e676e6f6c20, /* 2883 */
128'h732522203a717277000000000000002f, /* 2884 */
128'h0a64253d657a69736b636f6c62202c22, /* 2885 */
128'h20657669656365520000000000000000, /* 2886 */
128'h0000000000000a2e646e6520656c6966, /* 2887 */
128'h656c6c6163207172775f656c646e6168, /* 2888 */
128'h206c6167656c6c4900000000000a2e64, /* 2889 */
128'h0a2e6e6f6974617265706f2050544654, /* 2890 */
128'h75716572206e656c0000000000000000, /* 2891 */
128'h6175746361202c5825203d2064657269, /* 2892 */
128'h000000005c2d2f7c000a7825203d206c, /* 2893 */
128'h20646564616f6c2065687420746f6f42, /* 2894 */
128'h6572646461207461206d6172676f7270, /* 2895 */
128'h000000000000000a2e2e2e7025207373, /* 2896 */
128'h445320746e756f6d206f74206c696146, /* 2897 */
128'h000000000000000a2172657669726420, /* 2898 */
128'h6e69206e69622e746f6f622064616f4c, /* 2899 */
128'h0000000000000a79726f6d656d206f74, /* 2900 */
128'h00000000000000006e69622e746f6f62, /* 2901 */
128'h62206e65706f206f742064656c696146, /* 2902 */
128'h206f74206c6961660000000a21746f6f, /* 2903 */
128'h000000000021656c69662065736f6c63, /* 2904 */
128'h6420746e756f6d75206f74206c696166, /* 2905 */
128'h20746f6f622d750a00000000216b7369, /* 2906 */
128'h67617473207473726966206465736162, /* 2907 */
128'h00000a726564616f6c20746f6f622065, /* 2908 */
128'h696166207325206e6f69747265737361, /* 2909 */
128'h696c202c732520656c6966202c64656c, /* 2910 */
128'h206e6f6974636e7566202c642520656e, /* 2911 */
128'h3a4552554c49414600000000000a7325, /* 2912 */
128'h74612078257830203d21207825783020, /* 2913 */
128'h00000a2e782578302074657366666f20, /* 2914 */
128'h7025203d203270202c7025203d203170, /* 2915 */
128'h2020202020202020000000000000000a, /* 2916 */
128'h08080808080808080000000000202020, /* 2917 */
128'h20676e69747465730000000000080808, /* 2918 */
128'h20676e69747365740000000000007525, /* 2919 */
128'h3a4552554c4941460000000000007525, /* 2920 */
128'h64612064616220656c626973736f7020, /* 2921 */
128'h666f20746120656e696c207373657264, /* 2922 */
128'h00000000000a2e782578302074657366, /* 2923 */
128'h7478656e206f7420676e697070696b53, /* 2924 */
128'h000000000000000a2e2e2e7473657420, /* 2925 */
128'h20202020200808080808080808080808, /* 2926 */
128'h08080808080808080808202020202020, /* 2927 */
128'h00000000000820080000000000000008, /* 2928 */
128'h78302073692065676e61722074736574, /* 2929 */
128'h00000000000a70257830206f74207025, /* 2930 */
128'h000000000075252f00752520706f6f4c, /* 2931 */
128'h6441206b637574530000000000000a3a, /* 2932 */
128'h0000203a732520200000007373657264, /* 2933 */
128'h00000a2e656e6f4400000000000a6b6f, /* 2934 */
128'h4d415244206c6174656d20657261420a, /* 2935 */
128'h65747365746d656d00000a7473657420, /* 2936 */
128'h20302e332e34206e6f69737265762072, /* 2937 */
128'h000000000000000a297469622d642528, /* 2938 */
128'h30322029432820746867697279706f43, /* 2939 */
128'h2073656c7261684320323130322d3130, /* 2940 */
128'h000000000000000a2e6e6f62617a6143, /* 2941 */
128'h74207265646e75206465736e6563694c, /* 2942 */
128'h50206c6172656e654720554e47206568, /* 2943 */
128'h65762065736e6563694c2063696c6275, /* 2944 */
128'h0a2e29796c6e6f282032206e6f697372, /* 2945 */
128'h5f676e696b726f770000000000000000, /* 2946 */
128'h20646c25202c424b6425203d20746573, /* 2947 */
128'h6c25202c736e6f697463757274736e69, /* 2948 */
128'h203d20495043202c73656c6379632064, /* 2949 */
128'h00000000000000000a646c252e646c25, /* 2950 */
128'h46454443424139383736353433323130, /* 2951 */
128'h6f57206f6c6c65480000000000000000, /* 2952 */
128'h205d64255b70777300000a0d21646c72, /* 2953 */
128'h73206863746977530000000a5825203d, /* 2954 */
128'h000a58252c5825203d20676e69747465, /* 2955 */
128'h5825203d2064656573206d6f646e6152, /* 2956 */
128'h0a746f6f62204453000000000000000a, /* 2957 */
128'h6f6f6220495053510000000000000000, /* 2958 */
128'h736574204d4152440000000000000a74, /* 2959 */
128'h6f6f6220505446540000000000000a74, /* 2960 */
128'h65742065686361430000000000000a74, /* 2961 */
128'h00000a0d7061727400000000000a7473, /* 2962 */
128'h00000002464c457fcccccccccccccccd, /* 2963 */
128'h1032547698badcfeefcdab8967452301, /* 2964 */
128'h5851f42d4c957f2d1000000020000000, /* 2965 */
128'haaaaaaaaaaaaaaaa5555555555555555, /* 2966 */
128'h00000000000000000000000000000000, /* 2967 */
128'h00000000000000000000000000000000, /* 2968 */
128'h00000000000000000000000000000000, /* 2969 */
128'h00000000000000000000000000000000, /* 2970 */
128'h00000000000000000000000000000000, /* 2971 */
128'h00000000000000000000000000000000, /* 2972 */
128'h00000000000000000000000000000000, /* 2973 */
128'h00000000000000000000000000000000, /* 2974 */
128'h00000000000000000000000000000000, /* 2975 */
128'h00004b4d47545045000000030f060301, /* 2976 */
128'h000000003000000000000000004b4d47, /* 2977 */
128'h00000000ffffffff0000000000000000, /* 2978 */
128'h0000646d635f6473000000000c000000, /* 2979 */
128'h00000000ffffffff00006772615f6473, /* 2980 */
128'h000000002f7c5c2d0000000087feb1f8, /* 2981 */
128'h000000060000000087feb3b0cc33aa55, /* 2982 */
128'h87fe708a0000000000000000ffffffff, /* 2983 */
128'h00000000000000000000000000000000, /* 2984 */
128'h00000000000000000000000000000000, /* 2985 */
128'h00000000000000000000000000000000, /* 2986 */
128'h00000000000000000000000000000000, /* 2987 */
128'h00000000000000000000000000000000, /* 2988 */
128'h00000000000000000000000000000000, /* 2989 */
128'h00000000000000000000000000000000, /* 2990 */
128'h00000000000000000000000000000000, /* 2991 */
128'h00000000000000000000000000000000, /* 2992 */
128'h00000000000000000000000000000000, /* 2993 */
128'h00000000000000000000000000000000, /* 2994 */
128'h00000000000000000000000000000000, /* 2995 */
128'h00000000000000000000000000000000, /* 2996 */
128'h00000000000000000000000000000000, /* 2997 */
128'h00000000000000000000000000000000, /* 2998 */
128'h00000000000000000000000000000000, /* 2999 */
128'h00000000000000000000000000000000, /* 3000 */
128'h00000000000000000000000000000000, /* 3001 */
128'h00000000000000000000000000000000, /* 3002 */
128'h00000000000000000000000000000000, /* 3003 */
128'h00000000000000000000000000000000, /* 3004 */
128'h00000000000000000000000000000000, /* 3005 */
128'h00000000000000000000000000000000, /* 3006 */
128'h00000000000000000000000000000000, /* 3007 */
128'h00000000000000000000000000000000, /* 3008 */
128'h00000000000000000000000000000000, /* 3009 */
128'h00000000000000000000000000000000, /* 3010 */
128'h00000000000000000000000000000000, /* 3011 */
128'h00000000000000000000000000000000, /* 3012 */
128'h00000000000000000000000000000000, /* 3013 */
128'h00000000000000000000000000000000, /* 3014 */
128'h00000000000000000000000000000000, /* 3015 */
128'h00000000000000000000000000000000, /* 3016 */
128'h00000000000000000000000000000000, /* 3017 */
128'h00000000000000000000000000000000, /* 3018 */
128'h00000000000000000000000000000000, /* 3019 */
128'h00000000000000000000000000000000, /* 3020 */
128'h00000000000000000000000000000000, /* 3021 */
128'h00000000000000000000000000000000, /* 3022 */
128'h00000000000000000000000000000000, /* 3023 */
128'h00000000000000000000000000000000, /* 3024 */
128'h00000000000000000000000000000000, /* 3025 */
128'h00000000000000000000000000000000, /* 3026 */
128'h00000000000000000000000000000000, /* 3027 */
128'h00000000000000000000000000000000, /* 3028 */
128'h00000000000000000000000000000000, /* 3029 */
128'h00000000000000000000000000000000, /* 3030 */
128'h00000000000000000000000000000000, /* 3031 */
128'h00000000000000000000000000000000, /* 3032 */
128'h00000000000000000000000000000000, /* 3033 */
128'h00000000000000000000000000000000, /* 3034 */
128'h00000000000000000000000000000000, /* 3035 */
128'h00000000000000000000000000000000, /* 3036 */
128'h00000000000000000000000000000000, /* 3037 */
128'h00000000000000000000000000000000, /* 3038 */
128'h00000000000000000000000000000000, /* 3039 */
128'h00000000000000000000000000000000, /* 3040 */
128'h00000000000000000000000000000000, /* 3041 */
128'h00000000000000000000000000000000, /* 3042 */
128'h00000000000000000000000000000000, /* 3043 */
128'h00000000000000000000000000000000, /* 3044 */
128'h00000000000000000000000000000000, /* 3045 */
128'h00000000000000000000000000000000, /* 3046 */
128'h00000000000000000000000000000000, /* 3047 */
128'h00000000000000000000000000000000, /* 3048 */
128'h00000000000000000000000000000000, /* 3049 */
128'h00000000000000000000000000000000, /* 3050 */
128'h00000000000000000000000000000000, /* 3051 */
128'h00000000000000000000000000000000, /* 3052 */
128'h00000000000000000000000000000000, /* 3053 */
128'h00000000000000000000000000000000, /* 3054 */
128'h00000000000000000000000000000000, /* 3055 */
128'h00000000000000000000000000000000, /* 3056 */
128'h00000000000000000000000000000000, /* 3057 */
128'h00000000000000000000000000000000, /* 3058 */
128'h00000000000000000000000000000000, /* 3059 */
128'h00000000000000000000000000000000, /* 3060 */
128'h00000000000000000000000000000000, /* 3061 */
128'h00000000000000000000000000000000, /* 3062 */
128'h00000000000000000000000000000000, /* 3063 */
128'h00000000000000000000000000000000, /* 3064 */
128'h00000000000000000000000000000000, /* 3065 */
128'h00000000000000000000000000000000, /* 3066 */
128'h00000000000000000000000000000000, /* 3067 */
128'h00000000000000000000000000000000, /* 3068 */
128'h00000000000000000000000000000000, /* 3069 */
128'h00000000000000000000000000000000, /* 3070 */
128'h00000000000000000000000000000000, /* 3071 */
128'h00000000000000000000000000000000, /* 3072 */
128'h00000000000000000000000000000000, /* 3073 */
128'h00000000000000000000000000000000, /* 3074 */
128'h00000000000000000000000000000000, /* 3075 */
128'h00000000000000000000000000000000, /* 3076 */
128'h00000000000000000000000000000000, /* 3077 */
128'h00000000000000000000000000000000, /* 3078 */
128'h00000000000000000000000000000000, /* 3079 */
128'h00000000000000000000000000000000, /* 3080 */
128'h00000000000000000000000000000000, /* 3081 */
128'h00000000000000000000000000000000, /* 3082 */
128'h00000000000000000000000000000000, /* 3083 */
128'h00000000000000000000000000000000, /* 3084 */
128'h00000000000000000000000000000000, /* 3085 */
128'h00000000000000000000000000000000, /* 3086 */
128'h00000000000000000000000000000000, /* 3087 */
128'h00000000000000000000000000000000, /* 3088 */
128'h00000000000000000000000000000000, /* 3089 */
128'h00000000000000000000000000000000, /* 3090 */
128'h00000000000000000000000000000000, /* 3091 */
128'h00000000000000000000000000000000, /* 3092 */
128'h00000000000000000000000000000000, /* 3093 */
128'h00000000000000000000000000000000, /* 3094 */
128'h00000000000000000000000000000000, /* 3095 */
128'h00000000000000000000000000000000, /* 3096 */
128'h00000000000000000000000000000000, /* 3097 */
128'h00000000000000000000000000000000, /* 3098 */
128'h00000000000000000000000000000000, /* 3099 */
128'h00000000000000000000000000000000, /* 3100 */
128'h00000000000000000000000000000000, /* 3101 */
128'h00000000000000000000000000000000, /* 3102 */
128'h00000000000000000000000000000000, /* 3103 */
128'h00000000000000000000000000000000, /* 3104 */
128'h00000000000000000000000000000000, /* 3105 */
128'h00000000000000000000000000000000, /* 3106 */
128'h00000000000000000000000000000000, /* 3107 */
128'h00000000000000000000000000000000, /* 3108 */
128'h00000000000000000000000000000000, /* 3109 */
128'h00000000000000000000000000000000, /* 3110 */
128'h00000000000000000000000000000000, /* 3111 */
128'h00000000000000000000000000000000, /* 3112 */
128'h00000000000000000000000000000000, /* 3113 */
128'h00000000000000000000000000000000, /* 3114 */
128'h00000000000000000000000000000000, /* 3115 */
128'h00000000000000000000000000000000, /* 3116 */
128'h00000000000000000000000000000000, /* 3117 */
128'h00000000000000000000000000000000, /* 3118 */
128'h00000000000000000000000000000000, /* 3119 */
128'h00000000000000000000000000000000, /* 3120 */
128'h00000000000000000000000000000000, /* 3121 */
128'h00000000000000000000000000000000, /* 3122 */
128'h00000000000000000000000000000000, /* 3123 */
128'h00000000000000000000000000000000, /* 3124 */
128'h00000000000000000000000000000000, /* 3125 */
128'h00000000000000000000000000000000, /* 3126 */
128'h00000000000000000000000000000000, /* 3127 */
128'h00000000000000000000000000000000, /* 3128 */
128'h00000000000000000000000000000000, /* 3129 */
128'h00000000000000000000000000000000, /* 3130 */
128'h00000000000000000000000000000000, /* 3131 */
128'h00000000000000000000000000000000, /* 3132 */
128'h00000000000000000000000000000000, /* 3133 */
128'h00000000000000000000000000000000, /* 3134 */
128'h00000000000000000000000000000000, /* 3135 */
128'h00000000000000000000000000000000, /* 3136 */
128'h00000000000000000000000000000000, /* 3137 */
128'h00000000000000000000000000000000, /* 3138 */
128'h00000000000000000000000000000000, /* 3139 */
128'h00000000000000000000000000000000, /* 3140 */
128'h00000000000000000000000000000000, /* 3141 */
128'h00000000000000000000000000000000, /* 3142 */
128'h00000000000000000000000000000000, /* 3143 */
128'h00000000000000000000000000000000, /* 3144 */
128'h00000000000000000000000000000000, /* 3145 */
128'h00000000000000000000000000000000, /* 3146 */
128'h00000000000000000000000000000000, /* 3147 */
128'h00000000000000000000000000000000, /* 3148 */
128'h00000000000000000000000000000000, /* 3149 */
128'h00000000000000000000000000000000, /* 3150 */
128'h00000000000000000000000000000000, /* 3151 */
128'h00000000000000000000000000000000, /* 3152 */
128'h00000000000000000000000000000000, /* 3153 */
128'h00000000000000000000000000000000, /* 3154 */
128'h00000000000000000000000000000000, /* 3155 */
128'h00000000000000000000000000000000, /* 3156 */
128'h00000000000000000000000000000000, /* 3157 */
128'h00000000000000000000000000000000, /* 3158 */
128'h00000000000000000000000000000000, /* 3159 */
128'h00000000000000000000000000000000, /* 3160 */
128'h00000000000000000000000000000000, /* 3161 */
128'h00000000000000000000000000000000, /* 3162 */
128'h00000000000000000000000000000000, /* 3163 */
128'h00000000000000000000000000000000, /* 3164 */
128'h00000000000000000000000000000000, /* 3165 */
128'h00000000000000000000000000000000, /* 3166 */
128'h00000000000000000000000000000000, /* 3167 */
128'h00000000000000000000000000000000, /* 3168 */
128'h00000000000000000000000000000000, /* 3169 */
128'h00000000000000000000000000000000, /* 3170 */
128'h00000000000000000000000000000000, /* 3171 */
128'h00000000000000000000000000000000, /* 3172 */
128'h00000000000000000000000000000000, /* 3173 */
128'h00000000000000000000000000000000, /* 3174 */
128'h00000000000000000000000000000000, /* 3175 */
128'h00000000000000000000000000000000, /* 3176 */
128'h00000000000000000000000000000000, /* 3177 */
128'h00000000000000000000000000000000, /* 3178 */
128'h00000000000000000000000000000000, /* 3179 */
128'h00000000000000000000000000000000, /* 3180 */
128'h00000000000000000000000000000000, /* 3181 */
128'h00000000000000000000000000000000, /* 3182 */
128'h00000000000000000000000000000000, /* 3183 */
128'h00000000000000000000000000000000, /* 3184 */
128'h00000000000000000000000000000000, /* 3185 */
128'h00000000000000000000000000000000, /* 3186 */
128'h00000000000000000000000000000000, /* 3187 */
128'h00000000000000000000000000000000, /* 3188 */
128'h00000000000000000000000000000000, /* 3189 */
128'h00000000000000000000000000000000, /* 3190 */
128'h00000000000000000000000000000000, /* 3191 */
128'h00000000000000000000000000000000, /* 3192 */
128'h00000000000000000000000000000000, /* 3193 */
128'h00000000000000000000000000000000, /* 3194 */
128'h00000000000000000000000000000000, /* 3195 */
128'h00000000000000000000000000000000, /* 3196 */
128'h00000000000000000000000000000000, /* 3197 */
128'h00000000000000000000000000000000, /* 3198 */
128'h00000000000000000000000000000000, /* 3199 */
128'h00000000000000000000000000000000, /* 3200 */
128'h00000000000000000000000000000000, /* 3201 */
128'h00000000000000000000000000000000, /* 3202 */
128'h00000000000000000000000000000000, /* 3203 */
128'h00000000000000000000000000000000, /* 3204 */
128'h00000000000000000000000000000000, /* 3205 */
128'h00000000000000000000000000000000, /* 3206 */
128'h00000000000000000000000000000000, /* 3207 */
128'h00000000000000000000000000000000, /* 3208 */
128'h00000000000000000000000000000000, /* 3209 */
128'h00000000000000000000000000000000, /* 3210 */
128'h00000000000000000000000000000000, /* 3211 */
128'h00000000000000000000000000000000, /* 3212 */
128'h00000000000000000000000000000000, /* 3213 */
128'h00000000000000000000000000000000, /* 3214 */
128'h00000000000000000000000000000000, /* 3215 */
128'h00000000000000000000000000000000, /* 3216 */
128'h00000000000000000000000000000000, /* 3217 */
128'h00000000000000000000000000000000, /* 3218 */
128'h00000000000000000000000000000000, /* 3219 */
128'h00000000000000000000000000000000, /* 3220 */
128'h00000000000000000000000000000000, /* 3221 */
128'h00000000000000000000000000000000, /* 3222 */
128'h00000000000000000000000000000000, /* 3223 */
128'h00000000000000000000000000000000, /* 3224 */
128'h00000000000000000000000000000000, /* 3225 */
128'h00000000000000000000000000000000, /* 3226 */
128'h00000000000000000000000000000000, /* 3227 */
128'h00000000000000000000000000000000, /* 3228 */
128'h00000000000000000000000000000000, /* 3229 */
128'h00000000000000000000000000000000, /* 3230 */
128'h00000000000000000000000000000000, /* 3231 */
128'h00000000000000000000000000000000, /* 3232 */
128'h00000000000000000000000000000000, /* 3233 */
128'h00000000000000000000000000000000, /* 3234 */
128'h00000000000000000000000000000000, /* 3235 */
128'h00000000000000000000000000000000, /* 3236 */
128'h00000000000000000000000000000000, /* 3237 */
128'h00000000000000000000000000000000, /* 3238 */
128'h00000000000000000000000000000000, /* 3239 */
128'h00000000000000000000000000000000, /* 3240 */
128'h00000000000000000000000000000000, /* 3241 */
128'h00000000000000000000000000000000, /* 3242 */
128'h00000000000000000000000000000000, /* 3243 */
128'h00000000000000000000000000000000, /* 3244 */
128'h00000000000000000000000000000000, /* 3245 */
128'h00000000000000000000000000000000, /* 3246 */
128'h00000000000000000000000000000000, /* 3247 */
128'h00000000000000000000000000000000, /* 3248 */
128'h00000000000000000000000000000000, /* 3249 */
128'h00000000000000000000000000000000, /* 3250 */
128'h00000000000000000000000000000000, /* 3251 */
128'h00000000000000000000000000000000, /* 3252 */
128'h00000000000000000000000000000000, /* 3253 */
128'h00000000000000000000000000000000, /* 3254 */
128'h00000000000000000000000000000000, /* 3255 */
128'h00000000000000000000000000000000, /* 3256 */
128'h00000000000000000000000000000000, /* 3257 */
128'h00000000000000000000000000000000, /* 3258 */
128'h00000000000000000000000000000000, /* 3259 */
128'h00000000000000000000000000000000, /* 3260 */
128'h00000000000000000000000000000000, /* 3261 */
128'h00000000000000000000000000000000, /* 3262 */
128'h00000000000000000000000000000000, /* 3263 */
128'h00000000000000000000000000000000, /* 3264 */
128'h00000000000000000000000000000000, /* 3265 */
128'h00000000000000000000000000000000, /* 3266 */
128'h00000000000000000000000000000000, /* 3267 */
128'h00000000000000000000000000000000, /* 3268 */
128'h00000000000000000000000000000000, /* 3269 */
128'h00000000000000000000000000000000, /* 3270 */
128'h00000000000000000000000000000000, /* 3271 */
128'h00000000000000000000000000000000, /* 3272 */
128'h00000000000000000000000000000000, /* 3273 */
128'h00000000000000000000000000000000, /* 3274 */
128'h00000000000000000000000000000000, /* 3275 */
128'h00000000000000000000000000000000, /* 3276 */
128'h00000000000000000000000000000000, /* 3277 */
128'h00000000000000000000000000000000, /* 3278 */
128'h00000000000000000000000000000000, /* 3279 */
128'h00000000000000000000000000000000, /* 3280 */
128'h00000000000000000000000000000000, /* 3281 */
128'h00000000000000000000000000000000, /* 3282 */
128'h00000000000000000000000000000000, /* 3283 */
128'h00000000000000000000000000000000, /* 3284 */
128'h00000000000000000000000000000000, /* 3285 */
128'h00000000000000000000000000000000, /* 3286 */
128'h00000000000000000000000000000000, /* 3287 */
128'h00000000000000000000000000000000, /* 3288 */
128'h00000000000000000000000000000000, /* 3289 */
128'h00000000000000000000000000000000, /* 3290 */
128'h00000000000000000000000000000000, /* 3291 */
128'h00000000000000000000000000000000, /* 3292 */
128'h00000000000000000000000000000000, /* 3293 */
128'h00000000000000000000000000000000, /* 3294 */
128'h00000000000000000000000000000000, /* 3295 */
128'h00000000000000000000000000000000, /* 3296 */
128'h00000000000000000000000000000000, /* 3297 */
128'h00000000000000000000000000000000, /* 3298 */
128'h00000000000000000000000000000000, /* 3299 */
128'h00000000000000000000000000000000, /* 3300 */
128'h00000000000000000000000000000000, /* 3301 */
128'h00000000000000000000000000000000, /* 3302 */
128'h00000000000000000000000000000000, /* 3303 */
128'h00000000000000000000000000000000, /* 3304 */
128'h00000000000000000000000000000000, /* 3305 */
128'h00000000000000000000000000000000, /* 3306 */
128'h00000000000000000000000000000000, /* 3307 */
128'h00000000000000000000000000000000, /* 3308 */
128'h00000000000000000000000000000000, /* 3309 */
128'h00000000000000000000000000000000, /* 3310 */
128'h00000000000000000000000000000000, /* 3311 */
128'h00000000000000000000000000000000, /* 3312 */
128'h00000000000000000000000000000000, /* 3313 */
128'h00000000000000000000000000000000, /* 3314 */
128'h00000000000000000000000000000000, /* 3315 */
128'h00000000000000000000000000000000, /* 3316 */
128'h00000000000000000000000000000000, /* 3317 */
128'h00000000000000000000000000000000, /* 3318 */
128'h00000000000000000000000000000000, /* 3319 */
128'h00000000000000000000000000000000, /* 3320 */
128'h00000000000000000000000000000000, /* 3321 */
128'h00000000000000000000000000000000, /* 3322 */
128'h00000000000000000000000000000000, /* 3323 */
128'h00000000000000000000000000000000, /* 3324 */
128'h00000000000000000000000000000000, /* 3325 */
128'h00000000000000000000000000000000, /* 3326 */
128'h00000000000000000000000000000000, /* 3327 */
128'h00000000000000000000000000000000, /* 3328 */
128'h00000000000000000000000000000000, /* 3329 */
128'h00000000000000000000000000000000, /* 3330 */
128'h00000000000000000000000000000000, /* 3331 */
128'h00000000000000000000000000000000, /* 3332 */
128'h00000000000000000000000000000000, /* 3333 */
128'h00000000000000000000000000000000, /* 3334 */
128'h00000000000000000000000000000000, /* 3335 */
128'h00000000000000000000000000000000, /* 3336 */
128'h00000000000000000000000000000000, /* 3337 */
128'h00000000000000000000000000000000, /* 3338 */
128'h00000000000000000000000000000000, /* 3339 */
128'h00000000000000000000000000000000, /* 3340 */
128'h00000000000000000000000000000000, /* 3341 */
128'h00000000000000000000000000000000, /* 3342 */
128'h00000000000000000000000000000000, /* 3343 */
128'h00000000000000000000000000000000, /* 3344 */
128'h00000000000000000000000000000000, /* 3345 */
128'h00000000000000000000000000000000, /* 3346 */
128'h00000000000000000000000000000000, /* 3347 */
128'h00000000000000000000000000000000, /* 3348 */
128'h00000000000000000000000000000000, /* 3349 */
128'h00000000000000000000000000000000, /* 3350 */
128'h00000000000000000000000000000000, /* 3351 */
128'h00000000000000000000000000000000, /* 3352 */
128'h00000000000000000000000000000000, /* 3353 */
128'h00000000000000000000000000000000, /* 3354 */
128'h00000000000000000000000000000000, /* 3355 */
128'h00000000000000000000000000000000, /* 3356 */
128'h00000000000000000000000000000000, /* 3357 */
128'h00000000000000000000000000000000, /* 3358 */
128'h00000000000000000000000000000000, /* 3359 */
128'h00000000000000000000000000000000, /* 3360 */
128'h00000000000000000000000000000000, /* 3361 */
128'h00000000000000000000000000000000, /* 3362 */
128'h00000000000000000000000000000000, /* 3363 */
128'h00000000000000000000000000000000, /* 3364 */
128'h00000000000000000000000000000000, /* 3365 */
128'h00000000000000000000000000000000, /* 3366 */
128'h00000000000000000000000000000000, /* 3367 */
128'h00000000000000000000000000000000, /* 3368 */
128'h00000000000000000000000000000000, /* 3369 */
128'h00000000000000000000000000000000, /* 3370 */
128'h00000000000000000000000000000000, /* 3371 */
128'h00000000000000000000000000000000, /* 3372 */
128'h00000000000000000000000000000000, /* 3373 */
128'h00000000000000000000000000000000, /* 3374 */
128'h00000000000000000000000000000000, /* 3375 */
128'h00000000000000000000000000000000, /* 3376 */
128'h00000000000000000000000000000000, /* 3377 */
128'h00000000000000000000000000000000, /* 3378 */
128'h00000000000000000000000000000000, /* 3379 */
128'h00000000000000000000000000000000, /* 3380 */
128'h00000000000000000000000000000000, /* 3381 */
128'h00000000000000000000000000000000, /* 3382 */
128'h00000000000000000000000000000000, /* 3383 */
128'h00000000000000000000000000000000, /* 3384 */
128'h00000000000000000000000000000000, /* 3385 */
128'h00000000000000000000000000000000, /* 3386 */
128'h00000000000000000000000000000000, /* 3387 */
128'h00000000000000000000000000000000, /* 3388 */
128'h00000000000000000000000000000000, /* 3389 */
128'h00000000000000000000000000000000, /* 3390 */
128'h00000000000000000000000000000000, /* 3391 */
128'h00000000000000000000000000000000, /* 3392 */
128'h00000000000000000000000000000000, /* 3393 */
128'h00000000000000000000000000000000, /* 3394 */
128'h00000000000000000000000000000000, /* 3395 */
128'h00000000000000000000000000000000, /* 3396 */
128'h00000000000000000000000000000000, /* 3397 */
128'h00000000000000000000000000000000, /* 3398 */
128'h00000000000000000000000000000000, /* 3399 */
128'h00000000000000000000000000000000, /* 3400 */
128'h00000000000000000000000000000000, /* 3401 */
128'h00000000000000000000000000000000, /* 3402 */
128'h00000000000000000000000000000000, /* 3403 */
128'h00000000000000000000000000000000, /* 3404 */
128'h00000000000000000000000000000000, /* 3405 */
128'h00000000000000000000000000000000, /* 3406 */
128'h00000000000000000000000000000000, /* 3407 */
128'h00000000000000000000000000000000, /* 3408 */
128'h00000000000000000000000000000000, /* 3409 */
128'h00000000000000000000000000000000, /* 3410 */
128'h00000000000000000000000000000000, /* 3411 */
128'h00000000000000000000000000000000, /* 3412 */
128'h00000000000000000000000000000000, /* 3413 */
128'h00000000000000000000000000000000, /* 3414 */
128'h00000000000000000000000000000000, /* 3415 */
128'h00000000000000000000000000000000, /* 3416 */
128'h00000000000000000000000000000000, /* 3417 */
128'h00000000000000000000000000000000, /* 3418 */
128'h00000000000000000000000000000000, /* 3419 */
128'h00000000000000000000000000000000, /* 3420 */
128'h00000000000000000000000000000000, /* 3421 */
128'h00000000000000000000000000000000, /* 3422 */
128'h00000000000000000000000000000000, /* 3423 */
128'h00000000000000000000000000000000, /* 3424 */
128'h00000000000000000000000000000000, /* 3425 */
128'h00000000000000000000000000000000, /* 3426 */
128'h00000000000000000000000000000000, /* 3427 */
128'h00000000000000000000000000000000, /* 3428 */
128'h00000000000000000000000000000000, /* 3429 */
128'h00000000000000000000000000000000, /* 3430 */
128'h00000000000000000000000000000000, /* 3431 */
128'h00000000000000000000000000000000, /* 3432 */
128'h00000000000000000000000000000000, /* 3433 */
128'h00000000000000000000000000000000, /* 3434 */
128'h00000000000000000000000000000000, /* 3435 */
128'h00000000000000000000000000000000, /* 3436 */
128'h00000000000000000000000000000000, /* 3437 */
128'h00000000000000000000000000000000, /* 3438 */
128'h00000000000000000000000000000000, /* 3439 */
128'h00000000000000000000000000000000, /* 3440 */
128'h00000000000000000000000000000000, /* 3441 */
128'h00000000000000000000000000000000, /* 3442 */
128'h00000000000000000000000000000000, /* 3443 */
128'h00000000000000000000000000000000, /* 3444 */
128'h00000000000000000000000000000000, /* 3445 */
128'h00000000000000000000000000000000, /* 3446 */
128'h00000000000000000000000000000000, /* 3447 */
128'h00000000000000000000000000000000, /* 3448 */
128'h00000000000000000000000000000000, /* 3449 */
128'h00000000000000000000000000000000, /* 3450 */
128'h00000000000000000000000000000000, /* 3451 */
128'h00000000000000000000000000000000, /* 3452 */
128'h00000000000000000000000000000000, /* 3453 */
128'h00000000000000000000000000000000, /* 3454 */
128'h00000000000000000000000000000000, /* 3455 */
128'h00000000000000000000000000000000, /* 3456 */
128'h00000000000000000000000000000000, /* 3457 */
128'h00000000000000000000000000000000, /* 3458 */
128'h00000000000000000000000000000000, /* 3459 */
128'h00000000000000000000000000000000, /* 3460 */
128'h00000000000000000000000000000000, /* 3461 */
128'h00000000000000000000000000000000, /* 3462 */
128'h00000000000000000000000000000000, /* 3463 */
128'h00000000000000000000000000000000, /* 3464 */
128'h00000000000000000000000000000000, /* 3465 */
128'h00000000000000000000000000000000, /* 3466 */
128'h00000000000000000000000000000000, /* 3467 */
128'h00000000000000000000000000000000, /* 3468 */
128'h00000000000000000000000000000000, /* 3469 */
128'h00000000000000000000000000000000, /* 3470 */
128'h00000000000000000000000000000000, /* 3471 */
128'h00000000000000000000000000000000, /* 3472 */
128'h00000000000000000000000000000000, /* 3473 */
128'h00000000000000000000000000000000, /* 3474 */
128'h00000000000000000000000000000000, /* 3475 */
128'h00000000000000000000000000000000, /* 3476 */
128'h00000000000000000000000000000000, /* 3477 */
128'h00000000000000000000000000000000, /* 3478 */
128'h00000000000000000000000000000000, /* 3479 */
128'h00000000000000000000000000000000, /* 3480 */
128'h00000000000000000000000000000000, /* 3481 */
128'h00000000000000000000000000000000, /* 3482 */
128'h00000000000000000000000000000000, /* 3483 */
128'h00000000000000000000000000000000, /* 3484 */
128'h00000000000000000000000000000000, /* 3485 */
128'h00000000000000000000000000000000, /* 3486 */
128'h00000000000000000000000000000000, /* 3487 */
128'h00000000000000000000000000000000, /* 3488 */
128'h00000000000000000000000000000000, /* 3489 */
128'h00000000000000000000000000000000, /* 3490 */
128'h00000000000000000000000000000000, /* 3491 */
128'h00000000000000000000000000000000, /* 3492 */
128'h00000000000000000000000000000000, /* 3493 */
128'h00000000000000000000000000000000, /* 3494 */
128'h00000000000000000000000000000000, /* 3495 */
128'h00000000000000000000000000000000, /* 3496 */
128'h00000000000000000000000000000000, /* 3497 */
128'h00000000000000000000000000000000, /* 3498 */
128'h00000000000000000000000000000000, /* 3499 */
128'h00000000000000000000000000000000, /* 3500 */
128'h00000000000000000000000000000000, /* 3501 */
128'h00000000000000000000000000000000, /* 3502 */
128'h00000000000000000000000000000000, /* 3503 */
128'h00000000000000000000000000000000, /* 3504 */
128'h00000000000000000000000000000000, /* 3505 */
128'h00000000000000000000000000000000, /* 3506 */
128'h00000000000000000000000000000000, /* 3507 */
128'h00000000000000000000000000000000, /* 3508 */
128'h00000000000000000000000000000000, /* 3509 */
128'h00000000000000000000000000000000, /* 3510 */
128'h00000000000000000000000000000000, /* 3511 */
128'h00000000000000000000000000000000, /* 3512 */
128'h00000000000000000000000000000000, /* 3513 */
128'h00000000000000000000000000000000, /* 3514 */
128'h00000000000000000000000000000000, /* 3515 */
128'h00000000000000000000000000000000, /* 3516 */
128'h00000000000000000000000000000000, /* 3517 */
128'h00000000000000000000000000000000, /* 3518 */
128'h00000000000000000000000000000000, /* 3519 */
128'h00000000000000000000000000000000, /* 3520 */
128'h00000000000000000000000000000000, /* 3521 */
128'h00000000000000000000000000000000, /* 3522 */
128'h00000000000000000000000000000000, /* 3523 */
128'h00000000000000000000000000000000, /* 3524 */
128'h00000000000000000000000000000000, /* 3525 */
128'h00000000000000000000000000000000, /* 3526 */
128'h00000000000000000000000000000000, /* 3527 */
128'h00000000000000000000000000000000, /* 3528 */
128'h00000000000000000000000000000000, /* 3529 */
128'h00000000000000000000000000000000, /* 3530 */
128'h00000000000000000000000000000000, /* 3531 */
128'h00000000000000000000000000000000, /* 3532 */
128'h00000000000000000000000000000000, /* 3533 */
128'h00000000000000000000000000000000, /* 3534 */
128'h00000000000000000000000000000000, /* 3535 */
128'h00000000000000000000000000000000, /* 3536 */
128'h00000000000000000000000000000000, /* 3537 */
128'h00000000000000000000000000000000, /* 3538 */
128'h00000000000000000000000000000000, /* 3539 */
128'h00000000000000000000000000000000, /* 3540 */
128'h00000000000000000000000000000000, /* 3541 */
128'h00000000000000000000000000000000, /* 3542 */
128'h00000000000000000000000000000000, /* 3543 */
128'h00000000000000000000000000000000, /* 3544 */
128'h00000000000000000000000000000000, /* 3545 */
128'h00000000000000000000000000000000, /* 3546 */
128'h00000000000000000000000000000000, /* 3547 */
128'h00000000000000000000000000000000, /* 3548 */
128'h00000000000000000000000000000000, /* 3549 */
128'h00000000000000000000000000000000, /* 3550 */
128'h00000000000000000000000000000000, /* 3551 */
128'h00000000000000000000000000000000, /* 3552 */
128'h00000000000000000000000000000000, /* 3553 */
128'h00000000000000000000000000000000, /* 3554 */
128'h00000000000000000000000000000000, /* 3555 */
128'h00000000000000000000000000000000, /* 3556 */
128'h00000000000000000000000000000000, /* 3557 */
128'h00000000000000000000000000000000, /* 3558 */
128'h00000000000000000000000000000000, /* 3559 */
128'h00000000000000000000000000000000, /* 3560 */
128'h00000000000000000000000000000000, /* 3561 */
128'h00000000000000000000000000000000, /* 3562 */
128'h00000000000000000000000000000000, /* 3563 */
128'h00000000000000000000000000000000, /* 3564 */
128'h00000000000000000000000000000000, /* 3565 */
128'h00000000000000000000000000000000, /* 3566 */
128'h00000000000000000000000000000000, /* 3567 */
128'h00000000000000000000000000000000, /* 3568 */
128'h00000000000000000000000000000000, /* 3569 */
128'h00000000000000000000000000000000, /* 3570 */
128'h00000000000000000000000000000000, /* 3571 */
128'h00000000000000000000000000000000, /* 3572 */
128'h00000000000000000000000000000000, /* 3573 */
128'h00000000000000000000000000000000, /* 3574 */
128'h00000000000000000000000000000000, /* 3575 */
128'h00000000000000000000000000000000, /* 3576 */
128'h00000000000000000000000000000000, /* 3577 */
128'h00000000000000000000000000000000, /* 3578 */
128'h00000000000000000000000000000000, /* 3579 */
128'h00000000000000000000000000000000, /* 3580 */
128'h00000000000000000000000000000000, /* 3581 */
128'h00000000000000000000000000000000, /* 3582 */
128'h00000000000000000000000000000000, /* 3583 */
128'h00000000000000000000000000000000, /* 3584 */
128'h00000000000000000000000000000000, /* 3585 */
128'h00000000000000000000000000000000, /* 3586 */
128'h00000000000000000000000000000000, /* 3587 */
128'h00000000000000000000000000000000, /* 3588 */
128'h00000000000000000000000000000000, /* 3589 */
128'h00000000000000000000000000000000, /* 3590 */
128'h00000000000000000000000000000000, /* 3591 */
128'h00000000000000000000000000000000, /* 3592 */
128'h00000000000000000000000000000000, /* 3593 */
128'h00000000000000000000000000000000, /* 3594 */
128'h00000000000000000000000000000000, /* 3595 */
128'h00000000000000000000000000000000, /* 3596 */
128'h00000000000000000000000000000000, /* 3597 */
128'h00000000000000000000000000000000, /* 3598 */
128'h00000000000000000000000000000000, /* 3599 */
128'h00000000000000000000000000000000, /* 3600 */
128'h00000000000000000000000000000000, /* 3601 */
128'h00000000000000000000000000000000, /* 3602 */
128'h00000000000000000000000000000000, /* 3603 */
128'h00000000000000000000000000000000, /* 3604 */
128'h00000000000000000000000000000000, /* 3605 */
128'h00000000000000000000000000000000, /* 3606 */
128'h00000000000000000000000000000000, /* 3607 */
128'h00000000000000000000000000000000, /* 3608 */
128'h00000000000000000000000000000000, /* 3609 */
128'h00000000000000000000000000000000, /* 3610 */
128'h00000000000000000000000000000000, /* 3611 */
128'h00000000000000000000000000000000, /* 3612 */
128'h00000000000000000000000000000000, /* 3613 */
128'h00000000000000000000000000000000, /* 3614 */
128'h00000000000000000000000000000000, /* 3615 */
128'h00000000000000000000000000000000, /* 3616 */
128'h00000000000000000000000000000000, /* 3617 */
128'h00000000000000000000000000000000, /* 3618 */
128'h00000000000000000000000000000000, /* 3619 */
128'h00000000000000000000000000000000, /* 3620 */
128'h00000000000000000000000000000000, /* 3621 */
128'h00000000000000000000000000000000, /* 3622 */
128'h00000000000000000000000000000000, /* 3623 */
128'h00000000000000000000000000000000, /* 3624 */
128'h00000000000000000000000000000000, /* 3625 */
128'h00000000000000000000000000000000, /* 3626 */
128'h00000000000000000000000000000000, /* 3627 */
128'h00000000000000000000000000000000, /* 3628 */
128'h00000000000000000000000000000000, /* 3629 */
128'h00000000000000000000000000000000, /* 3630 */
128'h00000000000000000000000000000000, /* 3631 */
128'h00000000000000000000000000000000, /* 3632 */
128'h00000000000000000000000000000000, /* 3633 */
128'h00000000000000000000000000000000, /* 3634 */
128'h00000000000000000000000000000000, /* 3635 */
128'h00000000000000000000000000000000, /* 3636 */
128'h00000000000000000000000000000000, /* 3637 */
128'h00000000000000000000000000000000, /* 3638 */
128'h00000000000000000000000000000000, /* 3639 */
128'h00000000000000000000000000000000, /* 3640 */
128'h00000000000000000000000000000000, /* 3641 */
128'h00000000000000000000000000000000, /* 3642 */
128'h00000000000000000000000000000000, /* 3643 */
128'h00000000000000000000000000000000, /* 3644 */
128'h00000000000000000000000000000000, /* 3645 */
128'h00000000000000000000000000000000, /* 3646 */
128'h00000000000000000000000000000000, /* 3647 */
128'h00000000000000000000000000000000, /* 3648 */
128'h00000000000000000000000000000000, /* 3649 */
128'h00000000000000000000000000000000, /* 3650 */
128'h00000000000000000000000000000000, /* 3651 */
128'h00000000000000000000000000000000, /* 3652 */
128'h00000000000000000000000000000000, /* 3653 */
128'h00000000000000000000000000000000, /* 3654 */
128'h00000000000000000000000000000000, /* 3655 */
128'h00000000000000000000000000000000, /* 3656 */
128'h00000000000000000000000000000000, /* 3657 */
128'h00000000000000000000000000000000, /* 3658 */
128'h00000000000000000000000000000000, /* 3659 */
128'h00000000000000000000000000000000, /* 3660 */
128'h00000000000000000000000000000000, /* 3661 */
128'h00000000000000000000000000000000, /* 3662 */
128'h00000000000000000000000000000000, /* 3663 */
128'h00000000000000000000000000000000, /* 3664 */
128'h00000000000000000000000000000000, /* 3665 */
128'h00000000000000000000000000000000, /* 3666 */
128'h00000000000000000000000000000000, /* 3667 */
128'h00000000000000000000000000000000, /* 3668 */
128'h00000000000000000000000000000000, /* 3669 */
128'h00000000000000000000000000000000, /* 3670 */
128'h00000000000000000000000000000000, /* 3671 */
128'h00000000000000000000000000000000, /* 3672 */
128'h00000000000000000000000000000000, /* 3673 */
128'h00000000000000000000000000000000, /* 3674 */
128'h00000000000000000000000000000000, /* 3675 */
128'h00000000000000000000000000000000, /* 3676 */
128'h00000000000000000000000000000000, /* 3677 */
128'h00000000000000000000000000000000, /* 3678 */
128'h00000000000000000000000000000000, /* 3679 */
128'h00000000000000000000000000000000, /* 3680 */
128'h00000000000000000000000000000000, /* 3681 */
128'h00000000000000000000000000000000, /* 3682 */
128'h00000000000000000000000000000000, /* 3683 */
128'h00000000000000000000000000000000, /* 3684 */
128'h00000000000000000000000000000000, /* 3685 */
128'h00000000000000000000000000000000, /* 3686 */
128'h00000000000000000000000000000000, /* 3687 */
128'h00000000000000000000000000000000, /* 3688 */
128'h00000000000000000000000000000000, /* 3689 */
128'h00000000000000000000000000000000, /* 3690 */
128'h00000000000000000000000000000000, /* 3691 */
128'h00000000000000000000000000000000, /* 3692 */
128'h00000000000000000000000000000000, /* 3693 */
128'h00000000000000000000000000000000, /* 3694 */
128'h00000000000000000000000000000000, /* 3695 */
128'h00000000000000000000000000000000, /* 3696 */
128'h00000000000000000000000000000000, /* 3697 */
128'h00000000000000000000000000000000, /* 3698 */
128'h00000000000000000000000000000000, /* 3699 */
128'h00000000000000000000000000000000, /* 3700 */
128'h00000000000000000000000000000000, /* 3701 */
128'h00000000000000000000000000000000, /* 3702 */
128'h00000000000000000000000000000000, /* 3703 */
128'h00000000000000000000000000000000, /* 3704 */
128'h00000000000000000000000000000000, /* 3705 */
128'h00000000000000000000000000000000, /* 3706 */
128'h00000000000000000000000000000000, /* 3707 */
128'h00000000000000000000000000000000, /* 3708 */
128'h00000000000000000000000000000000, /* 3709 */
128'h00000000000000000000000000000000, /* 3710 */
128'h00000000000000000000000000000000, /* 3711 */
128'h00000000000000000000000000000000, /* 3712 */
128'h00000000000000000000000000000000, /* 3713 */
128'h00000000000000000000000000000000, /* 3714 */
128'h00000000000000000000000000000000, /* 3715 */
128'h00000000000000000000000000000000, /* 3716 */
128'h00000000000000000000000000000000, /* 3717 */
128'h00000000000000000000000000000000, /* 3718 */
128'h00000000000000000000000000000000, /* 3719 */
128'h00000000000000000000000000000000, /* 3720 */
128'h00000000000000000000000000000000, /* 3721 */
128'h00000000000000000000000000000000, /* 3722 */
128'h00000000000000000000000000000000, /* 3723 */
128'h00000000000000000000000000000000, /* 3724 */
128'h00000000000000000000000000000000, /* 3725 */
128'h00000000000000000000000000000000, /* 3726 */
128'h00000000000000000000000000000000, /* 3727 */
128'h00000000000000000000000000000000, /* 3728 */
128'h00000000000000000000000000000000, /* 3729 */
128'h00000000000000000000000000000000, /* 3730 */
128'h00000000000000000000000000000000, /* 3731 */
128'h00000000000000000000000000000000, /* 3732 */
128'h00000000000000000000000000000000, /* 3733 */
128'h00000000000000000000000000000000, /* 3734 */
128'h00000000000000000000000000000000, /* 3735 */
128'h00000000000000000000000000000000, /* 3736 */
128'h00000000000000000000000000000000, /* 3737 */
128'h00000000000000000000000000000000, /* 3738 */
128'h00000000000000000000000000000000, /* 3739 */
128'h00000000000000000000000000000000, /* 3740 */
128'h00000000000000000000000000000000, /* 3741 */
128'h00000000000000000000000000000000, /* 3742 */
128'h00000000000000000000000000000000, /* 3743 */
128'h00000000000000000000000000000000, /* 3744 */
128'h00000000000000000000000000000000, /* 3745 */
128'h00000000000000000000000000000000, /* 3746 */
128'h00000000000000000000000000000000, /* 3747 */
128'h00000000000000000000000000000000, /* 3748 */
128'h00000000000000000000000000000000, /* 3749 */
128'h00000000000000000000000000000000, /* 3750 */
128'h00000000000000000000000000000000, /* 3751 */
128'h00000000000000000000000000000000, /* 3752 */
128'h00000000000000000000000000000000, /* 3753 */
128'h00000000000000000000000000000000, /* 3754 */
128'h00000000000000000000000000000000, /* 3755 */
128'h00000000000000000000000000000000, /* 3756 */
128'h00000000000000000000000000000000, /* 3757 */
128'h00000000000000000000000000000000, /* 3758 */
128'h00000000000000000000000000000000, /* 3759 */
128'h00000000000000000000000000000000, /* 3760 */
128'h00000000000000000000000000000000, /* 3761 */
128'h00000000000000000000000000000000, /* 3762 */
128'h00000000000000000000000000000000, /* 3763 */
128'h00000000000000000000000000000000, /* 3764 */
128'h00000000000000000000000000000000, /* 3765 */
128'h00000000000000000000000000000000, /* 3766 */
128'h00000000000000000000000000000000, /* 3767 */
128'h00000000000000000000000000000000, /* 3768 */
128'h00000000000000000000000000000000, /* 3769 */
128'h00000000000000000000000000000000, /* 3770 */
128'h00000000000000000000000000000000, /* 3771 */
128'h00000000000000000000000000000000, /* 3772 */
128'h00000000000000000000000000000000, /* 3773 */
128'h00000000000000000000000000000000, /* 3774 */
128'h00000000000000000000000000000000, /* 3775 */
128'h00000000000000000000000000000000, /* 3776 */
128'h00000000000000000000000000000000, /* 3777 */
128'h00000000000000000000000000000000, /* 3778 */
128'h00000000000000000000000000000000, /* 3779 */
128'h00000000000000000000000000000000, /* 3780 */
128'h00000000000000000000000000000000, /* 3781 */
128'h00000000000000000000000000000000, /* 3782 */
128'h00000000000000000000000000000000, /* 3783 */
128'h00000000000000000000000000000000, /* 3784 */
128'h00000000000000000000000000000000, /* 3785 */
128'h00000000000000000000000000000000, /* 3786 */
128'h00000000000000000000000000000000, /* 3787 */
128'h00000000000000000000000000000000, /* 3788 */
128'h00000000000000000000000000000000, /* 3789 */
128'h00000000000000000000000000000000, /* 3790 */
128'h00000000000000000000000000000000, /* 3791 */
128'h00000000000000000000000000000000, /* 3792 */
128'h00000000000000000000000000000000, /* 3793 */
128'h00000000000000000000000000000000, /* 3794 */
128'h00000000000000000000000000000000, /* 3795 */
128'h00000000000000000000000000000000, /* 3796 */
128'h00000000000000000000000000000000, /* 3797 */
128'h00000000000000000000000000000000, /* 3798 */
128'h00000000000000000000000000000000, /* 3799 */
128'h00000000000000000000000000000000, /* 3800 */
128'h00000000000000000000000000000000, /* 3801 */
128'h00000000000000000000000000000000, /* 3802 */
128'h00000000000000000000000000000000, /* 3803 */
128'h00000000000000000000000000000000, /* 3804 */
128'h00000000000000000000000000000000, /* 3805 */
128'h00000000000000000000000000000000, /* 3806 */
128'h00000000000000000000000000000000, /* 3807 */
128'h00000000000000000000000000000000, /* 3808 */
128'h00000000000000000000000000000000, /* 3809 */
128'h00000000000000000000000000000000, /* 3810 */
128'h00000000000000000000000000000000, /* 3811 */
128'h00000000000000000000000000000000, /* 3812 */
128'h00000000000000000000000000000000, /* 3813 */
128'h00000000000000000000000000000000, /* 3814 */
128'h00000000000000000000000000000000, /* 3815 */
128'h00000000000000000000000000000000, /* 3816 */
128'h00000000000000000000000000000000, /* 3817 */
128'h00000000000000000000000000000000, /* 3818 */
128'h00000000000000000000000000000000, /* 3819 */
128'h00000000000000000000000000000000, /* 3820 */
128'h00000000000000000000000000000000, /* 3821 */
128'h00000000000000000000000000000000, /* 3822 */
128'h00000000000000000000000000000000, /* 3823 */
128'h00000000000000000000000000000000, /* 3824 */
128'h00000000000000000000000000000000, /* 3825 */
128'h00000000000000000000000000000000, /* 3826 */
128'h00000000000000000000000000000000, /* 3827 */
128'h00000000000000000000000000000000, /* 3828 */
128'h00000000000000000000000000000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00000000000000000000000000000000, /* 3840 */
128'h00000000000000000000000000000000, /* 3841 */
128'h00000000000000000000000000000000, /* 3842 */
128'h00000000000000000000000000000000, /* 3843 */
128'h00000000000000000000000000000000, /* 3844 */
128'h00000000000000000000000000000000, /* 3845 */
128'h00000000000000000000000000000000, /* 3846 */
128'h00000000000000000000000000000000, /* 3847 */
128'h00000000000000000000000000000000, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule

