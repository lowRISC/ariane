/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'h011111133ff1011b0000413711249463, /*    1 */
128'h00008297000280e70482829300008297, /*    2 */
128'h000280e7130505130000051706e28293, /*    3 */
128'ha1c606130000c617fc05859300000597, /*    4 */
128'h000f4eb7011696933ff6869b000046b7, /*    5 */
128'h0085b703fffe8e930005b703240e8e9b, /*    6 */
128'hff81011301b111130110011bfe0e9ae3, /*    7 */
128'h0085b70300e6b0230005b7030006b703, /*    8 */
128'h0185b70300e6b8230105b70300e6b423, /*    9 */
128'hfcc5cce3020686930205859300e6bc23, /*   10 */
128'h40b787b300d787b30147879300000797, /*   11 */
128'h30579073090787930000079700078067, /*   12 */
128'h1c8606130000c617a30585930000c597, /*   13 */
128'h0005bc230005b8230005b4230005b023, /*   14 */
128'h020004b7650090effec5c6e302058593, /*   15 */
128'h02000937004484930124a02300100913, /*   16 */
128'h3440297310500073ff24c6e34009091b, /*   17 */
128'hf1402973020004b7fe090ae300897913, /*   18 */
128'h0004a903000920230099093300291913, /*   19 */
128'h4009091b0200093700448493fe091ee3, /*   20 */
128'h1050007334102373342022f3ff24c6e3, /*   21 */
128'h41206d6f7266206f6c6c6548ffdff06f, /*   22 */
128'h617720657361656c502021656e616972, /*   23 */
128'h000a2e2e2e746e656d6f6d2061207469, /*   24 */
128'h00000000000000000000000000000000, /*   25 */
128'h00000000000000000000000000000000, /*   26 */
128'h00000000000000000000000000000000, /*   27 */
128'h00000000000000000000000000000000, /*   28 */
128'h00000000000000000000000000000000, /*   29 */
128'h00000000000000000000000000000000, /*   30 */
128'h00000000000000000000000000000000, /*   31 */
128'hd963454c0005cc635735c28587ae6914, /*   32 */
128'he21c97b6470102a787b30a00051300b7, /*   33 */
128'h853e85b200030563018533038082853a, /*   34 */
128'h6f8686930000b697b7edfda007138302, /*   35 */
128'h87930000c7976294824707130000c717, /*   36 */
128'h87b30280069302d787bb878d8f9981a7, /*   37 */
128'h47148082853a470100e7956397ba02d7, /*   38 */
128'hf0efe4061141b7f502870713fea68de3, /*   39 */
128'hbfe545018082014160a26108c509fbbf, /*   40 */
128'hf0efe852ec4ef04af426f822fc067139, /*   41 */
128'h0000ba17440144814985892acd31f9bf, /*   42 */
128'hc091553500f44d6300c9278327ca0a13, /*   43 */
128'h61216a4269e2790274a2744270e24501, /*   44 */
128'h67a2ed19f29ff0ef854a85a200308082, /*   45 */
128'h50ef8552000995632485cb990087c783, /*   46 */
128'h0513bf6524051de080ef4981652245c0, /*   47 */
128'hf2dff0efe42ef406f0227179b7c1fda0, /*   48 */
128'h842aee7ff0ef083065a2c105fda00413, /*   49 */
128'h00f7096300c547030ff007936562e911, /*   50 */
128'h547980826145740270a285221a4080ef, /*   51 */
128'hf0efec4ef04af426f822fc067139bfd5, /*   52 */
128'h0000a9970ff00913440184aacd01eebf, /*   53 */
128'h74a2744270e200f4496344dc39498993, /*   54 */
128'hf0ef852685a200308082612169e27902, /*   55 */
128'h85a20127896300c7c78367a2ed09e83f, /*   56 */
128'hb7d9240513e080ef65223b8050ef854e, /*   57 */
128'he8dff0ef892eec26f406e84af0227179, /*   58 */
128'he45ff0ef84aa85ca0030c11dfda00413, /*   59 */
128'h338505130000a517864a608ced01842a, /*   60 */
128'h740270a28522100080ef652237a050ef, /*   61 */
128'hf406ec26f022717980826145694264e2, /*   62 */
128'h85a6842ac11dfda00413e47ff0ef84ae, /*   63 */
128'hcf63445c342050ef310505130000a517, /*   64 */
128'h54350c6080ef30e505130000a51700f4, /*   65 */
128'h003085228082614564e2740270a28522, /*   66 */
128'h09a080ef6522f565842adcfff0ef85a6, /*   67 */
128'h5479fcf71be30ff0079300c7c70367a2, /*   68 */
128'he50965a2de1ff0eff406e42e7179bfc1, /*   69 */
128'hf96dd97ff0ef08308082614570a24501, /*   70 */
128'he42eec064108842ae8221101bfc56562, /*   71 */
128'h852200030e6302053303c919db9ff0ef, /*   72 */
128'h60e2fda005138302610560e265a26442, /*   73 */
128'h0000b7977139bfdd4501808261056442, /*   74 */
128'h04130000b417f426f822639c48478793, /*   75 */
128'h043b840d8c055a2484930000b4975aa4, /*   76 */
128'h892afc06e852ec4ef04a0280079302f4, /*   77 */
128'h942602f4043324ea0a130000aa1789ae, /*   78 */
128'h69e2790274a2744270e2450100849b63, /*   79 */
128'h23e050ef855285ca6090808261216a42, /*   80 */
128'hbfc902848493c50164b060ef854a608c, /*   81 */
128'hb7e16522f569cdbff0ef852685ce0030, /*   82 */
128'h84b68432e42efc06f04af426f8227139, /*   83 */
128'hcb5ff0ef083065a2c115cf7ff0ef893a, /*   84 */
128'h70e2978285a2615c862686ca6562e519, /*   85 */
128'hbfc5fda0051380826121790274a27442, /*   86 */
128'h84b68432e42efc06f04af426f8227139, /*   87 */
128'hc75ff0ef083065a2c115cb7ff0ef893a, /*   88 */
128'h70e2978285a2655c862686ca6562e519, /*   89 */
128'hbfc5fda0051380826121790274a27442, /*   90 */
128'hc7dff0ef84b2e42ef822fc06f4267139, /*   91 */
128'h701ce509c39ff0ef842a083065a2c105, /*   92 */
128'h8082612174a2744270e2978285a66562, /*   93 */
128'h2785c3190017f713419cbfcdfda00513, /*   94 */
128'hd71b8e5927a106220086571b419cc19c, /*   95 */
128'h0ff77713c19c0087d7138ed906a20086, /*   96 */
128'h122300d5112300c510238fd90087979b, /*   97 */
128'hf022f4067179419c80820005132300f5, /*   98 */
128'h419c00f510230457879b6785c19c27d1, /*   99 */
128'h0087979b0ff777130087d713c632842a, /*  100 */
128'hc4360509084c57fd460900f11a238fd9, /*  101 */
128'h0513016105934609739060ef00f11b23, /*  102 */
128'h00041323082c462147c172b060ef0044, /*  103 */
128'h00f404a347c5717060efec3e00840513, /*  104 */
128'h701060ef00c4051300041523006c4611, /*  105 */
128'h014406936f5060ef01040513002c4611, /*  106 */
128'hfed79ce39f31ffe7d6030789470187a2, /*  107 */
128'h9fb94107d71b9fb9934117424107579b, /*  108 */
128'h80826145740270a200f41523fff7c793, /*  109 */
128'h97ba46a167856398338787930000b797, /*  110 */
128'hc7bb27850077e793fff6079b8007bc23, /*  111 */
128'h3823973e678500f547636805450102d7, /*  112 */
128'h010686bb0035169b0005b883808280c7, /*  113 */
128'he0221141bff105a125050116b02396ba, /*  114 */
128'hfa5ff0efe406450185aa86220005841b, /*  115 */
128'hec26f022717980820141640260a28522, /*  116 */
128'h641060efe436f4064619051984b2842a, /*  117 */
128'h162347a1635060ef85b64619852266a2, /*  118 */
128'h614564e200e4859b70a27402852200f4, /*  119 */
128'h3a8130236785737dc5010113fadff06f, /*  120 */
128'h3931342338913c233a11342339213823, /*  121 */
128'h377134233761382337513c2339413023, /*  122 */
128'h3507879335a1382335913c2337813023, /*  123 */
128'hce042023d00007b7943e747d978a911a, /*  124 */
128'hd0040023f0040023e0040023ca040b23, /*  125 */
128'ha51785aa00e7ea63892a5800073797aa, /*  126 */
128'h00054703a001755040eff52505130000, /*  127 */
128'h970a3507871374fd678526f711634789, /*  128 */
128'hcb848b13970a350787139abacd848a93, /*  129 */
128'h9c3a9b3a49818a368cb28baed0048c13, /*  130 */
128'hc7830015cd03013907b395ca0f098593, /*  131 */
128'h869b01a989bb058902a0071329890f07, /*  132 */
128'h24e78163471904f76b6326e78d630007, /*  133 */
128'hcc848513470d2ae78963470502f76263, /*  134 */
128'h40ef052505130000a51785b622e78963, /*  135 */
128'hfee794e3473d22e785634731b77d6cd0, /*  136 */
128'h953e866ae0048513978a350787936785, /*  137 */
128'h03600713b759e00d00234fb060ef9d22, /*  138 */
128'h22e780630330071300f76e6322e78363, /*  139 */
128'haad94605cb648513fae798e303500713, /*  140 */
128'hf8e79ce30ff0071324e7856303800713, /*  141 */
128'h24e781630007859b747d471500614783, /*  142 */
128'h000ca7833ae79d63470938e781634719, /*  143 */
128'h05134985978a350a87936a8516079263, /*  144 */
128'h60ef013ca023953e461101090593ce44, /*  145 */
128'h01490593ce840513978a350a879347f0, /*  146 */
128'he28505130000a517469060ef953e4611, /*  147 */
128'h978a350a8793605040efde0254e25a52, /*  148 */
128'h3ef060ef854a55fd4619993ecf840913, /*  149 */
128'h879346f115231350079300f103a3478d, /*  150 */
128'h85a6460594becb740493c2a6978a350a, /*  151 */
128'h06a303200793417060efc0d246c10513, /*  152 */
128'h4a1195becf040593978a350a879346f1, /*  153 */
128'h07933f3060ef4741072346f105134611, /*  154 */
128'hcf440593978a350a879346f109a30360, /*  155 */
128'h3d1060ef47410a2347510513461195be, /*  156 */
128'h03a346f10ca347b1051385a6460557fd, /*  157 */
128'h0613102007933b7060ef47310d230001, /*  158 */
128'h0793351060efde3e37a1051345810f00, /*  159 */
128'h3961051385de4799464136f11d231010, /*  160 */
128'h13232637879377e1389060ef36f10e23, /*  161 */
128'h350a879346f1142335378793679946f1, /*  162 */
128'h0440061304300693943ecec40413978a, /*  163 */
128'h85a2460156fdba1ff0ef3721051385a2, /*  164 */
128'h0e8885de86ca5672bd5ff0ef35e10513, /*  165 */
128'h3a0134033a813083911a6305cebff0ef, /*  166 */
128'h38013a03388139833901390339813483, /*  167 */
128'h36013c0336813b8337013b0337813a83, /*  168 */
128'h851380823b01011335013d0335813c83, /*  169 */
128'ha00d953e978a3507879367854611cd04, /*  170 */
128'h953e866af0048513978a350787936785, /*  171 */
128'h85564611b39df00d00232db060ef9d22, /*  172 */
128'h87936785bfdd855a4611bbb12cd060ef, /*  173 */
128'h2b1060ef4611953ece048513978a3507, /*  174 */
128'h00f40123ce14478300f401a3ce044783, /*  175 */
128'h00f40023ce34478300f400a3ce244783, /*  176 */
128'h866ab759cc048513bb29cef42023401c, /*  177 */
128'h2783b311d00d0023279060ef9d228562, /*  178 */
128'h0000a51700fa2023478512079a63000a, /*  179 */
128'h0e88010905934611407040efc3c50513, /*  180 */
128'hcb840513978a35048793648524d060ef, /*  181 */
128'h35314703235060ef014905934611953e, /*  182 */
128'h0000a517350145833511460335214683, /*  183 */
128'h00a14683350157833c7040efc0c50513, /*  184 */
128'h35215783fcf71e230000b71700914603, /*  185 */
128'h0000b717c0c505130000a51700814583, /*  186 */
128'h01b14703393040ef00b14703fcf71323, /*  187 */
128'h0000a517018145830191460301a14683, /*  188 */
128'h0121468301314703377040efc0c50513, /*  189 */
128'hc10505130000a5170101458301114603, /*  190 */
128'h05130000a51755c20101578335b040ef, /*  191 */
128'hb71701215783f6f713230000b717c1e5, /*  192 */
128'hf6bb02f5d63b03c00793f4f71e230000, /*  193 */
128'h02f5d5bbe107879b678502f6763b02f5, /*  194 */
128'h95bee0040593978a3504879331b040ef, /*  195 */
128'h35048793303040efbf8505130000a517, /*  196 */
128'hbf0505130000a51795be978af0040593, /*  197 */
128'h40efbfa505130000a517b5012eb040ef, /*  198 */
128'h20234785de0796e3000a2783bbcd2dd0, /*  199 */
128'ha5172c1040efbee505130000a51700fa, /*  200 */
128'h3507879367852b5040efbf2505130000, /*  201 */
128'hbf8505130000a51795be978ad0040593, /*  202 */
128'hb35d291040efbfe505130000a517bf45, /*  203 */
128'hf852fc4ee0cae4a6e8a2ec86711d737d, /*  204 */
128'h6a85c12505130000a517911a89aaf456, /*  205 */
128'h0493978a020a8793747d269040efca02, /*  206 */
128'hb797051060ef852655fd461994beff84, /*  207 */
128'hc83e4a05fef40913439cd02787930000, /*  208 */
128'h993e978a020a879312f11d2313500793, /*  209 */
128'h0793073060ef014107a31a68460585ca, /*  210 */
128'h020a879312f10f23479112f10ea30370, /*  211 */
128'h60ef13f10513461195beff040593978a, /*  212 */
128'h14f101a314510513460585ca57fd04f0, /*  213 */
128'h0fc00793035060ef000107a315410223, /*  214 */
128'h7ce060efca3e04a1051345810f000613, /*  215 */
128'h05134641479985ce04f1152310100793, /*  216 */
128'h2637879377e1007060ef04f106230661, /*  217 */
128'h879312f11c2335378793679912f11b23, /*  218 */
128'h06930421051385a2943e1451978a020a, /*  219 */
128'h02e1051385a2821ff0ef044006130430, /*  220 */
128'h85ce86a610084652855ff0ef460156fd, /*  221 */
128'h64a66446450160e6911a630596bff0ef, /*  222 */
128'ha51785aa808261257aa27a4279e26906, /*  223 */
128'h3423810101131450406fb02505130000, /*  224 */
128'h34237d2138237c913c237e8130237e11, /*  225 */
128'h893689b2e04605a1051384aa71597d31, /*  226 */
128'h10186785764060efd602e83eec3ae442, /*  227 */
128'h943e7fc404136762747d97ba81078793, /*  228 */
128'hf8aff0efd64e0521051385a2864a86ba, /*  229 */
128'hf0ef03e10513863e86c285a267c26822, /*  230 */
128'h8cfff0ef86c685a6180856326882fbaf, /*  231 */
128'h7d8134837e01340345017e8130836165, /*  232 */
128'h716d80827f0101137c8139837d013903, /*  233 */
128'h003547830045480300554883e222e606, /*  234 */
128'ha597842a000546030015468300254703, /*  235 */
128'h40efa52505130000a517a52585930000, /*  236 */
128'ha597860ac10d842adedff0ef852207d0, /*  237 */
128'h40efa5a505130000a517a32585930000, /*  238 */
128'h0000a51780826151641260b2852205d0, /*  239 */
128'h03f040efbe07ae230000b797a7450513, /*  240 */
128'hf85afc56e0d2e4ceeca6f0a27159b7cd, /*  241 */
128'h8a2ae46ee8caf486e86aec66f062f45e, /*  242 */
128'h718a8a930000aa974401ff05049389ae, /*  243 */
128'h0000ac1706000b93a48b0b130000ab17, /*  244 */
128'hfff58d1ba44c8c930000ac97a54c0c13, /*  245 */
128'h6a0669a6694664e6740670a603344163, /*  246 */
128'h61656da26d426ce27c027ba27b427ae2, /*  247 */
128'h7be040ef855ae7a9c42900f477938082, /*  248 */
128'hfe05879b0007c583012487b34dc14901, /*  249 */
128'h09057a0040ef856602fbe2630ff7f793, /*  250 */
128'h78e040ef574505130000a517ffb912e3, /*  251 */
128'hb7c5780040ef8562a031788040ef8556, /*  252 */
128'h40ef9d2505130000a5170104c583dbe5, /*  253 */
128'h00f979134d81fffd4913028d1d6376c0, /*  254 */
128'h855aff2dcce32d85756040ef8556a029, /*  255 */
128'h00f45b630009079bff04791374a040ef, /*  256 */
128'h04852405732040ef518505130000a517, /*  257 */
128'hf793fe05879b0007c583012a07b3b781, /*  258 */
128'hb7e90905712040ef856600fbe7630ff7, /*  259 */
128'he44ee84aec267179bfdd708040ef8562, /*  260 */
128'h86930000a697893289ae84b6f022f406, /*  261 */
128'h0000971794c686930000a697c50919e6, /*  262 */
128'h854a85a6944606130000a617dfc70713, /*  263 */
128'h85bb00955d6300098f63842a68a040ef, /*  264 */
128'h40ef954a92c606130000a61786ce40a4, /*  265 */
128'hffd4841b00f44463ffe4879b9c2966c0, /*  266 */
128'h224060ef8fc585930000a59700890533, /*  267 */
128'h8082614569a2694264e2854a740270a2, /*  268 */
128'h0613002c7115f73ff06f4581862e86b2, /*  269 */
128'h0000a517002cfebff0efed8645050c80, /*  270 */
128'h8082612d450160ee656040ef8e450513, /*  271 */
128'h47b704a76963862e9ff787133b9ad7b7, /*  272 */
128'hf7633e70079304a7676323f78713000f, /*  273 */
128'h8e8707130000b7173e80079346890ca7, /*  274 */
128'he426e822ec0600074903e04a97361101, /*  275 */
128'ha51785aa690264a260e2644202091663, /*  276 */
128'h879346815f20406f610588a505130000, /*  277 */
128'h02f57433bf7d240787934685b7d9a007, /*  278 */
128'h0287e66347293e800793c02102f555b3, /*  279 */
128'h0287746306300713c70502f4773347a9, /*  280 */
128'h0324341302e4743302f457b306400713, /*  281 */
128'h5433bfc102e45433a039943e00144413, /*  282 */
128'h40ef84b2834505130000a517f86102f4, /*  283 */
128'h40ef82a505130000a51785a2c80158c0, /*  284 */
128'ha517690264a285ca862660e2644257c0, /*  285 */
128'h951785aa5620406f610581a505130000, /*  286 */
128'h481958d94781862eb78d7ea505130000, /*  287 */
128'h1782cd8500e555b303c6871b02f886bb, /*  288 */
128'he42697c211017f6808130000a8179381, /*  289 */
128'h60e26442e495e04ae822ec060007c483, /*  290 */
128'h61057ca505130000951785aa690264a2, /*  291 */
128'h0000951785aafb079de3278550a0406f, /*  292 */
128'hfff7c79300e797b357fdb7f57b450513, /*  293 */
128'h03b6869b02f5053347a9c10d44018d7d, /*  294 */
128'hf46300e45433942a47a500d414334405, /*  295 */
128'h89327625051300009517058514590087, /*  296 */
128'h758505130000951785a2c8014ba040ef, /*  297 */
128'h64a2690285a6864a60e264424aa040ef, /*  298 */
128'h71514900406f61057605051300009517, /*  299 */
128'he96ae5cee9caf1a202c7073b8cbaed66, /*  300 */
128'he56ef162f55ef95afd56e1d2eda6f586, /*  301 */
128'h00e7f66384368d3289ae892a04000793, /*  302 */
128'hdcbb4cc1000c956302ccdcbb04000c93, /*  303 */
128'h0017849be03e020d1a13001d179b03ac, /*  304 */
128'h708b0b1300009b1703810a93020a5a13, /*  305 */
128'h5d8c0c1300008c17670b8b9300009b97, /*  306 */
128'h6a0e69ae694e64ee740e70ae4501e00d, /*  307 */
128'h616d6daa6d4a6cea7c0a7baa7b4a7aea, /*  308 */
128'h3ee040ef6c4505130000951785ca8082, /*  309 */
128'h470186ce000c8d9b008cf46300040d9b, /*  310 */
128'h971305b66c630007061b430948a14811, /*  311 */
128'h06bb0d9de66399ba034707339301020d, /*  312 */
128'h415705bb0006861b02e00813875603bd, /*  313 */
128'h05130000951785d6963e011c0ac5ed63, /*  314 */
128'h043b66a2392040effa060c23e43667e5, /*  315 */
128'h557dd13506e070ef99369281168241b4, /*  316 */
128'h260195d6002715934290030d1b63b795, /*  317 */
128'hec42f046f41a855a658292011602c190, /*  318 */
128'h96d27322674266a2356040efe436e83a, /*  319 */
128'h15936290011d1863bf85686278820705, /*  320 */
128'h0006d603006d1c63bfc1e19095d60037, /*  321 */
128'hbf6500c590239241164295d600171593, /*  322 */
128'h00c580230ff6761300ea85b30006c603, /*  323 */
128'h6ae32705672209a070efe43a855eb75d, /*  324 */
128'h053300074583bfdd4701bf1d3cfdfe97, /*  325 */
128'h0185959bc519097575130005450300bc, /*  326 */
128'hbf390705010700230005d4634185d59b, /*  327 */
128'h8082e21c00b7f4634501918187aa1582, /*  328 */
128'h89aa04000613fd4e7115bfd58f8d2505, /*  329 */
128'hf556f952e1cae5a6e9a2ed8600884581, /*  330 */
128'h577d67869982e16ae566e962ed5ef15a, /*  331 */
128'h55796318474707130000a7178ff98361, /*  332 */
128'h00009b174a8503800a13440106e79d63, /*  333 */
128'h80000c3758cb8b9300009b97554b0b13, /*  334 */
128'h07815783564d0d1300009d1708000cb7, /*  335 */
128'h06137786028a05bba091656600f46463, /*  336 */
128'h77c20957926347a299829dbd00280380, /*  337 */
128'h040908637922224040ef855a85a2cfbd, /*  338 */
128'h0000951785a60397e863018487b37482, /*  339 */
128'h64ae644e60ee5575206040ef50450513, /*  340 */
128'h6caa6c4a6bea7b0a7aaa7a4a79ea690e, /*  341 */
128'h40ef856a86ca85a666428082612d6d0a, /*  342 */
128'h77a274c2998285260009061b45c21dc0, /*  343 */
128'h855e85ca993e86268c9d79020097ff63, /*  344 */
128'h24057b1050ef854a458186261ba040ef, /*  345 */
128'ha7178082400005378082057e4505bfb1, /*  346 */
128'h869300756513157d631c57a707130000, /*  347 */
128'h057e450597aa20000537e30895360017, /*  348 */
128'h862a0ce507638207871367858082953e, /*  349 */
128'h4b050513000095178087871308a74463, /*  350 */
128'h000095178006079b04c7496306e60b63, /*  351 */
128'h0000951787f787936785c3ad48c50513, /*  352 */
128'h11417c07879b77fd04c7c96350c50513, /*  353 */
128'h05130000a5174fe58593000095979e3d, /*  354 */
128'h05130000a51760a20f2040efe4064de5, /*  355 */
128'h05130000951781078713808201414ce5, /*  356 */
128'h0513000095178187879300e60a6345e5, /*  357 */
128'h00009517830787138082faf612e345e5, /*  358 */
128'h8287879300c74963fee609e347c50513, /*  359 */
128'h951783878713bfe94585051300009517, /*  360 */
128'h951784078793fce608e346a505130000, /*  361 */
128'h4205051300009517bf7546a505130000, /*  362 */
128'h84ae892af406e84aec26f02271798082, /*  363 */
128'h942a9041144201045513029044634401, /*  364 */
128'h1542fff54513740270a2952201045513, /*  365 */
128'h0068460985ca808261459141694264e2, /*  366 */
128'h00f107a334f9090900c147836ad050ef, /*  367 */
128'hbf55943e00e1578300f1072300d14783, /*  368 */
128'h8793f44ef84afc26e486e0a26785715d, /*  369 */
128'h0e636dd7879367a13cf50563842e8067, /*  370 */
128'h082884b205e944079a638005079b0af5, /*  371 */
128'ha517461985ca0064091365b050ef4611, /*  372 */
128'h079301744583647050ef3d2505130000, /*  373 */
128'h1cf5826347b108b7e76332f5896302e0, /*  374 */
128'h478502b7e3631af58363479104b7e563, /*  375 */
128'h83633aa5051300009517478910f58463, /*  376 */
128'ha41d7b1030ef546505130000951702f5, /*  377 */
128'h3b0505130000951747a118f582634799, /*  378 */
128'h2cf5826347f5a431797030effef591e3, /*  379 */
128'h0000951747d916f58a6347c500b7ed63, /*  380 */
128'h866302100793bf6dfef580e33cc50513, /*  381 */
128'h051300009517faf596e3029007932af5, /*  382 */
128'h04b7e2632cf5826306200793b7c93e65, /*  383 */
128'h02f0079300b7ef632af5826303300793, /*  384 */
128'h3e850513000095170320079328f58763, /*  385 */
128'h079328f5846305c00793b7bdf8f58ae3, /*  386 */
128'hbf91f6f58de33fe505130000951705e0, /*  387 */
128'h0670079300b7ef6328f5866308400793, /*  388 */
128'h410505130000951706c0079326f58b63, /*  389 */
128'h079326f5886308900793b73df4f58ae3, /*  390 */
128'h9517f0f59ce30880079326f589630ff0, /*  391 */
128'h0000a79701e45703b73d41a505130000, /*  392 */
128'h12f714632dc989930000a9972e47d783, /*  393 */
128'h10f71c632ce7d7830000a79702045703, /*  394 */
128'h0000a59746194e7050ef852285ca4619, /*  395 */
128'h012301a457834d7050ef854a29c58593, /*  396 */
128'h859b01c4578300f41f23020412230204, /*  397 */
128'h1d230009d78302f4102302240513fde4, /*  398 */
128'h0ea3db9ff0ef00f41e230029d78300f4, /*  399 */
128'h1223862601c1578300a10e23812100a1, /*  400 */
128'h00009517a06ddcbfe0ef450185a202f4, /*  401 */
128'hb55922a5051300009517bd4121c50513, /*  402 */
128'h470302444783bdb52385051300009517, /*  403 */
128'h178300f10e230254478300f10ea30264, /*  404 */
128'h00e10e2327810274470300e10ea301c1, /*  405 */
128'h0234470300e10ea301c1190302244703, /*  406 */
128'h04e79b6301c156830450071300e10e23, /*  407 */
128'h0000a597461947e21ad79e230000a797, /*  408 */
128'h0000a71719c505130000a51719458593, /*  409 */
128'ha79766a247623f7050efe43618f72e23, /*  410 */
128'h450102a40593ff89061b172787930000, /*  411 */
128'h616179a2794274e2640660a6508060ef, /*  412 */
128'h0000a71747e204e69463043007138082, /*  413 */
128'hc799439c160787930000a79714f72e23, /*  414 */
128'h0000a697f7e9439c150787930000a797, /*  415 */
128'h0000a597140606130000a61714468693, /*  416 */
128'h0713b765d6dfe0ef02a4051314458593, /*  417 */
128'h30ef152505130000951702e798634d20, /*  418 */
128'h051300009517cdcff0ef852285a651d0, /*  419 */
128'hcc6ff0ef02a4051385ca509030ef14e5, /*  420 */
128'h67c101e45703f6e787e35fe00713bf95, /*  421 */
128'h4611f4f70de302045703f6f701e317fd, /*  422 */
128'hb799323050ef0868100585930000a597, /*  423 */
128'h051300009517b3351285051300009517, /*  424 */
128'h9517bb211445051300009517b30d12e5, /*  425 */
128'h1685051300009517b339152505130000, /*  426 */
128'h00009517b9ed16e5051300009517b311, /*  427 */
128'hb1dd19a5051300009517b9c518c50513, /*  428 */
128'h051300009517b9f11b05051300009517, /*  429 */
128'hd703b1e11e45051300009517b9c91d65, /*  430 */
128'h84930000a49707e7d7830000a7970265, /*  431 */
128'hd7830000a7970285d703ecf711e30764, /*  432 */
128'h89930205891320000793eaf719e30687, /*  433 */
128'h271050ef854a85ce461900f59a230165, /*  434 */
128'h261050ef854e026585930000a5974619, /*  435 */
128'h50ef00640513016585930000a5974619, /*  436 */
128'h01c45783245050ef852285ca461924f0, /*  437 */
128'h02f4142301e4578302f4132302a00613, /*  438 */
128'h00f41f230024d78300f41e230004d783, /*  439 */
128'h0000951785aab36900f4162360800793, /*  440 */
128'h300017b7bba546013b7030ef16c50513, /*  441 */
128'h74132601608130239f0101138307b603, /*  442 */
128'h8406871b0387759366850034171b00f6, /*  443 */
128'h3c23630c8387b783972a300005379f2d, /*  444 */
128'h5f200813ffc5849b2581601134235e91, /*  445 */
128'h00c5963b101005938a1d08b8696335b9, /*  446 */
128'h87930000a797cfb527818ff1fff7c793, /*  447 */
128'h869b7007f7930084179bea254390f4e7, /*  448 */
128'h00d100a3872646d496aa068e9ebd8006, /*  449 */
128'h00d100230086d69b0106d69b0106969b, /*  450 */
128'h806686936685c6918005069b00015503, /*  451 */
128'h67139fad377d8005859b658502d51a63, /*  452 */
128'h868a83f502d7473b1782270546a10077, /*  453 */
128'h862602e6446397c285b6300008378f95, /*  454 */
128'h30838287b823300017b70405aa1ff0ef, /*  455 */
128'h610101135f8134838526600134036081, /*  456 */
128'hbc2306a126050008380300d788338082, /*  457 */
128'he42643c0e8220c2007b71101b7e1ff06, /*  458 */
128'h16938304b703300014b747812401ec06, /*  459 */
128'h0485051300009517e7990206c1630337, /*  460 */
128'h64a2644260e2c3c00c2007b727b030ef, /*  461 */
128'hf0227179bfc14785eb9ff0ef80826105, /*  462 */
128'he78585930000a597461184ae8432ec26, /*  463 */
128'he30787930000a797099050eff4060068, /*  464 */
128'h88930000a89785a6862247b20007a803, /*  465 */
128'ha51704500693e1a757030000a717e168, /*  466 */
128'h740270a285228d4ff0efe22505130000, /*  467 */
128'h15428d5d05220085579b8082614564e2, /*  468 */
128'h8fd966c10185579b0185171b80829141, /*  469 */
128'h0085151b8fd98f750085571bf0068693, /*  470 */
128'h07b7715d808225018d5d8d7900ff0737, /*  471 */
128'h04b005134585460100740207879b0700, /*  472 */
128'hc63eec56f052f44ef84afc26e0a2e486, /*  473 */
128'h30eff8250513000095178a2a023070ef, /*  474 */
128'h99975ae14401d9e484930000a49719d0, /*  475 */
128'h854e85a2028a863b4919f7a989930000, /*  476 */
128'h0ff6761300ca56330286061b04852405, /*  477 */
128'ha5974611ff2410e3167030effec48fa3, /*  478 */
128'ha59746097a4050ef0048d64585930000, /*  479 */
128'hf0ef4512794050ef0028d52585930000, /*  480 */
128'h0087179bf0060613010006374722f47f, /*  481 */
128'h300016b78fd915020ff777138ff18321, /*  482 */
128'hb78380f6b42393c180a6b02317c29101, /*  483 */
128'h82f6b42347a1640660a68086b7838006, /*  484 */
128'h17b7808261616ae27a0279a2794274e2, /*  485 */
128'h0080073771398087b5838007b6033000, /*  486 */
128'hec4ef04af426f822fc068f4d91c115c2, /*  487 */
128'h05130000951780e7b423e05ae456e852, /*  488 */
128'ha797cbd747030000a7170b9030efec65, /*  489 */
128'ha697caf848030000a817cb67c7830000, /*  490 */
128'ha597c9b646030000a617ca46c6830000, /*  491 */
128'h30efe9a5051300009517c925c5830000, /*  492 */
128'h448100044783c7e404130000a41707d0, /*  493 */
128'hc6f708230000a717c58989930000a997, /*  494 */
128'ha7176a89c4ca0a130000aa1700144783, /*  495 */
128'h193700262b3700244783c4f70da30000, /*  496 */
128'ha71700344783c4f704230000a7173000, /*  497 */
128'h09230000a71700444783c2f70ea30000, /*  498 */
128'ha797c2f703a30000a71700544783c2f7, /*  499 */
128'ha797be07a9230000a797be079f230000, /*  500 */
128'ha797be07a7230000a797be07ad230000, /*  501 */
128'h8522e78d0009a783e4a9be07a1230000, /*  502 */
128'h03379713830937835a0b0493f2ffe0ef, /*  503 */
128'hfc075de3033797138309378302074563, /*  504 */
128'h4501dff154fd000a2783bfc5c0dff0ef, /*  505 */
128'hb7e9bf3ff0efbfc1710a849377d050ef, /*  506 */
128'h8f5d07a20005470300154783b7d914fd, /*  507 */
128'h8d5d05628fd907c20035450300254783, /*  508 */
128'hc703808200f61363367d57fd80822501, /*  509 */
128'h367d57fdb7f5fee50fa3058505050005, /*  510 */
128'h495cbfcd050500b50023808200f61363, /*  511 */
128'hcfa500958413e04ae426ec06e8221101, /*  512 */
128'h48a5481586ca02000513478101853903, /*  513 */
128'h00a70e6327850006c703462d02e00313, /*  514 */
128'h00640023011795630e50071301071463, /*  515 */
128'h4783fcc79ee30685040500e400230405, /*  516 */
128'hf59ff0ef00f5842384ae01c9051300b9, /*  517 */
128'h8fd90087979b0189470301994783c088, /*  518 */
128'h0087979b016947030179478300f49223, /*  519 */
128'h64a2644260e20004002300f493238fd9, /*  520 */
128'h02000593cf99873e611c808261056902, /*  521 */
128'h00c6986302d5fc630007468303a00613, /*  522 */
128'hb7dd0705a00d577d00d7066300178693, /*  523 */
128'h0ff6f593fd06869b577d46050007c683, /*  524 */
128'h8082853ae11c0006871b078900b66663, /*  525 */
128'hcb85611cc915bfd5aa8747030000a717, /*  526 */
128'h9063008557030067d683c70d0007c703, /*  527 */
128'h77933c4060ef0017c503e406114102e6, /*  528 */
128'h45258082014160a24525c39145010015, /*  529 */
128'h0087979b468d01a5c70301b5c7838082, /*  530 */
128'hc6830155c78300d51d630007079b8f5d, /*  531 */
128'h27818fd90107979b8fd50087979b0145, /*  532 */
128'hf4065904e44eec26f02271798082853e, /*  533 */
128'h468500154503842a03450993e052e84a, /*  534 */
128'h4c58505ce1312501352060ef85ce8626, /*  535 */
128'h70a2450100e7eb6340f487bb00040223, /*  536 */
128'h4903808261456a0269a2694264e27402, /*  537 */
128'h4685001445034c5cff2a74e34a050034, /*  538 */
128'h4505b7e5397d310060ef85ce86269cbd, /*  539 */
128'h80824501f8dff06fc39900454783b7f9, /*  540 */
128'h87634401e04ae426ec06e8221101591c, /*  541 */
128'hec190005041bfddff0ef892e84aa02b7, /*  542 */
128'h298060ef03448593864a46850014c503, /*  543 */
128'h60e285220324a823597d4405c1192501, /*  544 */
128'hec06e822110180826105690264a26442, /*  545 */
128'hf0ef842ad91c0005022357fde04ae426, /*  546 */
128'h45092324470323344783e52d2501fa3f, /*  547 */
128'h4107d79b776d0107979b8fd90087979b, /*  548 */
128'hd59ff0ef06a4051302f71f63a5570713, /*  549 */
128'h00544537fff50913010005370005079b, /*  550 */
128'h051300978c6345010127f7b314650493, /*  551 */
128'h35338d05012575332501d33ff0ef0864, /*  552 */
128'h450d80826105690264a2644260e200a0, /*  553 */
128'hf052fc26e0a2e486f44ef84a715dbfcd, /*  554 */
128'hf0ef8932852e89aa00053023e85aec56, /*  555 */
128'h0000a7970035171302054e6347addd9f, /*  556 */
128'hb023c01547b184aa638097ba8ac78793, /*  557 */
128'h1e2060ef00144503cb85000447830089, /*  558 */
128'h47a9c111891100090563e38d00157793, /*  559 */
128'h6b426ae27a0279a2794274e2640660a6, /*  560 */
128'h00a3000400230ff4f51380826161853e, /*  561 */
128'h0463fb71478d001577130f4060ef00a4, /*  562 */
128'h4785ee1ff0ef85224581f56989110009, /*  563 */
128'h89a623a40a131fa40913848a04f51a63, /*  564 */
128'h2501c5bff0ef854ac7894501ffc94783, /*  565 */
128'h01048913ff2a14e30991094100a9a023, /*  566 */
128'hf0ef852285d6000a876345090004aa83, /*  567 */
128'h19634785470dfe9915e30491c10de9df, /*  568 */
128'hc1194a81f6e504e34785470db7bd00e5, /*  569 */
128'h0087979b03f4470304044783bfb947b5, /*  570 */
128'h11e3200007134107d79b0107979b8fd9, /*  571 */
128'he9b30089999b04a4478304b44983fef7, /*  572 */
128'h01342e230444490329811a09866300f9, /*  573 */
128'h69e30ff7f793012401a3fff9079b4705, /*  574 */
128'h079bfa0b03e30164012304144b03faf7, /*  575 */
128'h0454478304644a03ffc900fb77b3fffb, /*  576 */
128'h00fa77930144142300fa6a33008a1a1b, /*  577 */
128'h8d450085151b0474448304844503f3c1, /*  578 */
128'h979b2501042447030434478314050e63, /*  579 */
128'h004a571b2781033906bbdfb18fd90087, /*  580 */
128'h40c504bbf4c564e3873200d7063b9f3d, /*  581 */
128'h3933664119556905dd8d84ae0364d5bb, /*  582 */
128'h00ea873b490d00b673630905165500b9, /*  583 */
128'hd05c03542023cc04d458015787bb2489, /*  584 */
128'hf0ef06040513f00a15e310e91263470d, /*  585 */
128'h0094d49b1ff4849b0024949bd408b17f, /*  586 */
128'hf8000793c45cc81c57fdee99e7e32481, /*  587 */
128'h47030654478308f91963478d00f402a3, /*  588 */
128'h4107d79b0107979b8fd90087979b0644, /*  589 */
128'hce5ff0ef8522001a859b06f71b634705, /*  590 */
128'h000402a32324470323344783e13d2501, /*  591 */
128'h4107d79b776d0107979b8fd90087979b, /*  592 */
128'ha99ff0ef0344051304f71263a5570713, /*  593 */
128'h051302f51763252787932501416157b7, /*  594 */
128'h272787932501614177b7a83ff0ef2184, /*  595 */
128'h0513c808a6dff0ef21c4051300f51c63, /*  596 */
128'h6327d78300009797c448a63ff0ef2204, /*  597 */
128'h132362f712230000971793c117c22785, /*  598 */
128'h0513b351478100042a230124002300f4, /*  599 */
128'h05440513b5b90005099ba33ff0ef0584, /*  600 */
128'h4789d41c9fb5e00a05e3b545a25ff0ef, /*  601 */
128'h029787bb478db7010014949b00f91563, /*  602 */
128'hec06e8221101bdc59cbd0017d79b8885, /*  603 */
128'h00044703ed692501bffff0ef842ae426, /*  604 */
128'h0af71b634785005447030cf71063478d, /*  605 */
128'ha01ff0ef852645812000061303440493, /*  606 */
128'h22f409a3faa0079322f4092305500793, /*  607 */
128'h0610079302f40aa302f40a2305200793, /*  608 */
128'h0ba304100713481c20f40da302f40b23, /*  609 */
128'h571b0107571b0107971b20e40d2302e4, /*  610 */
128'hd79b0107d71b20e40ea320f40e230087, /*  611 */
128'h971b501020e40f23445c20f40fa30187, /*  612 */
128'h0693001445030087571b0107571b0107, /*  613 */
128'h0107d71b260522e400a322f400230720, /*  614 */
128'h22e4012320d40ca320d40c230187d79b, /*  615 */
128'h02a363d050ef85a64685d81022f401a3, /*  616 */
128'h2501631050ef45814601001445030004, /*  617 */
128'h4d1c8082610564a2644260e200a03533, /*  618 */
128'h55480025458300f6f96337f9ffe5869b, /*  619 */
128'hf76347858082450180829d2d02d585bb, /*  620 */
128'he44eec26f022f406e84a71794d180eb7, /*  621 */
128'h0c63842e46890005470302e5f963892a, /*  622 */
128'h0015d49b00f71e6308d70e63468d06d7, /*  623 */
128'h2501ac7ff0ef9dbd0094d59b9cad515c, /*  624 */
128'h853e69a2694264e2740270a257fdc911, /*  625 */
128'h0099d59b0014899b0249278380826145, /*  626 */
128'hf0ef0344c483854a9dbd94ca1ff4f493, /*  627 */
128'h03494783994e1ff9f993f5792501a93f, /*  628 */
128'h6505bf658391c0198fc50087979b8805, /*  629 */
128'hf0ef9dbd0085d59b515cbf458fe9157d, /*  630 */
128'h99221fe474130014141bfd592501a63f, /*  631 */
128'hb7598fc90087979b0349450303594783, /*  632 */
128'hf9352501a39ff0ef9dbd0075d59b515c, /*  633 */
128'hf0ef954a034505131fc575130024151b, /*  634 */
128'h853e4785b76517fd2501100007b7807f, /*  635 */
128'hec4ef426fc06f04a4540f82271398082, /*  636 */
128'h00f41c63892a478500b51523e456e852, /*  637 */
128'h6aa26a4269e2790274a2744270e24509, /*  638 */
128'he02184aefee474e34f98611c80826121, /*  639 */
128'hd703eb15579800e69463470d0007c683, /*  640 */
128'hd79bd171008928235788fce4f7e30087, /*  641 */
128'h03478793049688bd000937839d3d0044, /*  642 */
128'h8722b75d450100993c2300a92a2394be, /*  643 */
128'h000935034a8509925a7d843a0027c983, /*  644 */
128'hf0efbf752501e59ff0ef0134f66385a2, /*  645 */
128'h3783f68afbe301440c630005041be6ff, /*  646 */
128'h4505bfc1413484bbf6f476e34f9c0009, /*  647 */
128'h842aec06e426e822110100a55583b78d, /*  648 */
128'hf0ef6008484ce4950005049bf33ff0ef, /*  649 */
128'h4581020006136c08ec990005049b933f, /*  650 */
128'h4705601c00e7802357156c1cf3cff0ef, /*  651 */
128'h8082610564a28526644260e200e78223, /*  652 */
128'he456ec4ef04af426f822fc06e8527139, /*  653 */
128'h0af5f063498984aa4d1c16ba75634a05, /*  654 */
128'h470d0ae78f63842e8932470900054783, /*  655 */
128'h0a3b515c0015da1b154794630ee78863, /*  656 */
128'h0005099b8b9ff0ef9dbd009a559b00ba, /*  657 */
128'h7a130ff97793001a0a9b880506099663, /*  658 */
128'h16c166850347c783014487b3cc191ffa, /*  659 */
128'h0ff7f7938fd98ff50049179b00f7f713, /*  660 */
128'hd59b50dc00f48223478502fa0a239a26, /*  661 */
128'h9f630005099b86bff0ef9dbd8526009a, /*  662 */
128'h0ff979130049591bc40d1ffafa930009, /*  663 */
128'h744270e200f482234785032a8a239aa6, /*  664 */
128'h808261216aa26a4269e2790274a2854e, /*  665 */
128'h00f979130089591b0347c783015487b3, /*  666 */
128'h9dbd0085d59b515cb7e90127e9339bc1, /*  667 */
128'h0014141bfc0992e30005099b811ff0ef, /*  668 */
128'h591b0109191b03240a2394261fe47413, /*  669 */
128'hbf790144822303240aa30089591b0109, /*  670 */
128'h0005099bfd8ff0ef9dbd0075d59b515c, /*  671 */
128'h03440a931fc474130024141bf80996e3, /*  672 */
128'h8d71f00006372501da0ff0ef85569aa6, /*  673 */
128'h0a230107d79b94260109179b01256933, /*  674 */
128'h591b0109579b00fa80a30087d79b0324, /*  675 */
128'hbf3d4989b745012a81a300fa81230189, /*  676 */
128'he456e852f04af822fc06ec4ef4267139, /*  677 */
128'h4d1c04090a6300c52903e19d89ae84aa, /*  678 */
128'h636324054c9c5afd4a05844a04f97763, /*  679 */
128'h041bc43ff0efa8214401052a606304f4, /*  680 */
128'h547d00f41d6357fd0887f86347850005, /*  681 */
128'h6aa26a4269e2790274a2744270e28522, /*  682 */
128'h4905b7d5faf47ee3894e4c9c80826121, /*  683 */
128'hc9012501c05ff0ef852685a24409bf55, /*  684 */
128'h0637b76dfb2411e305450863fd5507e3, /*  685 */
128'he9052501de9ff0ef852685a2167d1000, /*  686 */
128'h37fdfae783e3577dc4c0489c02099063, /*  687 */
128'hbf4900f482a30017e7930054c783c89c, /*  688 */
128'h4785dd612501dbbff0ef852685ce8622, /*  689 */
128'h00a55903f04a7139bfad4405f6f50fe3, /*  690 */
128'he852ec4ef426030917932905f822fc06, /*  691 */
128'h790274a2744270e24511eb9993c1e456, /*  692 */
128'h7993d7ed495c808261216aa26a4269e2, /*  693 */
128'h61082785480c00099d63842a8a2e00f9, /*  694 */
128'hfcf775e30009071b00855783e18dc85c, /*  695 */
128'hec1c97ce03478793012415230996601c, /*  696 */
128'hfab337fd00495a9b00254783bf5d4501, /*  697 */
128'h47850005049bb27ff0effc0a9fe30157, /*  698 */
128'h450500f4946357fdbf4945090097e463, /*  699 */
128'h480cf60a0ee306f4e0634d1c6008b761, /*  700 */
128'h8be34785d4bd451d0005049be81ff0ef, /*  701 */
128'h2501dd8ff0ef6008fcf48de357fdfcf4, /*  702 */
128'hf0ef034505134581200006136008f579, /*  703 */
128'h2823aa5ff0ef855285a600043a03beef, /*  704 */
128'h591c00faed630025478360084a0502aa, /*  705 */
128'ha83ff0ef85a6c8046008d91c415787bb, /*  706 */
128'hf1412501d1cff0ef01450223b7b9c848, /*  707 */
128'hf8227139b7e9db1c27855b1c2a856018, /*  708 */
128'hc783e05ae456e852ec4ef04afc06f426, /*  709 */
128'h071300e78663842e84aa02f007130005, /*  710 */
128'h000447030004a62304050ce7906305c0, /*  711 */
128'h099305c00a9302f00a130ae7fc6347fd, /*  712 */
128'h0d5780630d478263000447834b2102e0, /*  713 */
128'hb40ff0ef854a02000593462d0204b903, /*  714 */
128'h00144783013900230d37926300044783, /*  715 */
128'h0024478300f900a302e007930b379063, /*  716 */
128'h02000793943a09479763470d1b378e63, /*  717 */
128'h10632501adbff0ef8526458100f905a3, /*  718 */
128'h6c98e96d2501cdaff0ef608848cc1005, /*  719 */
128'h709cef918ba100b74783c7e500074783, /*  720 */
128'hfff74603078507050cb78d6300b78593, /*  721 */
128'hdfdff0ef85264581fed608e3fff7c683, /*  722 */
128'hf0ef85264581b791c55c4bdc611cbf75, /*  723 */
128'h790274a2744270e20004bc232501a85f, /*  724 */
128'hbf1d0405808261216b026aa26a4269e2, /*  725 */
128'h12f6e06302000693f7578be3bf954709, /*  726 */
128'h478145a147014681b7ad02400793943a, /*  727 */
128'h0027e793a8dd0505a0d1486502000313, /*  728 */
128'ha06d268500e50023954a910102069513, /*  729 */
128'h00d515630e50069300094503c6ed4711, /*  730 */
128'hf7930027979b0165966300d900234695, /*  731 */
128'h0107671300b6946345850037f6930ff7, /*  732 */
128'h920116020087671300d7946346918bb1, /*  733 */
128'h709c4511bf654701bdfd00e905a39432, /*  734 */
128'h0047f713f4e518e34711c50500b7c783, /*  735 */
128'h03e30004bc230004a623cb890207f793, /*  736 */
128'hfbf58b91b73d4515fb0dbf154501e807, /*  737 */
128'h0007c503609cdbe58bc100b5c7836c8c, /*  738 */
128'h0027979b05659a63bdb9c4c8af2ff0ef, /*  739 */
128'h17020017061b873245ad46a10ff7f793, /*  740 */
128'hf94706e3f4e374e30007470397229301, /*  741 */
128'h0187151b02b6f263fd370ae3f95704e3, /*  742 */
128'hf18505130000851700054c634185551b, /*  743 */
128'hbd6d4519f11710e30008866300054883, /*  744 */
128'hf9f7051beea87ae30ff57513fbf7051b, /*  745 */
128'h77130017e7933701eea866e30ff57513, /*  746 */
128'h842ae44ee84aec26f0227179bdf90ff7, /*  747 */
128'he199484c49bd0e500913451184aef406, /*  748 */
128'h6c1ce1292501afaff0ef6008a0b1c90d, /*  749 */
128'h026303f7f79300b7c783c3210007c703, /*  750 */
128'h9a630017b79317e18bfd033780630327, /*  751 */
128'h614569a2694264e2740270a245010097, /*  752 */
128'h2a23d9452501c13ff0ef852245818082, /*  753 */
128'hec06e82245811101bfe54511b7cd0004, /*  754 */
128'h0e500493e50d250188fff0ef842ae426, /*  755 */
128'hc7836c1ced092501a8cff0ef6008484c, /*  756 */
128'hbcdff0ef85224585cb9900978d630007, /*  757 */
128'h644260e2451d00f513634791dd792501, /*  758 */
128'h842aec06e426e82211018082610564a2, /*  759 */
128'hf0ef6008484ce49d0005049bfa9ff0ef, /*  760 */
128'h4581020006136c08e0850005049ba42f, /*  761 */
128'h601c82aff0ef462d6c08700c84cff0ef, /*  762 */
128'h610564a28526644260e200e782234705, /*  763 */
128'h70a245098082450900b7ed6347858082, /*  764 */
128'h4d1c808261456a0269a2694264e27402, /*  765 */
128'h842ae052e44ee84af406ec26f0227179, /*  766 */
128'h00f4fa634c1c59fd4a05fcf5fde384ae, /*  767 */
128'h000914630005091bec8ff0ef852285a6, /*  768 */
128'h85a6460103390763fb490ce3bf754501, /*  769 */
128'h01378a63481cf15d25018afff0ef8522, /*  770 */
128'h00f402a30017e79300544783c81c2785, /*  771 */
128'h1028ec2a7139b7594505bf5d0009049b, /*  772 */
128'h0405426383eff0eff42ee432e82efc06, /*  773 */
128'h631800a78733050eb187879300009797, /*  774 */
128'h00070023c319676200070023c3196622, /*  775 */
128'h460100f618634785cb114501e39897aa, /*  776 */
128'h8082612170e22501a0eff0ef0828080c, /*  777 */
128'hf4cefca6e122e506f8ca7175bfe5452d, /*  778 */
128'h302314050d634925e42ee8daecd6f0d2, /*  779 */
128'h9d6ff0ef1028002c8a7984aa89b20005, /*  780 */
128'he4be1028083c65a2140910630005091b, /*  781 */
128'hf7934519e011e11964062501b6dff0ef, /*  782 */
128'h00f516634791c54dc3e101f9fa1301c9, /*  783 */
128'h6406e949008a6a132501e75ff0ef1028, /*  784 */
128'h02100713046007937aa2cfcd008a7793, /*  785 */
128'h000407a30004072300f40ca300f408a3, /*  786 */
128'h00e40c2300040ba300040b2300e40823, /*  787 */
128'h00040f2300040ea300040e23000405a3, /*  788 */
128'h4785fc9fe0ef85a2000ac50300040fa3, /*  789 */
128'h00040aa300040a2300040da300040d23, /*  790 */
128'h855685ce04098b6300fa82230005099b, /*  791 */
128'h39fd7522e9112501e3fff0ef030aab03, /*  792 */
128'h892ac90d250183aff0ef0135262385da, /*  793 */
128'h81e30049f993e3d98bc500b44783a895, /*  794 */
128'h0107f71300b44783f565a0854921f609, /*  795 */
128'h7793e3ad8b85000984630029f993e72d, /*  796 */
128'h0309a78385a279a2020a6a13c399008a, /*  797 */
128'h0009c503000485a3d09c01448523f480, /*  798 */
128'hd783dbbfe0ef01c40513c8c8f33fe0ef, /*  799 */
128'h0134b0230004ae230004a623c8880069, /*  800 */
128'h79a6794674e6854a640a60aa00f49423, /*  801 */
128'h491db7e54911808261496b466ae67a06, /*  802 */
128'hf4a6fc86e4d6e8d2eccef8a27119b7d5, /*  803 */
128'ha023ec6ef06af466f862fc5ee0daf0ca, /*  804 */
128'h099be91fe0ef8ab6e4328a2e842a0006, /*  805 */
128'h899bc39d662200b44783000998630005, /*  806 */
128'h6a4669e6790674a6854e744670e60007, /*  807 */
128'h61096de27d027ca27c427be26b066aa6, /*  808 */
128'h01042903160789638b8500a447838082, /*  809 */
128'h0006091b00f67463893e40f907bb445c, /*  810 */
128'h4458fa090ce35c7d03040b1320000b93, /*  811 */
128'h478300975c9b6008120790631ff77793, /*  812 */
128'h020c99630ffcfc930197fcb337fd0025, /*  813 */
128'h00f405a3478900a7ec6347854848eb11, /*  814 */
128'h1763b7e52501bd6ff0ef4c0cb7414989, /*  815 */
128'h3d83cc08b7a5498500f405a347850185, /*  816 */
128'h861bd5792501b98ff0ef856e4c0c0004, /*  817 */
128'h8d3a0007849b00a6073b0099579b000c, /*  818 */
128'h419684bb00f6f4639fb1002dc683c4b5, /*  819 */
128'h250114a050ef85d2863a86a6001dc503, /*  820 */
128'h07bb4c48c3850407f79300a44783f94d, /*  821 */
128'h0613910115020097951b0097fc6341a5, /*  822 */
128'h97930094949bc5ffe0ef955285da2000, /*  823 */
128'hc45c9fa54099093b445c9a3e93810204, /*  824 */
128'h01634c50b70500faa0239fa5000aa783, /*  825 */
128'h001dc503c38d0407f79300a4478304e6, /*  826 */
128'h4783f1392501110050efe43a85da4685, /*  827 */
128'h4685601c00f40523fbf7f793672200a4, /*  828 */
128'hf11525010bc050ef85da0017c503863a, /*  829 */
128'h87bb1ff5f5930009049b444c01a42e23, /*  830 */
128'h8626030585930007849b0127f46340bb, /*  831 */
128'h7159b59d499dbf9dbd1fe0ef855295a2, /*  832 */
128'hf85aeca6f486fc56e0d2e4cee8caf0a2, /*  833 */
128'h842a0006a023e46ee86aec66f062f45e, /*  834 */
128'h97630005099bcb5fe0ef8ab689328a2e, /*  835 */
128'h740670a60007899bc39d00b447830009, /*  836 */
128'h7ba27b427ae26a0669a6694664e6854e, /*  837 */
128'h00a44783808261656da26d426ce27c02, /*  838 */
128'h04f76c630127873b445c18078f638b89, /*  839 */
128'h0409046344585c7d03040b1320000b93, /*  840 */
128'h478300975c9b6008140793631ff77793, /*  841 */
128'h040c9a630ffcfc930197fcb337fd0025, /*  842 */
128'h478902e798634705cb914581485cef01, /*  843 */
128'h079bd86ff0ef4c0cb759498900f405a3, /*  844 */
128'h00a4478312f76a634818445cf3fd0005, /*  845 */
128'h478501879763b79500f405230207e793, /*  846 */
128'hc85ce311cc1c4858bf99498500f405a3, /*  847 */
128'h46854c50601cc38d0407f79300a44783, /*  848 */
128'h4783f96925017b1040ef85da0017c503, /*  849 */
128'h4c0c00043d8300f40523fbf7f79300a4, /*  850 */
128'h579b000c869bd159250197cff0ef856e, /*  851 */
128'hc703c4b58d320007849b00a6863b0099, /*  852 */
128'h001dc503419704bb00f774639fb5002d, /*  853 */
128'h87bb4c4cf1512501763040ef85d286a6, /*  854 */
128'h0613918115820097959b0297f26341a5, /*  855 */
128'hf79300a44783a4ffe0ef855a95d22000, /*  856 */
128'h9381020497930094949b00f40523fbf7, /*  857 */
128'h000aa783c45c9fa54099093b445c9a3e, /*  858 */
128'h481800c78e634c5cbdd100faa0239fa5, /*  859 */
128'h40ef85da4685001dc50300e7fa63445c, /*  860 */
128'h0009049b444801a42e23fd0925016c70, /*  861 */
128'h0007849b0127f46340ab87bb1ff57513, /*  862 */
128'h47839dbfe0ef952285d2862603050513, /*  863 */
128'hb5f9c81cbf4100f405230407e79300a4, /*  864 */
128'hacffe0ef842ae406e0221141bd2d499d, /*  865 */
128'hf793cf690207f71300a44783e1752501, /*  866 */
128'h05930017c50346854c50601cc3950407, /*  867 */
128'hf79300a44783ed552501685040ef0304, /*  868 */
128'h2501b77fe0ef6008500c00f40523fbf7, /*  869 */
128'h00e785a30207671300b7c703741ce15d, /*  870 */
128'h8e230086d69b0106d69b0107169b4818, /*  871 */
128'h8f230187571b0107569b00d78ea300e7, /*  872 */
128'h00078ba300078b23485800e78fa300d7, /*  873 */
128'h8a2327010107571b0107169b00e78d23, /*  874 */
128'h8aa30087571b0107571b0107171b00e7, /*  875 */
128'hd69b00e78c23021007130106d69b00e7, /*  876 */
128'h892300e78ca300d78da3046007130086, /*  877 */
128'hfdf7f793600800a44783000789a30007, /*  878 */
128'h014160a2640200f50223478500f40523, /*  879 */
128'h114180820141640260a24505ebbfe06f, /*  880 */
128'h8522e9012501effff0ef842ae406e022, /*  881 */
128'h640260a200043023e11925019cbfe0ef, /*  882 */
128'h95bfe0efec060028e42a110180820141, /*  883 */
128'h60e2450144a782230000879700054a63, /*  884 */
128'h002c4601e42a7159bfe5452d80826105, /*  885 */
128'h0005041bb3bfe0efeca6f486f0a21028, /*  886 */
128'h041bcd2ff0efe4be1028083c65a2ec19, /*  887 */
128'h8522cbd8575277a2e9916586e41d0005, /*  888 */
128'h8bc100b5c7838082616564e6740670a6, /*  889 */
128'hb7c5c8c897bfe0ef0004c50374a2cb99, /*  890 */
128'he42afca67175bfd94415fcf41ee34791, /*  891 */
128'h84ae00050023f0d2f4cef8cae122e506, /*  892 */
128'h081ce5292501acdfe0ef1828002c4601, /*  893 */
128'hc2be02f009934bdc597d842677e2ecbe, /*  894 */
128'h00008717e50567a24501040a12634a16, /*  895 */
128'h03a0071300e780230307071b38c74703, /*  896 */
128'h00e7812302f007130e94186300e780a3, /*  897 */
128'h79a6794674e6640a60aa00078023078d, /*  898 */
128'h2501f89fe0ef18284585808261497a06, /*  899 */
128'h77e2f5552501e6eff0ef18284581fd45, /*  900 */
128'h18284581c2aa8cdfe0ef0007c50365c6, /*  901 */
128'he48ff0ef18284581f9492501f63fe0ef, /*  902 */
128'h8a7fe0ef0007c50365c677e2e1052501, /*  903 */
128'h2501a9eff0ef1828458101450e632501, /*  904 */
128'h100cb7594509f8e516e367a24711dd61, /*  905 */
128'h10949301020797134781f5cfe0ef1828, /*  906 */
128'h04e462630037871beb05fc9747039736, /*  907 */
128'h0206961300e586bb40f405bbfff7871b, /*  908 */
128'h8023fff7c79301271a6396b2920166a2, /*  909 */
128'h920102071613b7c12785b7319c3d0136, /*  910 */
128'hb7e900c68023377dfc964603962a1088, /*  911 */
128'h973692810204169367220789bddd4545, /*  912 */
128'hfe9465e3fee78fa32405078500074703, /*  913 */
128'he852ec4efc06f04af426f8227139b709, /*  914 */
128'h17630005091bfb4fe0ef84ae842ae456, /*  915 */
128'h744270e20007891bcf8900b447830009, /*  916 */
128'h808261216aa26a4269e2790274a2854a, /*  917 */
128'h84bae3918b8900a44783009777634818, /*  918 */
128'hfcf778e34818445ce4bd000426234458, /*  919 */
128'hbf7d00f405230207e79300a44783c81c, /*  920 */
128'hfc960ee34c50d3e51ff7f793445c4481, /*  921 */
128'h601cc3850407f7930304099300a44783, /*  922 */
128'hed51250130f040ef0017c50385ce4685, /*  923 */
128'h4685601c00f40523fbf7f79300a44783, /*  924 */
128'hed3525012bd040ef85ce0017c5038626, /*  925 */
128'hc7290097999b002547836008bf59cc44, /*  926 */
128'hed630337563b0336d6bbfff4869b377d, /*  927 */
128'h9c9dc45c27814c0c8ff9413007bb02c6, /*  928 */
128'hc45c9fa5445c0499ea634a855a7dd1c1, /*  929 */
128'hcd112501c87fe0ef6008d7b51ff4f793, /*  930 */
128'h814ff0efe595484cbfb19ca90094d49b, /*  931 */
128'h00f405a3478900f5976347850005059b, /*  932 */
128'h00f405a3478500f5976357fdbded4909, /*  933 */
128'h600800a44783b765cc0cc84cb5ed4905, /*  934 */
128'h84cee5990005059bfddfe0efcb818b89, /*  935 */
128'hfee3fd4588e30005059bc4bfe0efbf69, /*  936 */
128'h84bbcc0c445cfaf5fae34f9c601cfaba, /*  937 */
128'hf822fc067139b7bdc45c013787bb4134, /*  938 */
128'hfe6fe0ef0828002c4601842ac52de42e, /*  939 */
128'hf01c101ce01c852265a267e2e1152501, /*  940 */
128'h00b5c783cd996c0ce529250197cff0ef, /*  941 */
128'hc50367e2a02d000430234515e7898bc1, /*  942 */
128'hd7838522458167e2c448e30fe0ef0007, /*  943 */
128'h0be347912501cbdfe0ef00f414230067, /*  944 */
128'hbfdd452580826121744270e2f971fcf5, /*  945 */
128'h842ae406e0221141b7c1fcf501e34791, /*  946 */
128'h640260a200043023e1192501dbafe0ef, /*  947 */
128'h842af406e84aec26f022717980820141, /*  948 */
128'h00091f63e8890005049bd98fe0ef892e, /*  949 */
128'h740270a20005049bc5ffe0ef85224581, /*  950 */
128'h4581022430238082614564e269428526, /*  951 */
128'h2a2302f5136347912501b32ff0ef8522, /*  952 */
128'he0ef85224581c68fe0ef852285ca0004, /*  953 */
128'hbf7d00042a2300f5166347912501f8bf, /*  954 */
128'h460184aee42aeca67159bf6584aad16d, /*  955 */
128'h0005041bedafe0eff486f0a21028002c, /*  956 */
128'h041b872ff0efe4be1028083c65a2e00d, /*  957 */
128'he0ef102885a6c489cf816786e8010005, /*  958 */
128'h44198082616564e6740670a68522c10f, /*  959 */
128'h46018b2ee42af85a8432f0a27159bfcd, /*  960 */
128'hfc56e4cee8caeca6f486e0d28522002c, /*  961 */
128'h1c6300050a1be7cfe0efec66f062f45e, /*  962 */
128'h6263ffec871b481c01842c836000000a, /*  963 */
128'h694664e68552740670a600fb202302f7, /*  964 */
128'h61656ce27c027ba27b427ae26a0669a6, /*  965 */
128'h4481490902fb9f63478500044b838082, /*  966 */
128'h08632501a55fe0ef852285ca4a8559fd, /*  967 */
128'h63e329054c1c2485e111095508630935, /*  968 */
128'h00f402a30017e793c80400544783fef9, /*  969 */
128'h4981490110000ab7504cb74d009b2023, /*  970 */
128'h0015899b852200099e631afd4c094481, /*  971 */
128'h09930344091385cee9212501d10fe0ef, /*  972 */
128'h979b0009470300194783038b91632000, /*  973 */
128'h94e33cfd39f909092485e3918fd90087, /*  974 */
128'h75332501abcfe0efe02e854ab745fc0c, /*  975 */
128'h4a05b7c539f109112485e11165820155, /*  976 */
128'he426e8221101bfad8a2abfbd4a09b749, /*  977 */
128'he4910005049bbc4fe0ef842ae04aec06, /*  978 */
128'h8526644260e20007849bcb9100b44783, /*  979 */
128'h0027f71300a447838082610564a26902, /*  980 */
128'hc8180207e793fed772e348144458cf39, /*  981 */
128'h2501a58ff0ef484cef01600800f40523, /*  982 */
128'h4c0cbf7d84aa00a405a3c53900042a23, /*  983 */
128'h450502f9146357fd0005091b94dfe0ef, /*  984 */
128'h2501b37fe0ef167d100006374c0cb7dd, /*  985 */
128'h449db7e12501a1cff0ef85ca6008f979, /*  986 */
128'h6ae34d1c6008fcf900e345094785b769, /*  987 */
128'h4c50601cdba50407f79300a44783fcf9, /*  988 */
128'h25016ec040ef030405930017c5034685, /*  989 */
128'hb7b100f40523fbf7f79300a44783f55d, /*  990 */
128'hfca6e122e5061008002c4605e42a7175, /*  991 */
128'h1008081c65a2e9052501ca0fe0eff8ca, /*  992 */
128'hc78345196786e1052501e3bfe0efe0be, /*  993 */
128'h00b5c483c59975e2eb890207f79300b7, /*  994 */
128'h794674e6640a60aa451dcb810014f793, /*  995 */
128'h041bad8fe0ef00094503790280826149, /*  996 */
128'hfc878de301492783c89d88c1cc0d0005, /*  997 */
128'h00a8458996cfe0ef00a8100c02800613, /*  998 */
128'hf0ef00a84581f1612501951fe0efcaa2, /*  999 */
128'he0ef1008faf518e34791d94d2501836f, /* 1000 */
128'h2501f20fe0ef7502e411f15525019f5f, /* 1001 */
128'hb769d575250191cff0ef85a27502bf61, /* 1002 */
128'hed26f506f1221028002c4605e42a7171, /* 1003 */
128'hece6f0e2f4def8dafcd6e152e54ee94a, /* 1004 */
128'h65a21c0414630005041bbd0fe0efe8ea, /* 1005 */
128'h09630005041bd67fe0efe4be1028083c, /* 1006 */
128'h00b7c783441967a61af4176347911c04, /* 1007 */
128'hb45fe0ef4581752218079f630207f793, /* 1008 */
128'h16f90f6344094785180902630005091b, /* 1009 */
128'h041ba98fe0ef752216f90b63440557fd, /* 1010 */
128'h85220109549b85ca7422160414630005, /* 1011 */
128'h0c1b45812000061303440a13f6efe0ef, /* 1012 */
128'h855202000593462d898fe0ef85520005, /* 1013 */
128'h0109199b0ff4fb1347c1248188cfe0ef, /* 1014 */
128'h021007930109d99b02f40fa30104949b, /* 1015 */
128'h0ff97a9304f4062302e00b930104d49b, /* 1016 */
128'h04f406a30084d49b0089d99b04600793, /* 1017 */
128'h040405a30404052303740a2302000613, /* 1018 */
128'h049404a305640423053407a305540723, /* 1019 */
128'h05740aa3772280efe0ef0544051385d2, /* 1020 */
128'h9363571400d6166357d200074603468d, /* 1021 */
128'h0107d79b0107969b06f40723478100f6, /* 1022 */
128'hd79b0106d69b0107979b06f404232781, /* 1023 */
128'h04a306d407a30087d79b0086d69b0107, /* 1024 */
128'he0ef1028040b99634c8500274b8306f4, /* 1025 */
128'h85a3752247416786e8350005041bf59f, /* 1026 */
128'h8b230460071300e78c230210071300e7, /* 1027 */
128'h8da301578d2300e78ca300078ba30007, /* 1028 */
128'h00f50223478500978aa301678a230137, /* 1029 */
128'h001c0d1b7522a82d0005041bd5afe0ef, /* 1030 */
128'h0005041b8dcfe0ef0195022303852823, /* 1031 */
128'hf61fd0ef3bfd8552458120000613ec09, /* 1032 */
128'he0ef85ca7522441db7498c6a0ffbfb93, /* 1033 */
128'h6a0a69aa694a64ea740a70aa8522f25f, /* 1034 */
128'h8082614d6d466ce67c067ba67b467ae6, /* 1035 */
128'h843284aee42aeca6f0a27159b7c54421, /* 1036 */
128'he13125019cafe0eff48610284605002c, /* 1037 */
128'he9152501b65fe0efe4be1028083c65a2, /* 1038 */
128'h6706e39d0207f79300b7c783451967a6, /* 1039 */
128'h027474138c658cbd752200b74783c30d, /* 1040 */
128'hc9efe0ef00f502234785008705a38c3d, /* 1041 */
128'he42a71718082616564e6740670a62501, /* 1042 */
128'he0efed26f122f5060088002c4605e02e, /* 1043 */
128'h008865a26786120796630005079b964f, /* 1044 */
128'h9a630005079baf7fe0eff0be083cf4be, /* 1045 */
128'h126302077713479900b7c70377861007, /* 1046 */
128'h102805ad46550e058e63479165e61007, /* 1047 */
128'he49fd0ef10a8008c02800613e55fd0ef, /* 1048 */
128'h10a865820c054d6347adf05fd0ef850a, /* 1049 */
128'h0ce793634711cbf90005079baadfe0ef, /* 1050 */
128'h464d648aefc50005079bdc5fe0ef10a8, /* 1051 */
128'h02814783e0dfd0ef00d4851302a10593, /* 1052 */
128'h00f40223478500f485a30207e7936406, /* 1053 */
128'h06f7086357d64736cbbd8bc100b4c783, /* 1054 */
128'h85220005059bf2dfd0ef85a600044503, /* 1055 */
128'hd0ef8522c5a547890005059bcaefe0ef, /* 1056 */
128'h468302e007936706efb10005079bfc3f, /* 1057 */
128'h06f707230107969b57d602f69d630557, /* 1058 */
128'hd79b0107979b06f7042327810107d79b, /* 1059 */
128'h04a30086d69b0106d69b0087d79b0107, /* 1060 */
128'he0ef008800f7022306d707a3478506f7, /* 1061 */
128'h079bb50fe0ef6506e7910005079be24f, /* 1062 */
128'h47a18082614d853e64ea740a70aa0005, /* 1063 */
128'h1028002c4605842ee42ae8a2711dbfcd, /* 1064 */
128'h1028083c65a2e9292501810fe0efec86, /* 1065 */
128'hc783451967a6e12925019abfe0efe4be, /* 1066 */
128'h00645703cb856786eb950207f79300b7, /* 1067 */
128'h570300e78ba30087571b00e78b237522, /* 1068 */
128'h478500e78ca30087571b00e78c230044, /* 1069 */
128'h6125644660e62501ad6fe0ef00f50223, /* 1070 */
128'h002c893284aee42ae0cae4a6711d8082, /* 1071 */
128'h0005041bf9bfd0efec86e8a208284601, /* 1072 */
128'h2501ca8fe0efd20208284581c4b9e051, /* 1073 */
128'h75c2e93d2501b8ffe0ef08284585e559, /* 1074 */
128'h061346ad00b48713ca1fd0ef8526462d, /* 1075 */
128'h0007869bfff6879bce89000700230200, /* 1076 */
128'hfec783e3177d0007c78397a693811782, /* 1077 */
128'h0005041be69fd0ef510c656202090a63, /* 1078 */
128'h84630005468304300793470d6562e015, /* 1079 */
128'hc29fd0ef953e034787930270079300e6, /* 1080 */
128'h6125690664a6644660e6852200a92023, /* 1081 */
128'h842abf550004802300f5156347918082, /* 1082 */
128'hec86e8a21028002c4605e42a711db7d5, /* 1083 */
128'h00010c2366a2ec550005041bee3fd0ef, /* 1084 */
128'heba10007c78397b69381020617934601, /* 1085 */
128'hbd6fe0efda0210284581ea2902000593, /* 1086 */
128'h2501abbfe0ef10284585e8410005041b, /* 1087 */
128'hd0ef082c462dc3dd650601814783e179, /* 1088 */
128'h0460071300e78c23021007136786bc7f, /* 1089 */
128'h2605a06100e78ca300078ba300078b23, /* 1090 */
128'h930102079713fff6079bbf45863eb74d, /* 1091 */
128'h8e2e4781082cfeb706e3000747039736, /* 1092 */
128'h051b27850006c70348b107f00e934365, /* 1093 */
128'h93411742370100a36c6391411542f9f7, /* 1094 */
128'hf863a82100070f1b9305051300007517, /* 1095 */
128'hf36d80826125644660e68522441900ee, /* 1096 */
128'hffe81be306080563000548030505bfcd, /* 1097 */
128'h5795a885078500c6802300fe06b3b7cd, /* 1098 */
128'h8fefe0ef00f502234785752200f50023, /* 1099 */
128'h0181478302f51b634791b7c10005041b, /* 1100 */
128'h6506f4450005041ba55fe0ef1028dbd5, /* 1101 */
128'h082c462d6506b07fd0ef458102000613, /* 1102 */
128'h842abf1900e785a347216786ae5fd0ef, /* 1103 */
128'he5e30585068500e58023f91780e3b751, /* 1104 */
128'h0007869b02000613472993811782f4c7, /* 1105 */
128'heaf71de30e50079301814703f8d771e3, /* 1106 */
128'h28830585230305452e0305052e83bf89, /* 1107 */
128'h040502938f2ae44ae826ec22110105c5, /* 1108 */
128'h4a8f8f9300005f97887687f2869a8646, /* 1109 */
128'h2583000fa38300b647338dfd00c6c5b3, /* 1110 */
128'ha3839db9007585bb0fc1008fa403000f, /* 1111 */
128'h581b0078159b0105883b004f2703ff4f, /* 1112 */
128'h9f3100f805bb0077073b0105e8330198, /* 1113 */
128'h171b9e39008f23838e358e6d00f6c633, /* 1114 */
128'h00c5873b008383bb8e590146561b00c6, /* 1115 */
128'h8ebd00cf24038ef900b7c6b300d383bb, /* 1116 */
128'h00d3e6b30116969b00f6d39b007686bb, /* 1117 */
128'h8f2d0007061b00d703bbffcfa4039fa1, /* 1118 */
128'h171b00a7579b9f3d8f2d9fa100777733, /* 1119 */
128'h87bb0003869b0005881b0f418f5d0167, /* 1120 */
128'h5f974ea5859300005597f45f17e300e3, /* 1121 */
128'hcf334ea2829300005297422f8f930000, /* 1122 */
128'hc383000faf0301e6c73300cf7f3300d7, /* 1123 */
128'h038a0005c70300ef0f3b0025c4030015, /* 1124 */
128'h00ef0f3b942a040a4318972a070a93aa, /* 1125 */
128'h581b9e3900581f1b010f083b004fa703, /* 1126 */
128'h9f3100f80f3b010f68330003a70301b8, /* 1127 */
128'h139b008fa7039e398e3d8e7501e7c633, /* 1128 */
128'h03bb00c3e63340189eb90176561b0096, /* 1129 */
128'hfff5c4838efd007f46b305919f3500cf, /* 1130 */
128'h94aa048affcfa7039eb90fc101e6c6b3, /* 1131 */
128'h843b8ec140980126d69b9fb900e6941b, /* 1132 */
128'h0077473301e777330083c7339fb900d3, /* 1133 */
128'h000f081b8f5d0147171b00c7579b9f3d, /* 1134 */
128'hf25599e300e407bb0004069b0003861b, /* 1135 */
128'h8393000053978ffa400f0f1300005f17, /* 1136 */
128'h040a00d7c2b30003a703010fc4033763, /* 1137 */
128'h9f21011fc4839f25400000c2c4b3942a, /* 1138 */
128'h0107083b40809e2194aa048a0043a403, /* 1139 */
128'h0107683301c8581b0048171b012fc483, /* 1140 */
128'h00e2c2b3048a00f8073b0083a4039e21, /* 1141 */
128'hc90300b6129b408000c2863b9ea194aa, /* 1142 */
128'h00c702bb03c100c2e6330156561b013f, /* 1143 */
128'h090a0056c6b300e7c6b3ffc3a4839c35, /* 1144 */
128'h24830106d69b9fa50106941b992a9ea1, /* 1145 */
128'h005747330007081b00d2843b8ec10009, /* 1146 */
128'h8f5d0177171b0097579b9f3d8f219fa5, /* 1147 */
128'h92e300e407bb0004069b0002861b0f91, /* 1148 */
128'h8f5dfff647132ee2829300005297f5f5, /* 1149 */
128'h022f4403021f43830002a70300d745b3, /* 1150 */
128'h418c95aa058a93aa038a020f45839f2d, /* 1151 */
128'h171b0107083b0042a5839f2d942a040a, /* 1152 */
128'h0107683301a8581b0003a5839e2d0068, /* 1153 */
128'h9e2d8e3d8e59fff6c6139db100f8073b, /* 1154 */
128'h400c9ead0166561b00a6139b0082a583, /* 1155 */
128'hc593023f44839ead00c703bb00c3e633, /* 1156 */
128'h9db5ffc2a4038db902c10075e5b3fff7, /* 1157 */
128'h9fa18dd50115d59b94aa00f5969b048a, /* 1158 */
128'h8f4dfff747130007081b00b385bb4080, /* 1159 */
128'h0157171b00b7579b9f3d007747339fa1, /* 1160 */
128'h00e587bb0005869b0003861b0f118f5d, /* 1161 */
128'h06bb00fe07bb010e883b6462f3ef9de3, /* 1162 */
128'hcd70cd34c97c0505282300c8863b00d3, /* 1163 */
128'hfc26e0a2715d653c80826105692264c2, /* 1164 */
128'hf413ec56f052e486e45ee85af44ef84a, /* 1165 */
128'h04000b13e53c893289ae84aa97b203f7, /* 1166 */
128'h9381178200078a1b408b07bb04000b93, /* 1167 */
128'h020ada93020a1a9300090a1b00f97463, /* 1168 */
128'h481020ef0144043b86560084853385ce, /* 1169 */
128'h4401852660bc0174176399d641590933, /* 1170 */
128'h7a0279a2794274e2640660a6b7c99782, /* 1171 */
128'hf0227179653c808261616ba26b426ae2, /* 1172 */
128'h8513e84af406e44eec26842a03f7f793, /* 1173 */
128'h0400099300e7802397a2f80007130017, /* 1174 */
128'h4581920116020006091b40a9863b449d, /* 1175 */
128'hfc1c078e643c0124f5633c9020ef9522, /* 1176 */
128'h740270a2fd24fde3450197828522603c, /* 1177 */
128'h8793000077978082614569a2694264e2, /* 1178 */
128'h879300007797e93c04053423639cf967, /* 1179 */
128'he13cb6c7879300000797ed3c639cf8e7, /* 1180 */
128'h20efec06850a46410505059311018082, /* 1181 */
128'h000065971ac686930000769747013bf0, /* 1182 */
128'h06890007c78300e107b345413c458593, /* 1183 */
128'h97ae000646038bbd962e0047d6130705, /* 1184 */
128'hfca71de3fef68fa3fec68f230007c783, /* 1185 */
128'h71758082610516e505130000751760e2, /* 1186 */
128'h6622f71ff0efe42ee5060808842ae122, /* 1187 */
128'h0808f01ff0ef0808e85ff0ef080885a2, /* 1188 */
128'h46a1595880826149640a60aaf83ff0ef, /* 1189 */
128'h0200071300d71763469100d70d63711c, /* 1190 */
128'h8082556dbfe50007ac2380824501cf98, /* 1191 */
128'h84ae842a200007b7ec06e426e8221101, /* 1192 */
128'h0880061309c686930000569702f50263, /* 1193 */
128'h33850513000065173285859300006597, /* 1194 */
128'h8082610564a2644260e2fc2419b030ef, /* 1195 */
128'h84ae200007b7ec06e4266100e8221101, /* 1196 */
128'h02f00613074686930000569702f40263, /* 1197 */
128'h2f850513000065172e85859300006597, /* 1198 */
128'h8082610564a2644260e2e00415b030ef, /* 1199 */
128'h84ae200007b7ec06e4266100e8221101, /* 1200 */
128'h03600613044686930000569702f40263, /* 1201 */
128'h2b850513000065172a85859300006597, /* 1202 */
128'h8082610564a2644260e2e40411b030ef, /* 1203 */
128'h842e200007b7ec06e8226104e4261101, /* 1204 */
128'h03e00613eec686930000769702f48263, /* 1205 */
128'h27850513000065172685859300006597, /* 1206 */
128'h64a2644260e2e880900114020db030ef, /* 1207 */
128'h07b7ec06e8226104e426110180826105, /* 1208 */
128'hea0686930000769702f48263842e2000, /* 1209 */
128'h00006517224585930000659704500613, /* 1210 */
128'h60e2ec8090011402097030ef23450513, /* 1211 */
128'he4266100e82211018082610564a26442, /* 1212 */
128'h0000569702f4026384ae200007b7ec06, /* 1213 */
128'h1e0585930000659704c00613f8c68693, /* 1214 */
128'h60e2f004053030ef1f05051300006517, /* 1215 */
128'he4266100e82211018082610564a26442, /* 1216 */
128'h0000569702f4026384ae200007b7ec06, /* 1217 */
128'h1a0585930000659705300613f5c68693, /* 1218 */
128'h60e2f404013030ef1b05051300006517, /* 1219 */
128'h00053983ec4e71398082610564a26442, /* 1220 */
128'h893284ae200007b7fc06f04af426f822, /* 1221 */
128'h0613f22686930000569702f984638436, /* 1222 */
128'h051300006517156585930000659705a0, /* 1223 */
128'h89890014159b67227c6030efe43a1665, /* 1224 */
128'h0034949b8dd9004979130029191b8b05, /* 1225 */
128'h02b9b8238dc5744270e288a10125e5b3, /* 1226 */
128'h7100e02211418082612169e2790274a2, /* 1227 */
128'hf7dff0efe40645818522460546814705, /* 1228 */
128'h4605468547058522f35ff0ef45818522, /* 1229 */
128'h60a2d97ff0ef45816008f67ff0ef4581, /* 1230 */
128'h4705e022e40611418082014145016402, /* 1231 */
128'h842a45810405302302053c2346054681, /* 1232 */
128'h45818522ef1ff0ef45818522f39ff0ef, /* 1233 */
128'h60a264026008f23ff0ef460546854705, /* 1234 */
128'he8226104e4261101d4dff06f01414581, /* 1235 */
128'h0000569702f48263842e200007b7ec06, /* 1236 */
128'h070585930000659706100613e4c68693, /* 1237 */
128'h904114426e2030ef0805051300006517, /* 1238 */
128'he42611018082610564a2644260e2fc80, /* 1239 */
128'h02f48263842e200007b7ec06e8226104, /* 1240 */
128'h0000659706800613e186869300005697, /* 1241 */
128'h69e030ef03c505130000651702c58593, /* 1242 */
128'h610564a2644260e2e0a08c7d17fd6785, /* 1243 */
128'h200007b7ec06e4266100e82211018082, /* 1244 */
128'h0613de2686930000569702f4026384ae, /* 1245 */
128'h051300006517fe6585930000659706f0, /* 1246 */
128'h610564a2644260e2e424658030efff65, /* 1247 */
128'hec06e426e82200053903e04a11018082, /* 1248 */
128'h0000569702f9026384ae842a200007b7, /* 1249 */
128'hfa0585930000659707600613dac68693, /* 1250 */
128'h04993c23612030effb05051300006517, /* 1251 */
128'h715980826105690264a2644260e2c844, /* 1252 */
128'hfc56e0d2e4cef486e8caeca67100f0a2, /* 1253 */
128'h0005d783020408a3ec66f062f45ef85a, /* 1254 */
128'h00c9051345814611d01ce03084b2892e, /* 1255 */
128'hbf5ff0ef458560080e049c636ca020ef, /* 1256 */
128'h16f99a6304043a03200007b700043983, /* 1257 */
128'h448d8b89c7090017f713448100492783, /* 1258 */
128'h000a09638cdd03243c234c1c4485e391, /* 1259 */
128'h47050144e493160786638b85008a2783, /* 1260 */
128'h85224581d71ff0ef8522458146054681, /* 1261 */
128'h0c1300005c17852200892583be1ff0ef, /* 1262 */
128'h00006a17852200095583c4fff0efd26c, /* 1263 */
128'hcbdff0ef852285a6c81ff0efecca0a13, /* 1264 */
128'h4581460546854705cf5ff0ef85224581, /* 1265 */
128'h852224058593000f45b7d27ff0ef8522, /* 1266 */
128'h0d89b583cd1ff0ef85224585e93ff0ef, /* 1267 */
128'heb7ff0ef25810015e593009899b78522, /* 1268 */
128'hefe9485ce8ca8a9300006a9768198993, /* 1269 */
128'h7b427ae26a0669a6694664e6740670a6, /* 1270 */
128'h852244cc8082616545016ce27c027ba2, /* 1271 */
128'h449cdf3ff0ef8522488cdb7ff0efe024, /* 1272 */
128'he683654100043883603cee079be38b85, /* 1273 */
128'h00ff0e37431147014781458163900107, /* 1274 */
128'h1f1b00064803ec0689e36e89f0050513, /* 1275 */
128'h060527810107e7b301e8183b07050037, /* 1276 */
128'h0187971b0187d81bf2e50067036316fd, /* 1277 */
128'h0087d79b01c878330087981b01076733, /* 1278 */
128'h1782170200be873b8fd98fe901076733, /* 1279 */
128'hb765470147812585e31c974693818375, /* 1280 */
128'h0000659714900613bc86869300005697, /* 1281 */
128'h41e030efdbc5051300006517dac58593, /* 1282 */
128'h3b7d20000bb78b4ebd6100c4e493bd85, /* 1283 */
128'h00006517bac5859300005597000b1d63, /* 1284 */
128'h096300043903b7116f6000efdac50513, /* 1285 */
128'h3de030ef855685d20f20061386e20179, /* 1286 */
128'h12048e6324818cfd4c81485c07093483, /* 1287 */
128'hc7817c1c00f76f630c89378302093703, /* 1288 */
128'h4581b6fff0ef85224581cc5cf9200793, /* 1289 */
128'h01442903c3950044f793b27ff0ef8522, /* 1290 */
128'hd47ff0ef85ca00896913ff3979138522, /* 1291 */
128'hf793680000efd4e505130000651785ca, /* 1292 */
128'h6913ff397913852201442903c3950084, /* 1293 */
128'h05130000651785cad1fff0ef85ca0049, /* 1294 */
128'h00043c83cfb50014f793658000efd4e5, /* 1295 */
128'hb186869300005697017c8c6303843903, /* 1296 */
128'hcba97c1c332030ef855685d209c00613, /* 1297 */
128'h9f630037f693470d02043c2300492783, /* 1298 */
128'h4591480d468100c90793018c871308e6, /* 1299 */
128'h01068763c3900086161bff8705136310, /* 1300 */
128'h0791872a2685c3988f518361ff873703, /* 1301 */
128'hc85c0027e793485ccbb5603cfeb690e3, /* 1302 */
128'h39036004cc9d4c858889c85c9bf9485c, /* 1303 */
128'h0613ab2686930000569701748c630404, /* 1304 */
128'h0963040430232b4030ef855685d20ca0, /* 1305 */
128'hb4dff0ef8522ef8d8b85008927830009, /* 1306 */
128'hc47ff0ef8522484cc85c9bf54c85485c, /* 1307 */
128'hdbd98b85bd95641020ef4505d80c8ee3, /* 1308 */
128'hb1dff0ef8522b77100f92623000cb783, /* 1309 */
128'h94be00093c830109648397a667a1bf41, /* 1310 */
128'h002c46218566639c00878913fa978de3, /* 1311 */
128'h41635535b7dd87ca0ca139a020efe43e, /* 1312 */
128'hf406e84aec26f02204800513717908b0, /* 1313 */
128'hcc1d5551842a1a4030ef892e84b2e44e, /* 1314 */
128'h89aa785010efa1e505130000551785a2, /* 1315 */
128'h4fe000efc1c5051300006517862285aa, /* 1316 */
128'hf40401242423e01c200007b702098b63, /* 1317 */
128'h740270a24501c45c4789cb990024f793, /* 1318 */
128'hd4fd450188858082614569a2694264e2, /* 1319 */
128'hbff9557d18c030ef8522b7e5c45c4785, /* 1320 */
128'h07b7f73ff06f20000537458146098082, /* 1321 */
128'h1141711c808225016108953e050e2000, /* 1322 */
128'h569702f40263200007b7e4066380e022, /* 1323 */
128'h85930000659734c006139ba686930000, /* 1324 */
128'h703c170030efb0e5051300006517afe5, /* 1325 */
128'h110180820141640260a2557de3914505, /* 1326 */
128'h85a24d3010efe42eec064501842ae822, /* 1327 */
128'h71797940006f6105468560e266226442, /* 1328 */
128'he052e44ee84aec26f022f40620000513, /* 1329 */
128'h30efb72505130000651784aa0aa030ef, /* 1330 */
128'h491010ef450144b010ef0001b5031b20, /* 1331 */
128'hb585051300006517681c206010ef842a, /* 1332 */
128'h05130000651706f445833f8000ef638c, /* 1333 */
128'hb605051300006517546c3e8000efb565, /* 1334 */
128'h4583583c3d2000ef91c115c20085d59b, /* 1335 */
128'hd69b0087d71bb56505130000651706c4, /* 1336 */
128'hf6930ff7f7930ff777130187d61b0107, /* 1337 */
128'h0513000065175c0c3a6000ef26010ff6, /* 1338 */
128'had05859300006597545c398000efb465, /* 1339 */
128'h051300006517abe5859300006597c789, /* 1340 */
128'h30efb425051300006517378000efb365, /* 1341 */
128'he0dfb0ef144585930000659774481020, /* 1342 */
128'he789a9a6061300006617584c19c42783, /* 1343 */
128'hb205051300006517df86061300006617, /* 1344 */
128'h4481ed5ff0ef84264581852633a000ef, /* 1345 */
128'hb209899300006997b20a0a1300006a17, /* 1346 */
128'h00ef855285a6e78901f4f79320000913, /* 1347 */
128'h819100f5f6132485854e0004458330c0, /* 1348 */
128'h051300006517fd249fe304052fa000ef, /* 1349 */
128'h69a2694264e2740270a22e8000ef0ce5, /* 1350 */
128'h0083b7830103b7038082614545016a02, /* 1351 */
128'hfe6393811782278540f707b30003b683, /* 1352 */
128'hb78300a7002300f3b8230017079300d7, /* 1353 */
128'hb7038082450180820007802345050103, /* 1354 */
128'hb7038f999201020596130103b7830083, /* 1355 */
128'hfff7059b00c6f5638e9dfff706930003, /* 1356 */
128'h00b6e6630103b70340a786bb87aa9d9d, /* 1357 */
128'h00d3b823001706938082852e00070023, /* 1358 */
128'h56634881bfe900d7002307850007c683, /* 1359 */
128'hc21906100693488540a0053be6810005, /* 1360 */
128'h061b385986ba4e250ff6f81304100693, /* 1361 */
128'h051b046e67630ff3751302b6733b0005, /* 1362 */
128'hfea68fa306850ff5751302b6563b0305, /* 1363 */
128'h02f5e9630300051340e685bbfe718532, /* 1364 */
128'h853b068500f6802302d0079300088763, /* 1365 */
128'h081b86ba2581000680230015559b40e6, /* 1366 */
128'h0685bf5d00a8053b808200b61b63fff5, /* 1367 */
128'h9381178240c807bbb7d92585fea68fa3, /* 1368 */
128'h0066802326050006c8830007c30397ba, /* 1369 */
128'h597d011cf0ca7119b7f1068501178023, /* 1370 */
128'h84b2e0dafc86e4d6e8d2eccef4a6f8a2, /* 1371 */
128'h0a1302500993f82af02ef42afc3e8436, /* 1372 */
128'hc50377a277420209591303000a9306c0, /* 1373 */
128'h9381178276820017079bc52d8f1d0004, /* 1374 */
128'hf0ef0201039304850135086304d7ff63, /* 1375 */
128'h4781048905450f630014c503bfe1e7bf, /* 1376 */
128'hf793fd07879bcb9d0004c78303551063, /* 1377 */
128'h04890014c503478100f6f36346a50ff7, /* 1378 */
128'h0580069302a6eb6306d50f6306400693, /* 1379 */
128'h70e6f55d08f509630630079304d50f63, /* 1380 */
128'h051b6b066aa66a4669e6790674a67446, /* 1381 */
128'h0713b74d048d0024c503808261090007, /* 1382 */
128'h1ee30700071300a76c6306e50e630730, /* 1383 */
128'h0713a00d46014685003800840b13f6e5, /* 1384 */
128'h0613f6e510e30780071302e500630750, /* 1385 */
128'h45c1001636134685003800840b13fa85, /* 1386 */
128'h0016b693003800840b13f8b50693a811, /* 1387 */
128'h03930005059be37ff0ef400845a94601, /* 1388 */
128'h039300044503a809ddbff0ef00280201, /* 1389 */
128'h0b13b5fd845ad93ff0ef00840b130201, /* 1390 */
128'h059b4db010ef85220124743360000084, /* 1391 */
128'h1034f436715db7f18522020103930005, /* 1392 */
128'he8dff0efe436e4c6e0c2fc3ef83aec06, /* 1393 */
128'h1014862ef436f032715d8082616160e2, /* 1394 */
128'he436e4c6e0c2fc3ef83aec0610000593, /* 1395 */
128'hfa32f62e710d8082616160e2e69ff0ef, /* 1396 */
128'hea22ee060808100005931234862afe36, /* 1397 */
128'h842ae3fff0efe436eec6eac2e6bee2ba, /* 1398 */
128'h80826135645260f28522129020ef0808, /* 1399 */
128'h45018302000303630087b303679c691c, /* 1400 */
128'h000047170205979304b7ee63479d8082, /* 1401 */
128'he822ec061101439c97ba83f951470713, /* 1402 */
128'h7540f55c08c52483795c878297bae426, /* 1403 */
128'h60e202f457b39381020497930c5010ef, /* 1404 */
128'hbfe97d5c808261054501e91c64a26442, /* 1405 */
128'hb7e9659c95aa058e05e135f1bfd9617c, /* 1406 */
128'h842ae406e02211418082557d8082557d, /* 1407 */
128'h0207b303679c681c00055e63ff5ff0ef, /* 1408 */
128'h45018302014160a26402852200030763, /* 1409 */
128'heb6347ad8082557d80820141640260a2, /* 1410 */
128'h953e817549c7879300004797150200a7, /* 1411 */
128'h691c808271c505130000551780826108, /* 1412 */
128'h02f1102347a1715d83020007b303679c, /* 1413 */
128'h0030e83ee42e078517824785d23e47d5, /* 1414 */
128'hfd3ff0efcc3ed402e486100c20000793, /* 1415 */
128'h00e6fe63400407374d148082616160a6, /* 1416 */
128'h34832301340323813083450180824501, /* 1417 */
128'h22813823dc0101138082240101132281, /* 1418 */
128'h22113c232291342385a2980101f10413, /* 1419 */
128'h47830a04c703f579f95ff0ef1a053483, /* 1420 */
128'h16630dd447830dd4c70302f71c630a04, /* 1421 */
128'hc70302f710630c0447830c04c70302f7, /* 1422 */
128'h0d440593461100f71a630e0447830e04, /* 1423 */
128'hb761fb600513d55156f010ef0d448513, /* 1424 */
128'h6ea020eff4063e800513842af0227179, /* 1425 */
128'hf0efc202c40200011023858a46018522, /* 1426 */
128'h85226cc020ef7d000513e509842af21f, /* 1427 */
128'h00f110234785717980826145740270a2, /* 1428 */
128'h6914c195842ac402c23ef406f0224785, /* 1429 */
128'h8ff58ff9f80787934ad4008007b74538, /* 1430 */
128'hc43e8fd98f55400006b78f75600006b7, /* 1431 */
128'hc43c47b2e119ec9ff0ef8522858a4601, /* 1432 */
128'h00f1102347b5711d80826145740270a2, /* 1433 */
128'h979bf852fc4ee0ca07c55783c23e47d5, /* 1434 */
128'hf456e4a6e8a26a056989fdf949370107, /* 1435 */
128'h8993080909134495c43e842e8aaaec86, /* 1436 */
128'he73ff0ef8556858a4601e00a0a13e009, /* 1437 */
128'h93630135f7b3c7891005f79345b2ed0d, /* 1438 */
128'h5785051300005517c78d0125f7b30547, /* 1439 */
128'h690664a6644660e6fba00513d4bff0ef, /* 1440 */
128'hfe04c6e334fd808261257aa27a4279e2, /* 1441 */
128'h20ef3e80051300f057630014079b347d, /* 1442 */
128'h051300005517fc8049e34501b7555d80, /* 1443 */
128'h19c52783bf7df9200513d09ff0ef54e5, /* 1444 */
128'h460147d5c42e00f1102347c17139e7a9, /* 1445 */
128'hde3ff0efc23e842af426fc06f822858a, /* 1446 */
128'h858a46014495cb918b891b842783c11d, /* 1447 */
128'h744270e2f8ed34fdc901dcdff0ef8522, /* 1448 */
128'h711d80824501bfd545018082612174a2, /* 1449 */
128'hf66384b6892a4785e8a2ec86e0cae4a6, /* 1450 */
128'h2783260102f1102302c9270347c906d7, /* 1451 */
128'h47850030cc3ee42e4755d432cf3108c9, /* 1452 */
128'h842ad75ff0efc83eca26d23a854a100c, /* 1453 */
128'h460102f1102347b10497f0634785e529, /* 1454 */
128'hc11dd55ff0efd23ed402854a100c47f5, /* 1455 */
128'h60e68522c43ff0ef4a85051300005517, /* 1456 */
128'h063bbf6147c580826125690664a66446, /* 1457 */
128'h7139b7c54401b7d50004841bb74d02f6, /* 1458 */
128'hce05e456e852ec4ef04af426f822fc06, /* 1459 */
128'h892a482010ef8ab684b28a2e4148842a, /* 1460 */
128'h00054d6391dfa0ef852200b44583c11d, /* 1461 */
128'h05130000551700b67a63014485b36810, /* 1462 */
128'h854a08c92583a0894481bd9ff0ef45e5, /* 1463 */
128'h0207e4030109378389a6f96decdff0ef, /* 1464 */
128'hf0ef854a85d6865286a2844e0089f363, /* 1465 */
128'h9a22408989b308c96783fc851ae3f01f, /* 1466 */
128'h8526744270e2fc0999e39aa202878433, /* 1467 */
128'h7139808261216aa26a4269e274a27902, /* 1468 */
128'h07b70086969bc23e47f500f110234799, /* 1469 */
128'hfc06f426f8228ed10106161b8edd0300, /* 1470 */
128'hc53ff0ef8526858a4601440dc43684aa, /* 1471 */
128'h744270e2d91ff0ef85263e800593e919, /* 1472 */
128'h01134d18bfcdfc79347d8082612174a2, /* 1473 */
128'h241134239fb923213823bffc07b7db01, /* 1474 */
128'h3ffc07372331342322913c2324813023, /* 1475 */
128'h84aa85a2980101f104131ce7f5634901, /* 1476 */
128'he7991a04b7831e051863892ac09ff0ef, /* 1477 */
128'h1a04b5031aa4b023766020ef20000513, /* 1478 */
128'h4783123010ef85a2200006131e050363, /* 1479 */
128'h04870713000047171cf76b6347210c04, /* 1480 */
128'hcc981ff78793400407b753b897ba078a, /* 1481 */
128'h07a68007071367050d44278300e7fd63, /* 1482 */
128'h49830a044783f8dc00d773630147d693, /* 1483 */
128'h4783e7810019f9938b8506f48f2309b4, /* 1484 */
128'h00098a6308f480a30b344783c7890e24, /* 1485 */
128'h06f48fa309c44783c7898b890a044783, /* 1486 */
128'hfcdc07c60c848613091407130e244783, /* 1487 */
128'h4783e0fc07c6468109d405130a844783, /* 1488 */
128'h9fad0105959b0087979b00074583fff7, /* 1489 */
128'h458300098c634685c39197aeffe74583, /* 1490 */
128'h07ce02b787b30dd4478302f585b30e04, /* 1491 */
128'h478304098f63fca714e30621070de21c, /* 1492 */
128'h0087171b0107979b468508d4470308e4, /* 1493 */
128'h02f707330e04470397ba08c447039fb9, /* 1494 */
128'h08b44783f8fc07ce02e787b30dd44783, /* 1495 */
128'h47039fb90107171b0187979b08a44703, /* 1496 */
128'h54d89fb9088447039fb90087171b0894, /* 1497 */
128'hc7898b850a044783f4fc07a6c319f4fc, /* 1498 */
128'h0af006134685ce81e3918bfd09c44783, /* 1499 */
128'h0af407a34785ed35e0bff0ef85264585, /* 1500 */
128'h00a6979bc7b98b850e0446830af44783, /* 1501 */
128'h0d44278300098663c79954dc08f4aa23, /* 1502 */
128'h02f686bb00a6969b0dd44783f8dc07a6, /* 1503 */
128'h2481308308f480230a74478308d4ac23, /* 1504 */
128'h39832301390323813483854a24013403, /* 1505 */
128'hd79b00a7d71b50fc8082250101132281, /* 1506 */
128'haa2302f707bb278527058bfd8b7d0057, /* 1507 */
128'h5c8020efd1691a04b503892abf4d08f4, /* 1508 */
128'h0113bf455929bf555951bf651a04b023, /* 1509 */
128'h3023229134232281382322113c23dc01, /* 1510 */
128'hc585468102b7e16302f5886347892321, /* 1511 */
128'h220139038526230134032381308354a9, /* 1512 */
128'h4705ffc5879b80822401011322813483, /* 1513 */
128'h892a45850b900613842e4685fef760e3, /* 1514 */
128'h258199f5ffe4059bf57184aad1fff0ef, /* 1515 */
128'h98dff0ef854a85a2980101f10413f1e9, /* 1516 */
128'h84aab75ddf400493f7d50b944783e519, /* 1517 */
128'h4783f022f406e44ee84aec267179b74d, /* 1518 */
128'h8edd892e9be10079f6930ff5f9930815, /* 1519 */
128'h57b5c519cc7ff0ef84aa45850b300613, /* 1520 */
128'hf0ef852685ca00091c6300f51e63842a, /* 1521 */
128'h8522013505a315e010ef8526842a875f, /* 1522 */
128'h01138082614569a2694264e2740270a2, /* 1523 */
128'h3023289134232881382328113c23d601, /* 1524 */
128'h3023275134232741382327313c232921, /* 1525 */
128'h3023259134232581382325713c232761, /* 1526 */
128'h07b74d180ac7e963478923b13c2325a1, /* 1527 */
128'hbfe787933ffc07b79f3dbff7879bbffc, /* 1528 */
128'heb63062505130000551784ae8b32892a, /* 1529 */
128'h00005517e7b90016779307e9460300e7, /* 1530 */
128'h30838522f8400413f96ff0ef08450513, /* 1531 */
128'h39832801390328813483290134032981, /* 1532 */
128'h3b8326013b0326813a8327013a032781, /* 1533 */
128'h3d8324013d0324813c8325013c032581, /* 1534 */
128'h000055170989270380822a0101132381, /* 1535 */
128'hf7bb060a81630045aa83db4505c50513, /* 1536 */
128'h5517cb8902ecf7bb0005ac83e79102ea, /* 1537 */
128'h2783bf415429f24ff0ef062505130000, /* 1538 */
128'h8c0a009c9c9be3994b8502eadabb02c9, /* 1539 */
128'h28834e114e85478189d6856200c48813, /* 1540 */
128'h551700030d6302e8f33b0017859b0008, /* 1541 */
128'h4a814c81b7c1ee4ff0ef05a505130000, /* 1542 */
128'h020880630065202302e8d33bb7f14b81, /* 1543 */
128'h00be96bbcb898b850107c78397a6078e, /* 1544 */
128'h05110821013309bb0ffbfb9300dbebb3, /* 1545 */
128'h000055178a09000b8963fbc596e387ae, /* 1546 */
128'hfe0a7a1302f10a13f00600e303c50513, /* 1547 */
128'h4603ee0519e3842af94ff0ef854a85d2, /* 1548 */
128'h9e3d0087979b0106161b09ea478309fa, /* 1549 */
128'h0000551785ce01367a63963e09da4783, /* 1550 */
128'h46830084c783b5c1e56ff0ef02c50513, /* 1551 */
128'h0fe6f9938b89c71989b60017f7130a7a, /* 1552 */
128'h0017059b4611450547010016e993c399, /* 1553 */
128'h0463001878130017581b4b189726070e, /* 1554 */
128'h999b0187979b0027571b00b517bb0208, /* 1555 */
128'he9b3c70d4189d99b4187d79b8b050189, /* 1556 */
128'h02d98263fcc592e3872e0ff9f99300f9, /* 1557 */
128'hfe05051300005517ef898b850a6a4783, /* 1558 */
128'hbfd100f9f9b3fff7c793b591370020ef, /* 1559 */
128'h0105051300005517cb898b8509ba4783, /* 1560 */
128'h0afa4783e20b02e3b51d547ddbaff0ef, /* 1561 */
128'hf0ef854a45850af006134685e3958b85, /* 1562 */
128'h979b0e0a47830afa07a34785e569a21f, /* 1563 */
128'h08c00d934d010880049308f92a2300a7, /* 1564 */
128'hf0ef854a458586260ff6f69301acd6bb, /* 1565 */
128'hffb492e32d210ff4f4932485ed499f1f, /* 1566 */
128'h86260ff6f693019ad6bb08f00d134c81, /* 1567 */
128'h0ff4f4932485e9359cbff0ef854a4585, /* 1568 */
128'h4c818aa609b00d934d61ffa492e32ca1, /* 1569 */
128'h0ff6f6930196d6bb45858656000c2683, /* 1570 */
128'h0ffafa932ca12a85e13999dff0ef854a, /* 1571 */
128'hfdb498e30c110ff4f493248dffac90e3, /* 1572 */
128'hed19975ff0ef854a458509c0061386de, /* 1573 */
128'h468501379b630a7a4783d4fb0de34785, /* 1574 */
128'hbb3d842a957ff0ef854a458509b00613, /* 1575 */
128'h842a945ff0ef854a45850a70061386ce, /* 1576 */
128'h810ff0ef842ae406e0221141b32ddd79, /* 1577 */
128'h000307630187b303679c681c00055e63, /* 1578 */
128'h640260a245058302014160a264028522, /* 1579 */
128'h4791f04af822fc06f426713980820141, /* 1580 */
128'h079304f592635529478500f5866384aa, /* 1581 */
128'h979b4955842e07c4d78300f110230370, /* 1582 */
128'hd52ff0efc43ec24a8526858a46010107, /* 1583 */
128'h00f41f634791c24a00f110234799ed19, /* 1584 */
128'h70e2d34ff0ef8526858a4601c43e4789, /* 1585 */
128'hfef414e3478580826121790274a27442, /* 1586 */
128'h87ae00f5f3634f5c6918ee09b7cdc402, /* 1587 */
128'hdd0c0007059b00e7f46385be27814f18, /* 1588 */
128'h0737691c80828082c2cff06f02c50823, /* 1589 */
128'hf0caf4a6fc86f8a2070d4b9c71191000, /* 1590 */
128'h8fd9f466f862fc5ee0dae4d6e8d2ecce, /* 1591 */
128'h6b9c679c681cc509f11ff0ef842ac17c, /* 1592 */
128'hf0efe22505130000551702042423eb8d, /* 1593 */
128'h74a679068526744670e6f8500493bacf, /* 1594 */
128'h61097ca27c427be26b066aa66a4669e6, /* 1595 */
128'h2c23478df93ff0eff3e54481541c8082, /* 1596 */
128'hf0ef852202042c2302f4082347851af4, /* 1597 */
128'h679c8522681c421010ef7d000513ba2f, /* 1598 */
128'h18042e2308842783f94584aa97826b9c, /* 1599 */
128'hf0ef8522d85c478508f422231a042823, /* 1600 */
128'hf0ef8522f1dff0ef852245814601b72f, /* 1601 */
128'h000505a345d000ef8522f14984aacf2f, /* 1602 */
128'h8ff94bdc00ff8737681c00f1102347a1, /* 1603 */
128'h858a460147d50aa00713e3991aa00713, /* 1604 */
128'h00c14703e911bf8ff0efc23ec43a8522, /* 1605 */
128'h0913cc1c800207b700f715630aa00793, /* 1606 */
128'h8bb74b0502900a934a55037009933e90, /* 1607 */
128'h8522858a460140000cb780020c3700ff, /* 1608 */
128'h681ce13dbb6ff0efc402c25201311023, /* 1609 */
128'hc43e0177f7b3c25a4bdc015110234c18, /* 1610 */
128'h8522858a4601c43e0197e7b301871563, /* 1611 */
128'h0863397d0007ca6347b2ed1db8eff0ef, /* 1612 */
128'h07374c14bf45331010ef3e8005130609, /* 1613 */
128'hd79bc43ccc188001073700e685638002, /* 1614 */
128'h18f40ca3478506041e23d45c8b8541e7, /* 1615 */
128'hc04ff0ef852202f51f63f9200793b55d, /* 1616 */
128'h0007d663443ced09c34ff0ef85224581, /* 1617 */
128'hc1cff0ef85224585bfd118f40c234785, /* 1618 */
128'h0493a10ff0efc9e5051300005517d965, /* 1619 */
128'hf706f3227161551cb58584aab595fa10, /* 1620 */
128'hf2e2f6defadafed6e352e74eeb4aef26, /* 1621 */
128'h10ef45018baae3b54401e6eeeaeaeee6, /* 1622 */
128'h180b8ca3198bc783c7b1199bc7831ff0, /* 1623 */
128'h855e008c479d460104f110234789e7b5, /* 1624 */
128'ha783120500e3842aabaff0efc482c2be, /* 1625 */
128'hf0ef855e008c46014495cf818b851b8b, /* 1626 */
128'h020ba423f4fd34fd100503e3842aaa0f, /* 1627 */
128'h70ba8522d55d842ad99ff0ef855ea031, /* 1628 */
128'h7bb67b567af66a1a69ba695a64fa741a, /* 1629 */
128'h048ba7838082615d6db66d566cf67c16, /* 1630 */
128'h4501b16ff0ef855e0407c163180b8c23, /* 1631 */
128'h45853e80091390810205149316d010ef, /* 1632 */
128'hcc63048ba783f155842ab36ff0ef855e, /* 1633 */
128'h0640051312a96ee3149010ef85260007, /* 1634 */
128'ha78300fbac23400007b7bfe91d7010ef, /* 1635 */
128'h9e23478502fba6238b8541e7d79b048b, /* 1636 */
128'h0ea61ee345111aa60f63450dbf0506fb, /* 1637 */
128'hac234006061b40010637a02940040637, /* 1638 */
128'h65898993000039978a9d0036d61b00cb, /* 1639 */
128'h1086a6830f86460396ce964e068a8a3d, /* 1640 */
128'h8a0500c7d61b02d606bb018ba8834505, /* 1641 */
128'h08dba42304cba823180bae231a0ba823, /* 1642 */
128'ha62300d5183b8abd0107d69b08dba223, /* 1643 */
128'h8e6302cba683090ba8231408dc63090b, /* 1644 */
128'h8ff50107571b003f06b70107979b1406, /* 1645 */
128'h00e797b3070907854721938117828fd9, /* 1646 */
128'h0c0bb4230c0bb0230a0bbc23030787b3, /* 1647 */
128'h0afbb8230e0bb0230c0bbc230c0bb823, /* 1648 */
128'h090ba70308fba6230107d46320000793, /* 1649 */
128'ha783c21508fba82300e7f46320000793, /* 1650 */
128'h46010107979b471100e78e63577d04cb, /* 1651 */
128'h902ff0efc282c4be04e11023855e008c, /* 1652 */
128'h979b4601495507cbd78304f11023479d, /* 1653 */
128'h842a8e4ff0efc4bec2ca855e008c0107, /* 1654 */
128'h08fb80a357fd08fbaa234785e40516e3, /* 1655 */
128'h00ef855ee2051ae3842ac9aff0ef855e, /* 1656 */
128'h1fe3842affbfe0ef855e00b545830f70, /* 1657 */
128'h2789100007b754075a63018ba703e005, /* 1658 */
128'h07cbd78306f110230370079304fba023, /* 1659 */
128'hf0efd4bed2ca855e0107979b108c4601, /* 1660 */
128'h033007930bf104934905d2caed05880f, /* 1661 */
128'h0a854a11d48206f11023988102091a93, /* 1662 */
128'hf0efd05aec56e826855e108c08104b21, /* 1663 */
128'h0637bb45842afe0a16e33a7dc131850f, /* 1664 */
128'h89bd0165d59bbd9940030637a7a94002, /* 1665 */
128'h979b16f16685b54d08bba82300b515bb, /* 1666 */
128'h00f7571b17828fd501e7569b8ff50027, /* 1667 */
128'h0187569b00ff05374098b5558b1d9381, /* 1668 */
128'h0087569b8e698fd50087161b0187179b, /* 1669 */
128'haa2327818fd58ef1f00706138fd16741, /* 1670 */
128'h159b8ecd0187169b0187559b40d804fb, /* 1671 */
128'hac238f558f718ecd0087571b8de90087, /* 1672 */
128'h02634689212700638b3d0187d71b04eb, /* 1673 */
128'h596302d7971300ebac238001073720d7, /* 1674 */
128'h04fba0238fd920000737040ba7830007, /* 1675 */
128'h000057971ef71863800107b7018ba703, /* 1676 */
128'ha783f0be4d05040ba903639c08478793, /* 1677 */
128'h79334724849300003497020d1a13044b, /* 1678 */
128'h0a05fe07fc1383f979130ff1079300f9, /* 1679 */
128'h8563278100f977b300e797bb47854098, /* 1680 */
128'h97d6109c840b0b1b4a81017d8b371607, /* 1681 */
128'h81630197f7b300f977b340dc0007ac83, /* 1682 */
128'h200007b700fc8d6345a1400007b71407, /* 1683 */
128'hb59340bc85b3100005b700fc88634591, /* 1684 */
128'h07370e051c638daa971ff0ef855e0015, /* 1685 */
128'h886347912000073700ec8d6347a14000, /* 1686 */
128'haa23001cb79340fc8cb3100007b700ec, /* 1687 */
128'h470d01a78663409cdfdfe0ef855e02fb, /* 1688 */
128'hd33e47d50af1102347994d850ce79163, /* 1689 */
128'h0110d53e00fde7b317c12d81810007b7, /* 1690 */
128'he0efc93ee552e162855e110c04000793, /* 1691 */
128'h409c09b794638bbd010c4783e941e91f, /* 1692 */
128'hb79317ed088ba58314079a631afba823, /* 1693 */
128'hf0ef855e460118fbae2308bba2230017, /* 1694 */
128'h102303700793fe07fd930ff10793947f, /* 1695 */
128'h110c0107979b4601475507cbd7830af1, /* 1696 */
128'he915e35fe0efd53ee03ad33a8cee855e, /* 1697 */
128'h07134791d502d33a0af1102347b56702, /* 1698 */
128'hc93ae552e16ee43e855e110c01100400, /* 1699 */
128'h37fd670267a20e050c63e0dfe0efe03a, /* 1700 */
128'h096ba2231afba823017d85b74785f3ed, /* 1701 */
128'h8c9ff0ef855e840585934601180bae23, /* 1702 */
128'h87930000379704a1eafa94e347a10a91, /* 1703 */
128'he0ef77a5051300004517e6f49fe32ee7, /* 1704 */
128'ha007071b80011737b61ddf400413cbdf, /* 1705 */
128'h5ee30307971300ebac2380020737b519, /* 1706 */
128'h0ab70ff104934905bbc580030737de07, /* 1707 */
128'h08633a7d09053ac54a15988119020100, /* 1708 */
128'h07931030c33e47d508f110234799020a, /* 1709 */
128'he0efdc3ef84af426c556855e010c0400, /* 1710 */
128'h44dcfbe18b8583a54cdcd0051ce3d61f, /* 1711 */
128'h8ff50087d79b0087961bf006869366c1, /* 1712 */
128'h6793da06d9e3040ba70302e796938fd1, /* 1713 */
128'heaf768e34581472db35d04fba0230087, /* 1714 */
128'h66c1b54511872583974e837902079713, /* 1715 */
128'h000da783f006869300ff0537040d8593, /* 1716 */
128'h0087961b8f510187971b0187d61b0d91, /* 1717 */
128'hfefdae238fd98ff58f510087d79b8e69, /* 1718 */
128'h8bbd00c7579b46a5008ca703fdb59ee3, /* 1719 */
128'h04d61c63800306b7018ba60300f6f863, /* 1720 */
128'h1487a78397b6078a1406869300003697, /* 1721 */
128'h17fd67c100cca68308fbae230087171b, /* 1722 */
128'h771327810126d71b8fd10186d61b8ff9, /* 1723 */
128'hd69b02e6073b3e800613c305c38d03f7, /* 1724 */
128'h0afba02302d606bb02f757bb8a8d0106, /* 1725 */
128'h19cba7831afbaa231b0ba7830adba223, /* 1726 */
128'h855e08fba82308fba62320000793c799, /* 1727 */
128'h08cba7030005062300051523484000ef, /* 1728 */
128'hccc68693aaa78793ccccd6b7aaaab7b7, /* 1729 */
128'h00f037b3068600d036b327818ef98ff9, /* 1730 */
128'h00d036b38ef90f068693f0f0f6b79fb5, /* 1731 */
128'h36b38ef9f0068693ff0106b79fb5068a, /* 1732 */
128'h37338f750207161376c19fb5068e00d0, /* 1733 */
128'hed1092010a8bb783d11c9fb9071200e0, /* 1734 */
128'h06fbc603074bd68307abd70302c7d7b3, /* 1735 */
128'h3623024505135b6585930000459784aa, /* 1736 */
128'hc603077bc883070ba803a95fe0effef5, /* 1737 */
128'hf7930188569b0108571b0088579b06cb, /* 1738 */
128'h0000459726810ff777130ff878130ff7, /* 1739 */
128'h074ba603a5ffe0ef04d4851359458593, /* 1740 */
128'h0106569b062485135905859300004597, /* 1741 */
128'h10ef8526a3ffe0ef8a3d8abd0146561b, /* 1742 */
128'h2785100007b7b8d102fba42347857e40, /* 1743 */
128'hecf76ce31a0bb683400407b704fba023, /* 1744 */
128'h70000737bb9550e5051300004517e691, /* 1745 */
128'h03f7f6930c46c78304fba0230017079b, /* 1746 */
128'hc68900c7f693ce910027f6931adba423, /* 1747 */
128'h01076713040ba70304eba0230217071b, /* 1748 */
128'h00c7e793040ba783c7998b8504eba023, /* 1749 */
128'h088ba583044ba783040baa0304fba023, /* 1750 */
128'hff0484930000349700fa7a33855e4601, /* 1751 */
128'h4c2d002b0b1300003b174a85db4ff0ef, /* 1752 */
128'h77b300fa97bb409c034c8c9300003c97, /* 1753 */
128'h0d37fe29091300003917cbb5278100fa, /* 1754 */
128'hb79317ed00494703409c10000db72000, /* 1755 */
128'h00fa77b30009270340dc04f718630017, /* 1756 */
128'hf69345850b70061300894683c3a18ff9, /* 1757 */
128'h0b7006134681c131debfe0ef855e0fb6, /* 1758 */
128'h1a0ba823088ba783ddbfe0ef855e4585, /* 1759 */
128'he0ef855e035baa2308fba223180bae23, /* 1760 */
128'h4517f7649fe304a1fb9911e30931973f, /* 1761 */
128'h00092783bb6d925fe0ef3e2505130000, /* 1762 */
128'h01a78663471100d789634721400006b7, /* 1763 */
128'he0ef855e02ebaa230017b71341b787b3, /* 1764 */
128'h00892683f941808ff0ef855e408c933f, /* 1765 */
128'ha583ef8d1afba823409ce79d0046f793, /* 1766 */
128'h18fbae2308bba2230017b79317ed088b, /* 1767 */
128'hfd319fdfe0ef855ecb0ff0ef855e4601, /* 1768 */
128'he0ef855e45850b7006130ff6f693bb91, /* 1769 */
128'h02079713fcfc65e34581b7c9f521d31f, /* 1770 */
128'h851300ec4641bf6d11872583974e8379, /* 1771 */
128'h07cbd78304f11023478d6da000ef06cb, /* 1772 */
128'hc2be47d5855ec4be0107979b008c4601, /* 1773 */
128'hd663018ba783ec051b63842a96ffe0ef, /* 1774 */
128'h04f1102347a506fb9e2304e157830007, /* 1775 */
128'h0107979b008c460107cbd783c2be479d, /* 1776 */
128'h46b6ea051163842a93bfe0efc4be855e, /* 1777 */
128'ha02304dbae23018ba50345e6475647c6, /* 1778 */
128'h1a634000063706bba42306eba22306fb, /* 1779 */
128'h43638ca602e345098a3d01a6d61bf2c5, /* 1780 */
128'h2006061b40010637f0a609634505f0c5, /* 1781 */
128'h4501c56ce54ff06ffa100413f0eff06f, /* 1782 */
128'h808218b50d238082557d8082557d8082, /* 1783 */
128'h47851141ef9d439cc347879300005797, /* 1784 */
128'h00efc0f72f2300005717842ae406e022, /* 1785 */
128'hf0ef852200055563aeefe0ef852212a0, /* 1786 */
128'h60a20dc000ef13e000ef02c00513fc5f, /* 1787 */
128'h00005717808245018082014145016402, /* 1788 */
128'h85aa114102e790636394631cbec70713, /* 1789 */
128'h60a2f60fe0efe4063905051300004517, /* 1790 */
128'h00a604630fc7a60380820141853e4781, /* 1791 */
128'he42eec06110141488082853ebfd187b6, /* 1792 */
128'h02b7006365a210354703c105fbdff0ef, /* 1793 */
128'h610560e200f70c630ff0079308154703, /* 1794 */
128'hbfe545018082610560e25535eb3fe06f, /* 1795 */
128'h84aee822ec06e4261101bfcdf8400513, /* 1796 */
128'h0413e501cf0ff0ef842acd09f7dff0ef, /* 1797 */
128'h55358082610564a2644260e2e0800f84, /* 1798 */
128'h0015071b43889d67879300005797bfd5, /* 1799 */
128'h87930000579780820f8505138082c398, /* 1800 */
128'hb2078793000057971101808243889be7, /* 1801 */
128'h60e20094176384beec06e4266380e822, /* 1802 */
128'h8522c78119a447838082610564a26442, /* 1803 */
128'haf07879300005797b7d56000a9cff0ef, /* 1804 */
128'he50880829607aa2300005797e79ce39c, /* 1805 */
128'he518e11ce7886798ad87879300005797, /* 1806 */
128'hac04849300005497e4a6711d8082e308, /* 1807 */
128'he862ec5ef05af456f852fc4e6080e8a2, /* 1808 */
128'h0a1300004a1789aae0caec86e06ae466, /* 1809 */
128'h0b1300004b1726ea8a9300004a9727ea, /* 1810 */
128'h4c9700050c1b276b8b9300004b97276b, /* 1811 */
128'h60e66446029415634d2985ac8c930000, /* 1812 */
128'h6c426be27b027aa27a4279e2690664a6, /* 1813 */
128'he06f61253c450513000045176d026ca2, /* 1814 */
128'h0007c36389524c1cc7914901541cddcf, /* 1815 */
128'hdbefe0ef638c855a0fc42603681c8956, /* 1816 */
128'h8e63601cdb2fe0ef855e85ca00090663, /* 1817 */
128'h351701a98863da4fe0ef856685e20097, /* 1818 */
128'h1101b771600032a010ef7e2505130000, /* 1819 */
128'h44014d1cc1414401e04ae426ec06e822, /* 1820 */
128'h639cc7bd651ccbad511ccbbd4d5ccfad, /* 1821 */
128'h200010ef45051c00059384aa892ec7ad, /* 1822 */
128'h47850ef52c234799c57c57fdcd21842a, /* 1823 */
128'hf0ef0405282303253023e90410f502a3, /* 1824 */
128'h179716f43c2391c78793fffff797e65f, /* 1825 */
128'h87930000179718f430232be787930000, /* 1826 */
128'hc78385220ea42e23681c18f434232ae7, /* 1827 */
128'h644260e28522e99ff0ef10f400230247, /* 1828 */
128'h000046971bc0106f80826105690264a2, /* 1829 */
128'h671302d786b365186294611c6fc68693, /* 1830 */
128'h93ed836d8f3d0127d713e11897360017, /* 1831 */
128'h25018d5d00f717bb40f007b300f7553b, /* 1832 */
128'h1141fc3ff06f93650513000055178082, /* 1833 */
128'h151bfe9ff0ef842afefff0efe022e406, /* 1834 */
128'h1141808201412501640260a28d410105, /* 1835 */
128'hf0ef14020005041bfdbff0efe022e406, /* 1836 */
128'h80820141640260a28d4115029001fd1f, /* 1837 */
128'hfb75fee78fa30785fff5c703058587aa, /* 1838 */
128'hfff5c703058500c7896387aa962a8082, /* 1839 */
128'h0007c70387aa8082fb65fee78fa30785, /* 1840 */
128'h8fa30785fff5c7030585eb0900178693, /* 1841 */
128'h8082e21987aab7d587b68082fb75fee7, /* 1842 */
128'h0585963efb7d001786930007c70387b6, /* 1843 */
128'h8082e291fed70fa300178713fff5c683, /* 1844 */
128'h0585b7cd87ba8082000780a300c71563, /* 1845 */
128'h0187979b40f707bbfff5c78300054703, /* 1846 */
128'h962e8082853ef37d0505e3994187d79b, /* 1847 */
128'hc783000547030585a839478100c59463, /* 1848 */
128'he3994187d79b0187979b40f707bbfff5, /* 1849 */
128'h000547830ff5f5938082853eff790505, /* 1850 */
128'h80824501bfcd0505c399808200b79363, /* 1851 */
128'hdffd808200b79363000547830ff5f593, /* 1852 */
128'h40a78533e7010007c70387aabfcd0505, /* 1853 */
128'hec06842ae42ee8221101bfcd07858082, /* 1854 */
128'h000547830ff5f593952265a2fe5ff0ef, /* 1855 */
128'h644260e24501fe857be3157d00b78663, /* 1856 */
128'h0007c70300b7856387aa95aa80826105, /* 1857 */
128'h87aa862ab7fd0785808240a78533e701, /* 1858 */
128'hfed80fe38082ea9940c785330007c683, /* 1859 */
128'h872eb7d50785fe081be3000748030705, /* 1860 */
128'hea1140d785330007c60387aa86aabfcd, /* 1861 */
128'hfe081be300074803070500c80a638082, /* 1862 */
128'heb1900054703bff90785bfd5872e8082, /* 1863 */
128'hfafd0007c6830785fee68fe380824501, /* 1864 */
128'hec06e426e8221101bfd587aeb7e50505, /* 1865 */
128'h63807327879300004797e519842a84ae, /* 1866 */
128'h00044783942af9dff0ef85a68522cc11, /* 1867 */
128'h60e2852244017007bb2300004797ef81, /* 1868 */
128'hf9fff0ef852285a68082610564a26442, /* 1869 */
128'h4797050500050023c78100054783c519, /* 1870 */
128'hec066104e4261101bfd96ea7b5230000, /* 1871 */
128'h0023c501f73ff0ef8526842ac891e822, /* 1872 */
128'h610564a28526644260e2e00805050005, /* 1873 */
128'h0007c68387aacf9900054783c11d8082, /* 1874 */
128'h80a300e780238082e3110017c703ce81, /* 1875 */
128'hcb9d0075779380824501b7e5078900d7, /* 1876 */
128'h377d8fd507a2808204c79063963e87aa, /* 1877 */
128'hef6340e88833469d00c508b3872aff6d, /* 1878 */
128'h97aa078e02e787335761003657930106, /* 1879 */
128'h3c230721bfd10ff5f6934725bfc1963a, /* 1880 */
128'h00b50a63bf6dfeb78fa30785bfe1fef7, /* 1881 */
128'h02c79e63963e87aacb9d8b9d00a5e7b3, /* 1882 */
128'h8833ff07bc2307a1ff87380307218082, /* 1883 */
128'h02f707b357e100365713ff06e8e340f8, /* 1884 */
128'h87aa872ebfc100e507b3963e95ba070e, /* 1885 */
128'h0785fff5c7030585bfe1469d00c508b3, /* 1886 */
128'hec26852e842af0227179bf65fee78fa3, /* 1887 */
128'h84aa6622dcdff0efe02ee84af406e432, /* 1888 */
128'h8522fff6091300c564636582892ace11, /* 1889 */
128'h740270a200040023f79ff0ef944a864a, /* 1890 */
128'he406e02211418082614564e269428526, /* 1891 */
128'h640260a28522f57ff0ef00a5e963842a, /* 1892 */
128'h87b340b6073300c506b395b280820141, /* 1893 */
128'h00f6802316fd0005c78315fdd7e500e5, /* 1894 */
128'h47838082853e478100c51563962ab7fd, /* 1895 */
128'hb7dd05850505fbed9f990005c7030005, /* 1896 */
128'hfeb78de300054783808200c51363962a, /* 1897 */
128'he44eec26852e842af0227179bfc50505, /* 1898 */
128'hc8890005049bd1fff0ef89aee84af406, /* 1899 */
128'h440100995b630005091bd13ff0ef8522, /* 1900 */
128'h8082614569a2694264e2740270a28522, /* 1901 */
128'h0405d175f8bff0ef397d852285ce8626, /* 1902 */
128'h8082450100c514630ff5f593962abfe9, /* 1903 */
128'hb7ed853efeb70be30015079300054703, /* 1904 */
128'he60187aa260100c7ef630ff5f59347c1, /* 1905 */
128'h0785feb71ce30007c7038082853e4781, /* 1906 */
128'h40e7873b47a1c31d00757713b7f5367d, /* 1907 */
128'h36fdfcb81ce30007c80387aa0007069b, /* 1908 */
128'h97938e1d953e938102071793faf50785, /* 1909 */
128'h020796938fd90107179300b7e7330085, /* 1910 */
128'hd24d8a1deb1187aa27018edd00365713, /* 1911 */
128'hb803bfcd367d0785f8b71fe30007c703, /* 1912 */
128'h12e30007c70300d80a63008785130007, /* 1913 */
128'hb7f1377d87aabfa5fef51be30785f8b7, /* 1914 */
128'h08f711630300079300054703e7a9419c, /* 1915 */
128'h00e786b313c787930000279700154703, /* 1916 */
128'h0ff777130207071bc6898a850006c683, /* 1917 */
128'hc78397ba0025470304d71b6307800693, /* 1918 */
128'h47c14198c19c47c1c3b10447f7930007, /* 1919 */
128'h02f71663030007930005470302f71c63, /* 1920 */
128'h4703973e0ec707130000271700154783, /* 1921 */
128'h07130ff7f7930207879bc7098b050007, /* 1922 */
128'h47a9bf7d47a18082050900e793630780, /* 1923 */
128'hf0efc632ec06006c842ee8221101bf6d, /* 1924 */
128'h0a88081300002817468100c16583f63f, /* 1925 */
128'h0006460300f806330007079b00054703, /* 1926 */
128'h8536644260e2ec050008986304467893, /* 1927 */
128'hfd07879b00088b630046789380826105, /* 1928 */
128'h8a09b7d196be050502d586b3feb7f4e3, /* 1929 */
128'hb7cdfc97879b0ff7f793fe07079bc609, /* 1930 */
128'h3023f04afc06f426f8227139b7e1e008, /* 1931 */
128'he90165a2b0dff0ef84b2842ae42e0006, /* 1932 */
128'h862e80826121790274a2744270e25529, /* 1933 */
128'hfe8782e367e2f5dff0ef8522082c892a, /* 1934 */
128'h47a9fd279be307858f81cb010007c703, /* 1935 */
128'h071300054683b7e94501e088fcf718e3, /* 1936 */
128'he40605051141f2dff06f00e6846302d0, /* 1937 */
128'h11418082014140a0053360a2f23ff0ef, /* 1938 */
128'h04b00693601cf0dff0ef842ee406e022, /* 1939 */
128'h0470069300e6ea6302d704630007c703, /* 1940 */
128'h04d0069380820141640260a202d70e63, /* 1941 */
128'h0017c683fed716e306b0069302d70763, /* 1942 */
128'h07130027c683fce69fe3052a06900713, /* 1943 */
128'h052a052ab7e9e01c078d00e698630420, /* 1944 */
128'hec06006c842ee8221101bfd50789bff1, /* 1945 */
128'h00002817468100c16583e0fff0efc632, /* 1946 */
128'h00f806330007079b00054703f5480813, /* 1947 */
128'h60e2ec05000898630446789300064603, /* 1948 */
128'h00088b63004678938082610585366442, /* 1949 */
128'h96be050502d586b3feb7f4e3fd07879b, /* 1950 */
128'h879b0ff7f793fe07079bc6098a09b7d1, /* 1951 */
128'h842ee406e0221141b7e1e008b7cdfc97, /* 1952 */
128'h04630007c70304b00693601cf87ff0ef, /* 1953 */
128'h60a202d70e630470069300e6ea6302d7, /* 1954 */
128'h069302d7076304d00693808201416402, /* 1955 */
128'h052a069007130017c683fed716e306b0, /* 1956 */
128'h00e69863042007130027c683fce69fe3, /* 1957 */
128'hbfd50789bff1052a052ab7e9e01c078d, /* 1958 */
128'h05b395bff0efe589842ae406e0221141, /* 1959 */
128'h8513e7a7879300002797fff5c70300a4, /* 1960 */
128'h640260a2e7198b1100074703973efff5, /* 1961 */
128'h00054703fea47ae3157d80820141557d, /* 1962 */
128'h462960a26402f77d8b1100074703973e, /* 1963 */
128'hfa5ff06f4581d7dff06f014105054581, /* 1964 */
128'h00e1550300a10723812100a107a31141, /* 1965 */
128'h1582639c30c787930000479780820141, /* 1966 */
128'h46254781aa5ff06f95be920116029181, /* 1967 */
128'hfd07069b8082853ee3190005470345a9, /* 1968 */
128'h879b9fb902f587bb00d667630ff6f693, /* 1969 */
128'h4563842ee406e0221141bff90505fd07, /* 1970 */
128'h357d02b455bb45a900b7f86347a500a0, /* 1971 */
128'h014160a2640202a4753b4529fe7ff0ef, /* 1972 */
128'h471707e2081007935000006f03050513, /* 1973 */
128'h808228f739230000471728f739230000, /* 1974 */
128'h862ee4262844041300004417e8221101, /* 1975 */
128'h60e2600ca15ff0efec06600885aa84ae, /* 1976 */
128'h479711018082610564a26442e00c95a6, /* 1977 */
128'h2484849300004497e42625a787930000, /* 1978 */
128'hec0680250513000045176380e8226090, /* 1979 */
128'he63fc0ef85a26088b87fd0ef85a29c11, /* 1980 */
128'hd0ef7fa5051300003517862286aa608c, /* 1981 */
128'h0517b61fd0ef8065051300004517b6df, /* 1982 */
128'h644200055e638a1f90efef6505130000, /* 1983 */
128'h7f8505130000351740a005b364a260e2, /* 1984 */
128'h006f610564a260e26442b39fd06f6105, /* 1985 */
128'h03638c2fa0ef8432e406e02211416680, /* 1986 */
128'h8082450180820141640260a2557d0085, /* 1987 */
128'hf606852289aae64e01258413f2227169, /* 1988 */
128'h00a404b30505f7eff0ef892eea4aee26, /* 1989 */
128'h071be93ff0ef95260505f72ff0ef8526, /* 1990 */
128'ha7230000479704e7ee631ff00793fff5, /* 1991 */
128'h05130000351784aaf50ff0ef852216a7, /* 1992 */
128'h04a7f2630ff007939526f42ff0ef56e5, /* 1993 */
128'h5505051300003517842af32ff0ef8522, /* 1994 */
128'h768505130000351700a405b3f24ff0ef, /* 1995 */
128'h615569b2695264f2741270b2a8bfd0ef, /* 1996 */
128'hb75510f7292300004717200007938082, /* 1997 */
128'h00003597863ff0ef850a458110000613, /* 1998 */
128'h079301294703deaff0ef850a50c58593, /* 1999 */
128'h850a73a585930000359700f7096302f0, /* 2000 */
128'h00004797df2ff0ef850a85a2dfaff0ef, /* 2001 */
128'h7205051300003517858a43900cc78793, /* 2002 */
128'h00004717451107e208100793a1bfd0ef, /* 2003 */
128'hd85ff0ef0af73a23000047170af73a23, /* 2004 */
128'h4797d77ff0ef4501e8a7982300004797, /* 2005 */
128'he7858593000045974611e8a792230000, /* 2006 */
128'h06f71a23000047174785eb1ff0ef854e, /* 2007 */
128'h8432478de04ae426ec06e8221101b791, /* 2008 */
128'hd783d37ff0ef84ae450d892a08c7df63, /* 2009 */
128'h044555030000451708a7956325010004, /* 2010 */
128'h059b06a79a6325010024d783d21ff0ef, /* 2011 */
128'hd05ff0ef4511dabff0ef00448513ffc4, /* 2012 */
128'h0145550300004517e0a7982300004797, /* 2013 */
128'h4597dea79e23000047974611cf1ff0ef, /* 2014 */
128'h00ef4535e2bff0ef854adf2585930000, /* 2015 */
128'hd1bff0ef4515fea5d583000045972560, /* 2016 */
128'hfd47879300004797240000ef02000513, /* 2017 */
128'h4797fcf713230000471727850007d783, /* 2018 */
128'h35170087cf63278d439cfba787930000, /* 2019 */
128'h64a260e26442905fd0ef62a505130000, /* 2020 */
128'h690264a2644260e2d49ff06f61056902, /* 2021 */
128'h47090105c783f022f406717980826105, /* 2022 */
128'h01e1578300f10f230115c78300f10fa3, /* 2023 */
128'h351770a2740202e78a63470d00e78e63, /* 2024 */
128'h3517842a8b3fd06f614560a505130000, /* 2025 */
128'h740285228a3fd0efe42e5e2505130000, /* 2026 */
128'h70a241907402d8bff06f614570a265a2, /* 2027 */
128'h22813823dc010113ebfff06f614505c1, /* 2028 */
128'h4581893284ae842a2321302322913423, /* 2029 */
128'h85a6e60ff0ef22113c23002821800613, /* 2030 */
128'h002cea2ff0efe802c44a082820400613, /* 2031 */
128'h34832301340323813083f63ff0ef8522, /* 2032 */
128'h00004797808224010113220139032281, /* 2033 */
128'hcb858593000045974611cb81ed07d783, /* 2034 */
128'he703504000efe40611418082cf3ff06f, /* 2035 */
128'ha02327051001a70300e57763878e1041, /* 2036 */
128'h1782150260a21007e78310a7a22310e1, /* 2037 */
128'hec06110180824501808201418d5d9101, /* 2038 */
128'h440000ef842afc1ff0ef84aae426e822, /* 2039 */
128'h644260e29101150202f407b33e800793, /* 2040 */
128'he40611418082610564a28d0502a7d533, /* 2041 */
128'h000f47b7414000ef842af95ff0efe022, /* 2042 */
128'h91011502640260a202f407b324078793, /* 2043 */
128'he426e822ec061101808202a7d5330141, /* 2044 */
128'h85333e2000ef892af63ff0ef84aae04a, /* 2045 */
128'h944a0285543324040413000f443702a4, /* 2046 */
128'h64a2644260e2fe856ee3f45ff0ef0405, /* 2047 */
128'he822009894b7e4261101808261056902, /* 2048 */
128'h0084f363892268048493842ae04aec06, /* 2049 */
128'h60e2f47dfa1ff0ef41240433854a8926, /* 2050 */
128'h808200b5002380826105690264a26442, /* 2051 */
128'h75130147c503100007b7808200054503, /* 2052 */
128'h0207f793014747831000073780820205, /* 2053 */
128'h00078223100007b7808200a70023dfe5, /* 2054 */
128'h822300e78023476d00e78623f8000713, /* 2055 */
128'h00e78423fc70071300e78623470d0007, /* 2056 */
128'he406e0221141808200e7882302000713, /* 2057 */
128'h80820141640260a2e50900044503842a, /* 2058 */
128'hda07879300002797b7f50405fa5ff0ef, /* 2059 */
128'hc7830007470397aa973e811100f57713, /* 2060 */
128'he8221101808200f5802300e580a30007, /* 2061 */
128'h00814503fd1ff0efec068121842a002c, /* 2062 */
128'h7513002cf5dff0ef00914503f65ff0ef, /* 2063 */
128'h4503f4bff0ef00814503fb7ff0ef0ff4, /* 2064 */
128'h717980826105644260e2f43ff0ef0091, /* 2065 */
128'h553b54e14461892af406e84aec26f022, /* 2066 */
128'h00814503f81ff0ef0ff57513002c0089, /* 2067 */
128'h10e3f0bff0ef00914503f13ff0ef3461, /* 2068 */
128'h717980826145694264e2740270a2fe94, /* 2069 */
128'h54e103800413892af406e84aec26f022, /* 2070 */
128'h4503f3fff0ef0ff57513002c00895533, /* 2071 */
128'hec9ff0ef00914503ed1ff0ef34610081, /* 2072 */
128'h80826145694264e2740270a2fe9410e3, /* 2073 */
128'hf0ef00814503f13ff0efec06002c1101, /* 2074 */
128'h8082610560e2e9fff0ef00914503ea7f, /* 2075 */
128'hf426f8227139439ce787879300004797, /* 2076 */
128'h02b7856384b2842e892aec4efc06f04a, /* 2077 */
128'hc10d2501f3afb0efc205051300004517, /* 2078 */
128'h790274a2744270e2e4a7a62300004797, /* 2079 */
128'he2f728230000471757fd8082612169e2, /* 2080 */
128'hb0efbea505130000451785ca86260074, /* 2081 */
128'h4632e0a7ab2300004797c50d2501814f, /* 2082 */
128'hd0ef282505130000351785a604967563, /* 2083 */
128'h4521b775def72c23000047174785d0cf, /* 2084 */
128'h000037970009099b00c4591be05ff0ef, /* 2085 */
128'hf0ef00094503993e0039791327c78793, /* 2086 */
128'h000047979c25bf5d320010ef854ede7f, /* 2087 */
128'h3517842a85aae0221141bf95da87ae23, /* 2088 */
128'h0000100fcb2fd0efe406252505130000, /* 2089 */
128'h259760a264028322f14025730ff0000f, /* 2090 */
128'h35974605114183020141c02585930000, /* 2091 */
128'he406d7a5051300004517f3a585930000, /* 2092 */
128'h051300003517c9112501d79fa0efe022, /* 2093 */
128'h00003517c62fd06f014160a264022365, /* 2094 */
128'h8593000035974605c56fd0ef24450513, /* 2095 */
128'h2501d9bfa0efafe50513000045172565, /* 2096 */
128'h00003517b7e124e5051300003517c511, /* 2097 */
128'he985051300000517c26fd0ef0cc50513, /* 2098 */
128'hd007a02300004797d007a62300004797, /* 2099 */
128'h87930000479700054863842a956f90ef, /* 2100 */
128'h351760a26402408005b3cf81439ccf27, /* 2101 */
128'h00004517be2fd06f01410a2505130000, /* 2102 */
128'h00003517c5112501b9afb0efa9450513, /* 2103 */
128'he7058593000035974605bfb91fc50513, /* 2104 */
128'h051300003517c5112501cb9fa0ef4501, /* 2105 */
128'h900200000023ee1ff0ef8522b7811f65, /* 2106 */
128'h000f4537a001d69ff0efe40625011141, /* 2107 */
128'h07130000471780824501808224050513, /* 2108 */
128'h95360017869300756513157d631cc667, /* 2109 */
128'h02b506338082953e055e10d00513e308, /* 2110 */
128'h842afd1ff0efe4328532ec06e8221101, /* 2111 */
128'h644260e28522944ff0ef45816622c509, /* 2112 */
128'h19050513000035171141808280826105, /* 2113 */
128'h60a2ee5fc0ef20000537b28fd0efe406, /* 2114 */
128'h25738082450180824501808201414501, /* 2115 */
128'h86b287361141808202f5553347a9b000, /* 2116 */
128'hd0efe40617c505130000351785aa862e, /* 2117 */
128'h842ae0221141a001cbbff0ef4505aecf, /* 2118 */
128'h60a29522408007b3f57ff0efe406952e, /* 2119 */
128'h8082450580824505808201418d7d6402, /* 2120 */
128'h84bb842ef406ec26f022717980824505, /* 2121 */
128'h6145450164e2740270a20096186300c6, /* 2122 */
128'h04136622e37fc0efe432852285b28082, /* 2123 */
128'h45098082450980824509bff926052004, /* 2124 */
128'h80824501808245018082808280828082, /* 2125 */
128'h96934781e426e822ec061101bbbff06f, /* 2126 */
128'h60e200c7986300d5043300d584b30037, /* 2127 */
128'h60980004380380826105450164a26442, /* 2128 */
128'h0f050513000035176090600c02e80363, /* 2129 */
128'h108505130000351785a28626a2afd0ef, /* 2130 */
128'h892ae0ca711dbf5d0785a001a1afd0ef, /* 2131 */
128'hf456f852fc4ee8a21085051300003517, /* 2132 */
128'h44018b2ee466e4a6ec86e862ec5ef05a, /* 2133 */
128'h00003b970f4a0a1300003a179eafd0ef, /* 2134 */
128'h100c0c1300003c17fff949930fcb8b93, /* 2135 */
128'h855e85e600040c9b9c6fd0ef85524ac1, /* 2136 */
128'hd0ef855203649863448187ca9bafd0ef, /* 2137 */
128'h9b63458187ca9a4fd0ef856285e69acf, /* 2138 */
128'h1285051300003517fd5417e3040502b4, /* 2139 */
128'h873e8a85008486b3a889450198afd0ef, /* 2140 */
128'h04856398e39840e9873300349713c689, /* 2141 */
128'hc689873e8a856390008586b3bf5d07a1, /* 2142 */
128'h3517058e02e60d6340e9873300359713, /* 2143 */
128'h051300003517944fd0ef08a505130000, /* 2144 */
128'h690664a6644660e6557d938fd0ef0b65, /* 2145 */
128'h61256ca26c426be27b027aa27a4279e2, /* 2146 */
128'h6a05fc56e0d27159bfa507a105858082, /* 2147 */
128'hf062f45ef85ae4ceeca6020005138aaa, /* 2148 */
128'h8bb28b2ee46ee86aec66e8caf0a2f486, /* 2149 */
128'h00003c179c4a0a134981b3fff0ef4481, /* 2150 */
128'h00fb0cb300fa8db3003497933ecc0c13, /* 2151 */
128'h8befd0ef084505130000351703749b63, /* 2152 */
128'h6ce27c027ba26a0669a6694670a67406, /* 2153 */
128'h7ae285567b4264e685da86266da26d42, /* 2154 */
128'hbd7fe0ef842abddfe0efe33ff06f6165, /* 2155 */
128'h0344f7b3bcbfe0ef892abd1fe0ef8d2a, /* 2156 */
128'h01a4643300a96533010d1d1b0105151b, /* 2157 */
128'h00adb02300acb0238d41910114021502, /* 2158 */
128'h97e20039f7930985aadff0ef4521ef81, /* 2159 */
128'he42e7139b7ad0485a9dff0ef0007c503, /* 2160 */
128'he0ef89aaec4ef04af426f822fc06e032, /* 2161 */
128'h84aab69fe0ef892ab6ffe0ef842ab75f, /* 2162 */
128'h8fc18d450109179b0105151bb63fe0ef, /* 2163 */
128'h971347818d5d9101178265a266021502, /* 2164 */
128'h70e2744200c79c63974e00e588330037, /* 2165 */
128'hd79ff06f6121863e69e2854e790274a2, /* 2166 */
128'h30238f2900083703e3148ea907856314, /* 2167 */
128'hf426f822fc06e032e42e7139b7f100e8, /* 2168 */
128'haf7fe0ef842aafdfe0ef89aaec4ef04a, /* 2169 */
128'h0105151baebfe0ef84aaaf1fe0ef892a, /* 2170 */
128'h178265a2660215028fc18d450109179b, /* 2171 */
128'h974e00e588330037971347818d5d9101, /* 2172 */
128'h69e2854e790274a270e2744200c79c63, /* 2173 */
128'he3148e8907856314d01ff06f6121863e, /* 2174 */
128'he42e7139b7f100e830238f0900083703, /* 2175 */
128'he0ef89aaec4ef04af426f822fc06e032, /* 2176 */
128'h84aaa79fe0ef892aa7ffe0ef842aa85f, /* 2177 */
128'h8fc18d450109179b0105151ba73fe0ef, /* 2178 */
128'h971347818d5d9101178265a266021502, /* 2179 */
128'h70e2744200c79c63974e00e588330037, /* 2180 */
128'hc89ff06f6121863e69e2854e790274a2, /* 2181 */
128'h073300083703e31402a686b307856314, /* 2182 */
128'hfc06e032e42e7139b7e100e8302302a7, /* 2183 */
128'h842aa09fe0ef89aaec4ef04af426f822, /* 2184 */
128'h9f7fe0ef84aa9fdfe0ef892aa03fe0ef, /* 2185 */
128'h660215028fc18d450109179b0105151b, /* 2186 */
128'h88330037971347818d5d9101178265a2, /* 2187 */
128'h790274a270e2744200c79c63974e00e5, /* 2188 */
128'h4505e111c0dff06f6121863e69e2854e, /* 2189 */
128'h573300083703e31402a6d6b307856314, /* 2190 */
128'hfc06e032e42e7139b7d100e8302302a7, /* 2191 */
128'h842a989fe0ef89aaec4ef04af426f822, /* 2192 */
128'h977fe0ef84aa97dfe0ef892a983fe0ef, /* 2193 */
128'h660215028fc18d450109179b0105151b, /* 2194 */
128'h88330037971347818d5d9101178265a2, /* 2195 */
128'h790274a270e2744200c79c63974e00e5, /* 2196 */
128'h07856314b8dff06f6121863e69e2854e, /* 2197 */
128'hb7f100e830238f4900083703e3148ec9, /* 2198 */
128'hec4ef04af426f822fc06e032e42e7139, /* 2199 */
128'he0ef892a90bfe0ef842a911fe0ef89aa, /* 2200 */
128'h0109179b0105151b8fffe0ef84aa905f, /* 2201 */
128'h8d5d9101178265a2660215028fc18d45, /* 2202 */
128'h00c79c63974e00e58833003797134781, /* 2203 */
128'h6121863e69e2854e790274a270e27442, /* 2204 */
128'h00083703e3148ee907856314b15ff06f, /* 2205 */
128'hfc06e032e42e7139b7f100e830238f69, /* 2206 */
128'h842a899fe0ef89aaec4ef04af426f822, /* 2207 */
128'h887fe0ef84aa88dfe0ef892a893fe0ef, /* 2208 */
128'h660214828fc18cc90109179b0105151b, /* 2209 */
128'h88330037169347018fc59081178265a2, /* 2210 */
128'h790274a270e2744200c71c6396ae00d9, /* 2211 */
128'h00f70533a9dff06f6121863a69e2854e, /* 2212 */
128'h892ae8ca7159bfc9070500a83023e288, /* 2213 */
128'hfc56e0d2e4cef0a2be85051300003517, /* 2214 */
128'h8b3289aeec66eca6f486f062f45ef85a, /* 2215 */
128'h3b97bd2a0a1300003a17cc9fc0ef4401, /* 2216 */
128'h0a93be2c0c1300003c17bdab8b930000, /* 2217 */
128'h855e85a2fff44493ca7fc0ef85520400, /* 2218 */
128'h179314fd460140900cb3c99fc0ef8885, /* 2219 */
128'he43285520566186397ce00f905b30036, /* 2220 */
128'h85ce6622c73fc0ef856285a2c7bfc0ef, /* 2221 */
128'hfb541be32405e12984aaa03ff0ef854a, /* 2222 */
128'h740670a6c53fc0efbf05051300003517, /* 2223 */
128'h7ba27b427ae26a0669a664e669468526, /* 2224 */
128'hc291876600167693808261656ce27c02, /* 2225 */
128'h7159bfc154fdbf590605e198e3988726, /* 2226 */
128'he8caf0a2b14505130000351784aaeca6, /* 2227 */
128'hf486ec66f062f45ef85afc56e0d2e4ce, /* 2228 */
128'h00003997bf3fc0ef44018ab2892ee86a, /* 2229 */
128'h00003b97dfcb0b1300003b17afc98993, /* 2230 */
128'h00003c97af4c0c1300003c17dfcb8b93, /* 2231 */
128'h7793bc1fc0ef854e04000a13afcc8c93, /* 2232 */
128'hbaffc0ef856285a2000bbd03cba50014, /* 2233 */
128'h97ca00f485b300361793fffd45134601, /* 2234 */
128'h856685a2b93fc0efe432854e05561c63, /* 2235 */
128'h8d2a91bff0ef852685ca6622b8bfc0ef, /* 2236 */
128'hb085051300003517fb441ae32405e529, /* 2237 */
128'h69a6694664e6856a740670a6b6bfc0ef, /* 2238 */
128'h61656d426ce27c027ba27b427ae26a06, /* 2239 */
128'hc291876a00167693bf49000b3d038082, /* 2240 */
128'h711db7e15d7db7790605e198e398872a, /* 2241 */
128'he0cae4a6a245051300003517842ae8a2, /* 2242 */
128'h84aefc4eec86e862ec5ef05af456f852, /* 2243 */
128'ha109091300003917b07fc0ef4c018ab2, /* 2244 */
128'ha20b8b9300003b97a18b0b1300003b17, /* 2245 */
128'h85ce000c099bae5fc0ef854a10000a13, /* 2246 */
128'h8fd9010c1793008c1713ad9fc0ef855a, /* 2247 */
128'h8fd9020c17138fd9018c17130187e7b3, /* 2248 */
128'h038c17138fd9030c17138fd9028c1713, /* 2249 */
128'h1763972600e406b30036171346018fd9, /* 2250 */
128'hc0ef855e85cea95fc0efe432854a0556, /* 2251 */
128'he91d89aa81dff0ef852285a66622a8df, /* 2252 */
128'hc0efa0a5051300003517f94c19e30c05, /* 2253 */
128'h7a4279e2690664a6854e644660e6a6df, /* 2254 */
128'he29ce31c808261256c426be27b027aa2, /* 2255 */
128'h351784aaf4a67119bff159fdb74d0605, /* 2256 */
128'he4d6e8d2eccef0caf8a293a505130000, /* 2257 */
128'h892eec6efc86f06af466f862fc5ee0da, /* 2258 */
128'h920a0a1300003a17a17fc0ef44018b32, /* 2259 */
128'h0c13498507f00b93928c8c9300003c97, /* 2260 */
128'h855208000a93926d0d1300003d1703f0, /* 2261 */
128'h408b873b9e3fc0ef856685a29ebfc0ef, /* 2262 */
128'h86b3003617934601008995b300e99733, /* 2263 */
128'h9bffc0efe432855205661a6397ca00f4, /* 2264 */
128'hf0ef852685ca66229b7fc0ef856a85a2, /* 2265 */
128'h00003517fb541be32405e1398daaf46f, /* 2266 */
128'h74a6856e744670e6997fc0ef93450513, /* 2267 */
128'h7ca27c427be26b066aa66a4669e67906, /* 2268 */
128'he28ce38c008c6663808261096de27d02, /* 2269 */
128'h7119b7f15dfdbfe5e298e398bf610605, /* 2270 */
128'hf0caf8a2854505130000351784aaf4a6, /* 2271 */
128'hf06af466f862fc5ee0dae4d6e8d2ecce, /* 2272 */
128'h3a17931fc0ef44018b32892eec6efc86, /* 2273 */
128'h0b93842c8c9300003c9783aa0a130000, /* 2274 */
128'h840d0d1300003d1703f00c13498507f0, /* 2275 */
128'hc0ef856685a2905fc0ef855208000a93, /* 2276 */
128'hc793008996b300f997b3408b87bb8fdf, /* 2277 */
128'h00e485b3003617134601fff6c693fff7, /* 2278 */
128'h85a28d1fc0efe432855205661a63974a, /* 2279 */
128'he58ff0ef852685ca66228c9fc0ef856a, /* 2280 */
128'h051300003517fb5417e32405e1398daa, /* 2281 */
128'h790674a6856e744670e68a9fc0ef8465, /* 2282 */
128'h7d027ca27c427be26b066aa66a4669e6, /* 2283 */
128'h0605e194e314008c6663808261096de2, /* 2284 */
128'hf4a67119b7f15dfdbfe5e19ce31cbf61, /* 2285 */
128'heccef0caf8a2766505130000251784aa, /* 2286 */
128'hfc86f06af466f862fc5ee0dae4d6e8d2, /* 2287 */
128'h00002997843fc0ef44018a32892eec6e, /* 2288 */
128'h07f00a93754c0c1300002c1774c98993, /* 2289 */
128'h8c9300002c9703f00b9308100b134d05, /* 2290 */
128'h80ffc0ef856285a2817fc0ef854e74ec, /* 2291 */
128'h00ed173300fd17b3408b07bb408a873b, /* 2292 */
128'h8fd5008d16b300fd17b30024079b8f5d, /* 2293 */
128'h8533003616934601fff7c313fff74893, /* 2294 */
128'hfcefc0efe432854e05461c6396ca00d4, /* 2295 */
128'hf0ef852685ca6622fc6fc0ef856685a2, /* 2296 */
128'hf8f41be3080007932405ed298daad56f, /* 2297 */
128'h744670e6fa2fc0ef7405051300002517, /* 2298 */
128'h7be26b066aa66a4669e6790674a6856e, /* 2299 */
128'h00167813808261096de27d027ca27c42, /* 2300 */
128'he10ce28c85be00081363859a008bea63, /* 2301 */
128'h5dfdbfc585bafe081be385c6b7610605, /* 2302 */
128'h6505051300002517892af0ca7119bf75, /* 2303 */
128'hf8a2fc86ec6ef06af466fc5ee8d2ecce, /* 2304 */
128'hc0ef4b81e03289aef862e0dae4d6f4a6, /* 2305 */
128'h8c9300002c97636a0a1300002a17f2cf, /* 2306 */
128'h9c3347854da1646d0d1300002d1763ec, /* 2307 */
128'h8b3bf00fc0ef85524401003b949b0177, /* 2308 */
128'h4601fffc4a93ef4fc0ef856685da0084, /* 2309 */
128'h06f61063974e00e90833003617136782, /* 2310 */
128'hecefc0ef856a85daed6fc0efe4328552, /* 2311 */
128'h2405e9318b2ac5eff0ef854a85ce6622, /* 2312 */
128'hfafb90e3040007932b85fbb41be38c56, /* 2313 */
128'h744670e6ea2fc0ef6405051300002517, /* 2314 */
128'h7be26b066aa66a4669e6790674a6855a, /* 2315 */
128'h00167513808261096de27d027ca27c42, /* 2316 */
128'hb749060500b83023e30c85d6e11185e2, /* 2317 */
128'h892e84aaf4cef8cafca67175b7e95b7d, /* 2318 */
128'he0e2e4dee8daecd6f0d2698502000513, /* 2319 */
128'hf0ef4a81e032f46ef86ae122e506fc66, /* 2320 */
128'h9c49899317cc0c1300003c174a01892f, /* 2321 */
128'h4d214d818bca8b26938c8c9300003c97, /* 2322 */
128'h85ca866e04fd956396da003d96936782, /* 2323 */
128'h2517020a0863ed45842aba2ff0ef8526, /* 2324 */
128'h640a60aa8522df4fc0ef5ba505130000, /* 2325 */
128'h6c066ba66b466ae67a0679a6794674e6, /* 2326 */
128'h8ba68b4a4a05808261497da27d427ce2, /* 2327 */
128'he82a908fe0ef842a90efe0efec36b775, /* 2328 */
128'h151b664267a28fcfe0efe42a902fe0ef, /* 2329 */
128'h9101140215028c510106161b8d5d0105, /* 2330 */
128'h4781e2880ca7be23000037978d4166e2, /* 2331 */
128'hf693078500fb86330006c683018786b3, /* 2332 */
128'h0ba1033df7b3ffa795e300d600230ff6, /* 2333 */
128'h00078a9b001a879bfbdfe0ef4521ef91, /* 2334 */
128'hbf0d0d85fa9fe0ef0007c50397e68b8d, /* 2335 */
128'h89ae892af0d2f4cef8ca7175bfa1547d, /* 2336 */
128'he0e2e4dee8daecd6fca66a0502000513, /* 2337 */
128'he0ef4b018cb2f46ee122e506f86afc66, /* 2338 */
128'h9c4a0a1306448493000034974a81f73f, /* 2339 */
128'h97934d818c4e8bca818d0d1300003d17, /* 2340 */
128'h85ce866e059d956397de00fc06b3003d, /* 2341 */
128'h2517020a8863e579842aa82ff0ef854a, /* 2342 */
128'h640a60aa8522cd4fc0ef49a505130000, /* 2343 */
128'h6c066ba66b466ae67a0679a6794674e6, /* 2344 */
128'h8c4a8bce4a85808261497da27d427ce2, /* 2345 */
128'hfe7fd0ef842afedfd0efe836ec3eb775, /* 2346 */
128'h67026622fdbfd0efe02afe1fd0efe42a, /* 2347 */
128'h140215028c518d590106161b0105151b, /* 2348 */
128'h66c267e2fca7b223000037978d419101, /* 2349 */
128'hd78300f6902393c117c20004d783e388, /* 2350 */
128'h17c20044d78300f6912393c117c20024, /* 2351 */
128'h932393c117c20064d78300f6922393c1, /* 2352 */
128'h079be87fe0ef4521ef91034df7b300f6, /* 2353 */
128'he0ef0007c50397ea8b8d00078b1b001b, /* 2354 */
128'h717580826505b789547dbf290d85e73f, /* 2355 */
128'h84ae842afca6e122fff586138932f8ca, /* 2356 */
128'hf0d2f4ce3bc505130000251785aa962a, /* 2357 */
128'he506f46ef86afc66e0e2e4dee8daecd6, /* 2358 */
128'he83e0014d9930044d793bd8fc0efec36, /* 2359 */
128'h00002b1744854a81e43e99a20034d793, /* 2360 */
128'h00002c173a4b8b9300002b973a4b0b13, /* 2361 */
128'h00002d173a4c8c9300002c973a4c0c13, /* 2362 */
128'h00003a173acd8d9300002d973acd0d13, /* 2363 */
128'h3a0505130000251702997863ebca0a13, /* 2364 */
128'h79a6794674e68556640a60aab7afc0ef, /* 2365 */
128'h7da27d427ce26c066ba66b466ae67a06, /* 2366 */
128'h00090663b52fc0ef855a85a680826149, /* 2367 */
128'h85e6b40fc0ef8562b46fc0ef855e85ca, /* 2368 */
128'hed15920ff0ef852265a2b38fc0ef856a, /* 2369 */
128'h02f749636762010a2783b28fc0ef856e, /* 2370 */
128'hc0ef3225051300002517c58d000a3583, /* 2371 */
128'h25179782852285ce6642008a3783b0cf, /* 2372 */
128'h2517b7e94a89af4fc0ef312505130000, /* 2373 */
128'h7179bfa10485ae4fc0ef0ca505130000, /* 2374 */
128'he84aec26f022f4063005051300002517, /* 2375 */
128'h05130000251704000593c19fe0efe44e, /* 2376 */
128'hc0ef31a5051300002517ab8fc0ef2fe5, /* 2377 */
128'h2517aa0fc0ef33e5051300002517aacf, /* 2378 */
128'h99934441a92fc0ef448507a505130000, /* 2379 */
128'h0135853346054685008495b3497901f4, /* 2380 */
128'h64e2740270a2ff2417e3e6dff0ef2405, /* 2381 */
128'h00c5131b460580828082614569a26942, /* 2382 */
128'h081387f245a901f61e13468148814701, /* 2383 */
128'h802397aa0007802397aa000780234000, /* 2384 */
128'hfe0813e397aa387d0007802397aa0007, /* 2385 */
128'hc00026f38e15c020267302b71d632705, /* 2386 */
128'h4000059302a68733411686b33e800513, /* 2387 */
128'h02a7473302a767b302b345bb02c74733, /* 2388 */
128'hfac710e39f2fc06f2d85051300002517, /* 2389 */
128'h4501e4061141bf51c00028f3c02026f3, /* 2390 */
128'hf6fff0ef4509f75ff0ef4505f7bff0ef, /* 2391 */
128'hf0ef4541f63ff0ef4521f69ff0ef4511, /* 2392 */
128'h8082e388400007b791011502bff1f5df, /* 2393 */
128'hb823400007b7808225016388400007b7, /* 2394 */
128'h25017b88400007b7808225016b880007, /* 2395 */
128'h400007b70106161b8d5d0085979b8082, /* 2396 */
128'h00b7ef634000073747812581f7888d51, /* 2397 */
128'h37fdc3198b097a98400006b73e800793, /* 2398 */
128'h27850006e60380827388400007b7ffe5, /* 2399 */
128'h842a4785e406e0221141bfe1f7100691, /* 2400 */
128'hfebff0ef250135fd0045551b00b7d863, /* 2401 */
128'h00044503943e24e7879300002797883d, /* 2402 */
128'h9d3d00b007b7a1ffe06f014160a26402, /* 2403 */
128'h3007071311010085151b67050185579b, /* 2404 */
128'h46010034842ec62ae8228fd905856513, /* 2405 */
128'h00344589f5bff0efec06c43e454d4589, /* 2406 */
128'h57610380079385a2f4fff0ef454d4601, /* 2407 */
128'hfee79ae3058537e100d5802300f556b3, /* 2408 */
128'hf84afc26e0a2715d80826105644260e2, /* 2409 */
128'h440189328a2e84aae486ec56f052f44e, /* 2410 */
128'h033466630144053b40000ab7ff86099b, /* 2411 */
128'h8526002c16024089063bf79ff0ef002c, /* 2412 */
128'h79a2794274e2640660a6ecbfd0ef9201, /* 2413 */
128'h2421f51ff0ef85a6808261616ae27a02, /* 2414 */
128'hbf6d00fab02304a19381178200c4579b, /* 2415 */
128'h83efc0efe406ce650513000025171141, /* 2416 */
128'h00055c63d7ff70eff885051300000517, /* 2417 */
128'h0141cda505130000251740a005b360a2, /* 2418 */
128'h00002517b4ffe06f014160a281afc06f, /* 2419 */
128'hf426f822fc067139957fe06f1ec50513, /* 2420 */
128'h251790ffe0efe05ae456e852ec4ef04a, /* 2421 */
128'h080009b74401935fe0ef12a505130000, /* 2422 */
128'h078e013407b344951289091300002917, /* 2423 */
128'h16e3fc1fb0ef0405854a0004059b6390, /* 2424 */
128'h2c8b0b1300002b174901deaf80effe94, /* 2425 */
128'h00002a17104a8a9300002a97400004b7, /* 2426 */
128'h85560007c783016907b34991114a0a13, /* 2427 */
128'hb0ef8622240125816080608ce09c0905, /* 2428 */
128'hf6ffb0ef25818552688c0004b823f7df, /* 2429 */
128'h646347190054579b0ff47413fd391be3, /* 2430 */
128'h439c97ba078a69e707130000071702f7, /* 2431 */
128'hf3ffb0ef0d45051300002517878297ba, /* 2432 */
128'h0d05051300002517a001aa9fe0ef8522, /* 2433 */
128'h00002517b7f5edbff0ef8522f2bfb0ef, /* 2434 */
128'h2517bfe9c37ff0eff17fb0ef0cc50513, /* 2435 */
128'hb7e1e14f80eff05fb0ef0ca505130000, /* 2436 */
128'hd0fff0efef3fb0ef0c85051300002517, /* 2437 */
128'h0000000000000000000000000000bf5d, /* 2438 */
128'h00000000000000000000000000000000, /* 2439 */
128'h00000000000000000000000000000000, /* 2440 */
128'h00000000000000000000000000000000, /* 2441 */
128'h00000000000000000000000000000000, /* 2442 */
128'h00000000000000000000000000000000, /* 2443 */
128'h00000000000000000000000000000000, /* 2444 */
128'h00000000000000000000000000000000, /* 2445 */
128'h00000000000000000000000000000000, /* 2446 */
128'h00000000000000000000000000000000, /* 2447 */
128'h08082828282828080808080808080808, /* 2448 */
128'h08080808080808080808080808080808, /* 2449 */
128'h101010101010101010101010101010a0, /* 2450 */
128'h10101010101004040404040404040404, /* 2451 */
128'h01010101010101010141414141414110, /* 2452 */
128'h10101010100101010101010101010101, /* 2453 */
128'h02020202020202020242424242424210, /* 2454 */
128'h08101010100202020202020202020202, /* 2455 */
128'h00000000000000000000000000000000, /* 2456 */
128'h00000000000000000000000000000000, /* 2457 */
128'h101010101010101010101010101010a0, /* 2458 */
128'h10101010101010101010101010101010, /* 2459 */
128'h01010101010101010101010101010101, /* 2460 */
128'h02010101010101011001010101010101, /* 2461 */
128'h02020202020202020202020202020202, /* 2462 */
128'h02020202020202021002020202020202, /* 2463 */
128'hc1bdceee242070dbe8c7b756d76aa478, /* 2464 */
128'hfd469501a83046134787c62af57c0faf, /* 2465 */
128'h895cd7beffff5bb18b44f7af698098d8, /* 2466 */
128'h49b40821a679438efd9871936b901122, /* 2467 */
128'he9b6c7aa265e5a51c040b340f61e2562, /* 2468 */
128'he7d3fbc8d8a1e68102441453d62f105d, /* 2469 */
128'h455a14edf4d50d87c33707d621e1cde6, /* 2470 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /* 2471 */
128'hfde5380c6d9d61228771f681fffa3942, /* 2472 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /* 2473 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /* 2474 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /* 2475 */
128'hfc93a039ab9423a7432aff97f4292244, /* 2476 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /* 2477 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /* 2478 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /* 2479 */
128'h0c07020d08030e09040f0a05000b0601, /* 2480 */
128'h020f0c090603000d0a0704010e0b0805, /* 2481 */
128'h09020b040d060f08010a030c050e0700, /* 2482 */
128'h6c5f7465735f64735f63736972776f6c, /* 2483 */
128'h6e67696c615f64730000000000006465, /* 2484 */
128'h645f6b6c635f64730000000000000000, /* 2485 */
128'h69747465735f64730000000000007669, /* 2486 */
128'h735f646d635f6473000000000000676e, /* 2487 */
128'h74657365725f64730000000074726174, /* 2488 */
128'h6e636b6c625f64730000000000000000, /* 2489 */
128'h69736b6c625f64730000000000000074, /* 2490 */
128'h6f656d69745f6473000000000000657a, /* 2491 */
128'h655f7172695f64730000000000007475, /* 2492 */
128'h5f63736972776f6c000000000000006e, /* 2493 */
128'h00000000646d635f74726174735f6473, /* 2494 */
128'h746e695f746961775f63736972776f6c, /* 2495 */
128'h000000000067616c665f747075727265, /* 2496 */
128'h00007172695f64735f63736972776f6c, /* 2497 */
128'h695f646d635f64735f63736972776f6c, /* 2498 */
128'h5f63736972776f6c0000000000007172, /* 2499 */
128'h007172695f646e655f617461645f6473, /* 2500 */
128'h0000000087fe9c880000000087feaf50, /* 2501 */
128'h004c4b40004c4b400030000020000000, /* 2502 */
128'h6d6d5f6472616f62000000020000ffff, /* 2503 */
128'h0000000087fe4e4e0064637465675f63, /* 2504 */
128'h0000000087fe4cba0000000087fe4a5c, /* 2505 */
128'h00000000000000000000000000000000, /* 2506 */
128'hffffbb30ffffbb2cffffbb2cffffbb06, /* 2507 */
128'hffffbb34ffffbb34ffffbb34ffffbb34, /* 2508 */
128'h0000000087feb2780000000087feb268, /* 2509 */
128'h0000000087feb2a00000000087feb288, /* 2510 */
128'h0000000087feb2d00000000087feb2b8, /* 2511 */
128'h0000000087feb3000000000087feb2e8, /* 2512 */
128'h0000000087feb3300000000087feb318, /* 2513 */
128'h0000000087feb3600000000087feb348, /* 2514 */
128'h40040300400402004004010040040000, /* 2515 */
128'h40050000400405004004040140040400, /* 2516 */
128'h30000000000000030000000040050100, /* 2517 */
128'h60000000000000053000000000000001, /* 2518 */
128'h70000000000000027000000000000004, /* 2519 */
128'h00000001400000007000000000000000, /* 2520 */
128'h00000005000000012000000000000006, /* 2521 */
128'h20000000000000020000000040000000, /* 2522 */
128'h00000000100000000000000100000000, /* 2523 */
128'h1e19140f0d0c0a000000000000000000, /* 2524 */
128'h000186a00000271050463c37322d2823, /* 2525 */
128'h017d7840017d784000989680000f4240, /* 2526 */
128'h031975000319750002faf080018cba80, /* 2527 */
128'h02faf08005f5e10002faf080017d7840, /* 2528 */
128'h00000020000000000bebc2000c65d400, /* 2529 */
128'h00000200000001000000008000000040, /* 2530 */
128'h00002000000010000000080000000400, /* 2531 */
128'h0000c000000080000000600000004000, /* 2532 */
128'h37363534333231300002000000010000, /* 2533 */
128'h2043534952776f4c4645444342413938, /* 2534 */
128'h746f6f622d7520646573696d696e696d, /* 2535 */
128'h00000000647261432d445320726f6620, /* 2536 */
128'hfffff986fffff99cfffff988fffff974, /* 2537 */
128'h00000000fffff9c0fffff986fffff9ae, /* 2538 */
128'he00600003800000039080000edfe0dd0, /* 2539 */
128'h00000000100000001100000028000000, /* 2540 */
128'h0000000000000000a806000059010000, /* 2541 */
128'h00000000010000000000000000000000, /* 2542 */
128'h02000000000000000400000003000000, /* 2543 */
128'h020000000f0000000400000003000000, /* 2544 */
128'h2c6874651b0000001400000003000000, /* 2545 */
128'h007665642d657261622d656e61697261, /* 2546 */
128'h2c687465260000001000000003000000, /* 2547 */
128'h0100000000657261622d656e61697261, /* 2548 */
128'h1a0000000300000000006e65736f6863, /* 2549 */
128'h303140747261752f636f732f2c000000, /* 2550 */
128'h0000003030323531313a303030303030, /* 2551 */
128'h00000000737570630100000002000000, /* 2552 */
128'h01000000000000000400000003000000, /* 2553 */
128'h000000000f0000000400000003000000, /* 2554 */
128'h40787d01380000000400000003000000, /* 2555 */
128'h03000000000000304075706301000000, /* 2556 */
128'h0300000080f0fa024b00000004000000, /* 2557 */
128'h03000000007570635b00000004000000, /* 2558 */
128'h03000000000000006700000004000000, /* 2559 */
128'h0000000079616b6f6b00000005000000, /* 2560 */
128'h7a6874651b0000001300000003000000, /* 2561 */
128'h0000766373697200656e61697261202c, /* 2562 */
128'h34367672720000000b00000003000000, /* 2563 */
128'h0b000000030000000000636466616d69, /* 2564 */
128'h0000393376732c76637369727c000000, /* 2565 */
128'h01000000850000000000000003000000, /* 2566 */
128'h6f72746e6f632d747075727265746e69, /* 2567 */
128'h04000000030000000000000072656c6c, /* 2568 */
128'h0000000003000000010000008f000000, /* 2569 */
128'h1b0000000f00000003000000a0000000, /* 2570 */
128'h000063746e692d7570632c7663736972, /* 2571 */
128'h01000000b50000000400000003000000, /* 2572 */
128'h01000000bb0000000400000003000000, /* 2573 */
128'h01000000020000000200000002000000, /* 2574 */
128'h0030303030303030384079726f6d656d, /* 2575 */
128'h6f6d656d5b0000000700000003000000, /* 2576 */
128'h67000000100000000300000000007972, /* 2577 */
128'h00000008000000000000008000000000, /* 2578 */
128'h0300000000636f730100000002000000, /* 2579 */
128'h03000000020000000000000004000000, /* 2580 */
128'h03000000020000000f00000004000000, /* 2581 */
128'h616972612c6874651b0000001f000000, /* 2582 */
128'h706d697300636f732d657261622d656e, /* 2583 */
128'h000000000300000000007375622d656c, /* 2584 */
128'h303240746e696c6301000000c3000000, /* 2585 */
128'h0d000000030000000000003030303030, /* 2586 */
128'h30746e696c632c76637369721b000000, /* 2587 */
128'hca000000100000000300000000000000, /* 2588 */
128'h07000000010000000300000001000000, /* 2589 */
128'h00000000670000001000000003000000, /* 2590 */
128'h0300000000000c000000000000000002, /* 2591 */
128'h006c6f72746e6f63de00000008000000, /* 2592 */
128'h7075727265746e690100000002000000, /* 2593 */
128'h3030634072656c6c6f72746e6f632d74, /* 2594 */
128'h04000000030000000000000030303030, /* 2595 */
128'h04000000030000000000000000000000, /* 2596 */
128'h0c00000003000000010000008f000000, /* 2597 */
128'h003063696c702c76637369721b000000, /* 2598 */
128'h03000000a00000000000000003000000, /* 2599 */
128'h0b00000001000000ca00000010000000, /* 2600 */
128'h10000000030000000900000001000000, /* 2601 */
128'h000000000000000c0000000067000000, /* 2602 */
128'he8000000040000000300000000000004, /* 2603 */
128'hfb000000040000000300000007000000, /* 2604 */
128'hb5000000040000000300000003000000, /* 2605 */
128'hbb000000040000000300000002000000, /* 2606 */
128'h75626564010000000200000002000000, /* 2607 */
128'h0000304072656c6c6f72746e6f632d67, /* 2608 */
128'h637369721b0000001000000003000000, /* 2609 */
128'h03000000003331302d67756265642c76, /* 2610 */
128'hffff000001000000ca00000008000000, /* 2611 */
128'h00000000670000001000000003000000, /* 2612 */
128'h03000000001000000000000000000000, /* 2613 */
128'h006c6f72746e6f63de00000008000000, /* 2614 */
128'h30303140747261750100000002000000, /* 2615 */
128'h08000000030000000000003030303030, /* 2616 */
128'h03000000003035373631736e1b000000, /* 2617 */
128'h00000010000000006700000010000000, /* 2618 */
128'h04000000030000000010000000000000, /* 2619 */
128'h040000000300000080f0fa024b000000, /* 2620 */
128'h040000000300000000c2010006010000, /* 2621 */
128'h04000000030000000200000014010000, /* 2622 */
128'h04000000030000000100000025010000, /* 2623 */
128'h04000000030000000200000030010000, /* 2624 */
128'h0100000002000000040000003a010000, /* 2625 */
128'h3030303240636d6d2d63736972776f6c, /* 2626 */
128'h10000000030000000000000030303030, /* 2627 */
128'h00000000000000200000000067000000, /* 2628 */
128'h14010000040000000300000000000100, /* 2629 */
128'h25010000040000000300000002000000, /* 2630 */
128'h1b0000000c0000000300000002000000, /* 2631 */
128'h0200000000636d6d2d63736972776f6c, /* 2632 */
128'h406874652d63736972776f6c01000000, /* 2633 */
128'h03000000000000003030303030303033, /* 2634 */
128'h2d63736972776f6c1b0000000c000000, /* 2635 */
128'h5b000000080000000300000000687465, /* 2636 */
128'h0400000003000000006b726f7774656e, /* 2637 */
128'h04000000030000000200000014010000, /* 2638 */
128'h06000000030000000300000025010000, /* 2639 */
128'h0300000000007fe3023e180047010000, /* 2640 */
128'h00000030000000006700000010000000, /* 2641 */
128'h01000000020000000080000000000000, /* 2642 */
128'h303440646e7277682d63736972776f6c, /* 2643 */
128'h0e000000030000000000303030303030, /* 2644 */
128'h6e7277682d63736972776f6c1b000000, /* 2645 */
128'h67000000100000000300000000000064, /* 2646 */
128'h00100000000000000000004000000000, /* 2647 */
128'h09000000020000000200000002000000, /* 2648 */
128'h2300736c6c65632d7373657264646123, /* 2649 */
128'h61706d6f6300736c6c65632d657a6973, /* 2650 */
128'h6f647473006c65646f6d00656c626974, /* 2651 */
128'h65736162656d697400687461702d7475, /* 2652 */
128'h6b636f6c630079636e6575716572662d, /* 2653 */
128'h63697665640079636e6575716572662d, /* 2654 */
128'h75746174730067657200657079745f65, /* 2655 */
128'h2d756d6d006173692c76637369720073, /* 2656 */
128'h230074696c70732d626c740065707974, /* 2657 */
128'h00736c6c65632d747075727265746e69, /* 2658 */
128'h6f72746e6f632d747075727265746e69, /* 2659 */
128'h646e6168702c78756e696c0072656c6c, /* 2660 */
128'h727265746e69007365676e617200656c, /* 2661 */
128'h6572006465646e657478652d73747075, /* 2662 */
128'h616d2c76637369720073656d616e2d67, /* 2663 */
128'h766373697200797469726f6972702d78, /* 2664 */
128'h70732d746e6572727563007665646e2c, /* 2665 */
128'h61702d747075727265746e6900646565, /* 2666 */
128'h0073747075727265746e6900746e6572, /* 2667 */
128'h6f692d6765720074666968732d676572, /* 2668 */
128'h63616d2d6c61636f6c0068746469772d, /* 2669 */
128'h0000000000000000737365726464612d, /* 2670 */
128'h0000000000203a642520656369766544, /* 2671 */
128'h00203a6425206563697665642073250a, /* 2672 */
128'h00000000203a6425206563697665440a, /* 2673 */
128'h000a656369766564206e776f6e6b6e75, /* 2674 */
128'h00000a2973252c73252870756b6f6f6c, /* 2675 */
128'h7265206c616e7265746e692070636864, /* 2676 */
128'h00000000000000000a7025202c726f72, /* 2677 */
128'h5145525f5043484420676e69646e6553, /* 2678 */
128'h4b434120504348440000000a54534555, /* 2679 */
128'h696c432050434844000000000000000a, /* 2680 */
128'h203a7373657264644120504920746e65, /* 2681 */
128'h0000000a64252e64252e64252e642520, /* 2682 */
128'h73657264644120504920726576726553, /* 2683 */
128'h0a64252e64252e64252e642520203a73, /* 2684 */
128'h6120726574756f520000000000000000, /* 2685 */
128'h252e64252e642520203a737365726464, /* 2686 */
128'h6b73616d2074654e0000000a64252e64, /* 2687 */
128'h64252e642520203a7373657264646120, /* 2688 */
128'h697420657361654c000a64252e64252e, /* 2689 */
128'h7364253a6d64253a686425203d20656d, /* 2690 */
128'h3d206e69616d6f44000000000000000a, /* 2691 */
128'h4820746e65696c4300000a2273252220, /* 2692 */
128'h000a22732522203d20656d616e74736f, /* 2693 */
128'h000000000a44455050494b53204b4341, /* 2694 */
128'h000000000000000a4b414e2050434844, /* 2695 */
128'h73657264646120646574736575716552, /* 2696 */
128'h0000000000000a646573756665722073, /* 2697 */
128'h000000000000000a732520726f727245, /* 2698 */
128'h6e6f6974706f2064656c646e61686e75, /* 2699 */
128'h656c646e61686e55000000000a642520, /* 2700 */
128'h64252065646f63706f20504348442064, /* 2701 */
128'h20676e69646e6553000000000000000a, /* 2702 */
128'h000a595245564f435349445f50434844, /* 2703 */
128'h00000000000a29732528726f72726570, /* 2704 */
128'h3a2043414d2073250000000030687465, /* 2705 */
128'h3a583230253a583230253a5832302520, /* 2706 */
128'h000a583230253a583230253a58323025, /* 2707 */
128'h484420646e65732074276e646c756f43, /* 2708 */
128'h206e6f20595245564f43534944205043, /* 2709 */
128'h00000a7325203a732520656369766564, /* 2710 */
128'h5043484420726f6620676e6974696157, /* 2711 */
128'h2020202020202020000a524546464f5f, /* 2712 */
128'h00000000000063250000000000000020, /* 2713 */
128'h0000005832302520000000000000002e, /* 2714 */
128'h00000000732573250000000000000a0a, /* 2715 */
128'h00000000007325203a646c697542202c, /* 2716 */
128'h73257a4820756c250000000000007325, /* 2717 */
128'h0000000000756c250000000000000000, /* 2718 */
128'h0073257a4863252000000000646c252e, /* 2719 */
128'h00000000007325736574794220756c25, /* 2720 */
128'h00003a786c3830250073254269632520, /* 2721 */
128'h000a73252020202000786c6c2a302520, /* 2722 */
128'h000000203a5d64255b6e6f6974636553, /* 2723 */
128'h727265207974696e6173207264646170, /* 2724 */
128'h2c7825286e666c6500000a702520726f, /* 2725 */
128'h000000000a3b29782578302c78257830, /* 2726 */
128'h782578302c302c7825287465736d656d, /* 2727 */
128'h464f5f4f4c43414d00000000000a3b29, /* 2728 */
128'h464f5f494843414d0000000054455346, /* 2729 */
128'h46464f5f524c50540000000054455346, /* 2730 */
128'h46464f5f534346540000000000544553, /* 2731 */
128'h4c5254434f49444d0000000000544553, /* 2732 */
128'h46464f5f534346520054455346464f5f, /* 2733 */
128'h5346464f5f5253520000000000544553, /* 2734 */
128'h46464f5f444142520000000000005445, /* 2735 */
128'h46464f5f524c50520000000000544553, /* 2736 */
128'h000000003f3f3f3f0000000000544553, /* 2737 */
128'h000064252b54455346464f5f524c5052, /* 2738 */
128'h6f746f72502050490000000000000047, /* 2739 */
128'h00000000000000000a50495049203d20, /* 2740 */
128'h6f746f72502050490000000000000054, /* 2741 */
128'h6f746f7250205049000a504745203d20, /* 2742 */
128'h6165682074736574000a505550203d20, /* 2743 */
128'h6e6f6320747365740000000a3a726564, /* 2744 */
128'h6f746f7250205049000a3a73746e6574, /* 2745 */
128'h6f746f7250205049000a504449203d20, /* 2746 */
128'h6f746f725020504900000a5054203d20, /* 2747 */
128'h00000000000000000a50434344203d20, /* 2748 */
128'h6f746f72502050490000000000000036, /* 2749 */
128'h00000000000000000a50565352203d20, /* 2750 */
128'h000a455247203d206f746f7250205049, /* 2751 */
128'h000a505345203d206f746f7250205049, /* 2752 */
128'h00000a4841203d206f746f7250205049, /* 2753 */
128'h000a50544d203d206f746f7250205049, /* 2754 */
128'h5054454542203d206f746f7250205049, /* 2755 */
128'h6f746f72502050490000000000000a48, /* 2756 */
128'h000000000000000a5041434e45203d20, /* 2757 */
128'h6f746f7250205049000000000000004d, /* 2758 */
128'h00000000000000000a504d4f43203d20, /* 2759 */
128'h0a50544353203d206f746f7250205049, /* 2760 */
128'h6f746f72502050490000000000000000, /* 2761 */
128'h00000000000a4554494c504455203d20, /* 2762 */
128'h0a534c504d203d206f746f7250205049, /* 2763 */
128'h6f746f72502050490000000000000000, /* 2764 */
128'h6f746f7270205049000a574152203d20, /* 2765 */
128'h2820646574726f707075736e75203d20, /* 2766 */
128'h79745f6f746f7270000000000a297825, /* 2767 */
128'h0000000000000a78257830203d206570, /* 2768 */
128'h727265746e692064656c646e61686e75, /* 2769 */
128'h414d2070757465530000000a21747075, /* 2770 */
128'h4d454f2049505351000a726464612043, /* 2771 */
128'h0000000000000a7825203d205d64255b, /* 2772 */
128'h00000a786c253a786c25203d2043414d, /* 2773 */
128'h3025203d20737365726464612043414d, /* 2774 */
128'h3230253a783230253a783230253a7832, /* 2775 */
128'h0000000a2e783230253a783230253a78, /* 2776 */
128'h00007f7c5d5b3f3e3d3c3b3a2c2b2a22, /* 2777 */
128'h007f7c5d5b3f3e3d3c3b3a2e2c2b2a22, /* 2778 */
128'h66656463626139383736353433323130, /* 2779 */
128'h72776f6c2f6372730000000000000000, /* 2780 */
128'h00000000000000632e636d6d5f637369, /* 2781 */
128'h61625f6473203d3d20657361625f6473, /* 2782 */
128'h5f63736972776f6c00726464615f6573, /* 2783 */
128'h000a74756f656d6974207325203a6473, /* 2784 */
128'h616d202c6465766f6d65722064726143, /* 2785 */
128'h6425206f74206465676e616863206b73, /* 2786 */
128'h736e692064726143000000000000000a, /* 2787 */
128'h6e616863206b73616d202c6465747265, /* 2788 */
128'h0000000000000a6425206f7420646567, /* 2789 */
128'h25207461206465746165726320636d6d, /* 2790 */
128'h0000000a7825203d2074736f68202c78, /* 2791 */
128'h0000000000006f4e0000000000736559, /* 2792 */
128'h002020203a434d4d0000000052444420, /* 2793 */
128'h00000000000a7325203a656369766544, /* 2794 */
128'h3a4449207265727574636166756e614d, /* 2795 */
128'h0a7825203a4d454f000000000a782520, /* 2796 */
128'h6325203a656d614e0000000000000000, /* 2797 */
128'h0000000000000a206325632563256325, /* 2798 */
128'h00000a6425203a646565705320737542, /* 2799 */
128'h25203a79746963617061432068676948, /* 2800 */
128'h79746963617061430000000000000a73, /* 2801 */
128'h7464695720737542000000000000203a, /* 2802 */
128'h000000000a73257469622d6425203a68, /* 2803 */
128'h0000007825782520000000203a78250a, /* 2804 */
128'h00000000000064735f63736972776f6c, /* 2805 */
128'h0000000065646f6d206e776f6e6b6e55, /* 2806 */
128'h7830203a726f72724520737574617453, /* 2807 */
128'h2074756f656d69540000000a58383025, /* 2808 */
128'h616572206472616320676e6974696177, /* 2809 */
128'h6c69616620636d6d00000000000a7964, /* 2810 */
128'h6d6320706f747320646e6573206f7420, /* 2811 */
128'h6f6c62203a434d4d0000000000000a64, /* 2812 */
128'h20786c257830207265626d756e206b63, /* 2813 */
128'h6c2578302878616d2073646565637865, /* 2814 */
128'h203d3e20434d4d6500000000000a2978, /* 2815 */
128'h726f6620646572697571657220342e34, /* 2816 */
128'h642072657375206465636e61686e6520, /* 2817 */
128'h000000000000000a6165726120617461, /* 2818 */
128'h757320746f6e2073656f642064726143, /* 2819 */
128'h696e6f697469747261702074726f7070, /* 2820 */
128'h656f64206472614300000000000a676e, /* 2821 */
128'h20434820656e6966656420746f6e2073, /* 2822 */
128'h00000a657a69732070756f7267205057, /* 2823 */
128'h636e61686e6520617461642072657355, /* 2824 */
128'h5720434820746f6e2061657261206465, /* 2825 */
128'h696c6120657a69732070756f72672050, /* 2826 */
128'h72617020692550470000000a64656e67, /* 2827 */
128'h505720434820746f6e206e6f69746974, /* 2828 */
128'h67696c6120657a69732070756f726720, /* 2829 */
128'h656f642064726143000000000a64656e, /* 2830 */
128'h6e652074726f7070757320746f6e2073, /* 2831 */
128'h657475626972747461206465636e6168, /* 2832 */
128'h6e65206c61746f54000000000000000a, /* 2833 */
128'h6563786520657a6973206465636e6168, /* 2834 */
128'h20752528206d756d6978616d20736465, /* 2835 */
128'h656f64206472614300000a297525203e, /* 2836 */
128'h6f682074726f7070757320746f6e2073, /* 2837 */
128'h61702064656c6c6f72746e6f63207473, /* 2838 */
128'h6572206574697277206e6f6974697472, /* 2839 */
128'h6e6974746573207974696c696261696c, /* 2840 */
128'h726c61206472614300000000000a7367, /* 2841 */
128'h64656e6f697469747261702079646165, /* 2842 */
128'h206f6e203a434d4d000000000000000a, /* 2843 */
128'h0000000a746e65736572702064726163, /* 2844 */
128'h73657220746f6e206469642064726143, /* 2845 */
128'h20656761746c6f76206f7420646e6f70, /* 2846 */
128'h00000000000000000a217463656c6573, /* 2847 */
128'h7463656c6573206f7420656c62616e75, /* 2848 */
128'h00000000000000000a65646f6d206120, /* 2849 */
128'h646e756f66206473635f747865206f4e, /* 2850 */
128'h78363025206e614d0000000000000a21, /* 2851 */
128'h000000783430257834302520726e5320, /* 2852 */
128'h00000000632563256325632563256325, /* 2853 */
128'h6167656c20434d4d00000064252e6425, /* 2854 */
128'h636167654c2044530000000000007963, /* 2855 */
128'h6867694820434d4d0000000000000079, /* 2856 */
128'h0000297a484d36322820646565705320, /* 2857 */
128'h35282064656570532068676948204453, /* 2858 */
128'h6867694820434d4d000000297a484d30, /* 2859 */
128'h0000297a484d32352820646565705320, /* 2860 */
128'h7a484d32352820323552444420434d4d, /* 2861 */
128'h31524453205348550000000000000029, /* 2862 */
128'h00000000000000297a484d3532282032, /* 2863 */
128'h7a484d30352820353252445320534855, /* 2864 */
128'h35524453205348550000000000000029, /* 2865 */
128'h000000000000297a484d303031282030, /* 2866 */
128'h7a484d30352820303552444420534855, /* 2867 */
128'h31524453205348550000000000000029, /* 2868 */
128'h0000000000297a484d38303228203430, /* 2869 */
128'h0000297a484d30303228203030325348, /* 2870 */
128'h6f6e2064252065636976654420434d4d, /* 2871 */
128'h00000000000000000a646e756f662074, /* 2872 */
128'h000000000000445300000000434d4d65, /* 2873 */
128'h000000297325282000006425203a7325, /* 2874 */
128'h6e656c20656c69460000000000636d6d, /* 2875 */
128'h000000000000000a6425203d20687467, /* 2876 */
128'h0a7325203d202964252c70252835646d, /* 2877 */
128'h666c652064616f6c0000000000000000, /* 2878 */
128'h000a79726f6d656d20524444206f7420, /* 2879 */
128'h2064656c696166206461657220666c65, /* 2880 */
128'h000000646c252065646f632068746977, /* 2881 */
128'h6f6f7420687461702074736575716552, /* 2882 */
128'h00000000000a646c25202e676e6f6c20, /* 2883 */
128'h732522203a717277000000000000002f, /* 2884 */
128'h0a64253d657a69736b636f6c62202c22, /* 2885 */
128'h20657669656365520000000000000000, /* 2886 */
128'h0000000000000a2e646e6520656c6966, /* 2887 */
128'h656c6c6163207172775f656c646e6168, /* 2888 */
128'h206c6167656c6c4900000000000a2e64, /* 2889 */
128'h0a2e6e6f6974617265706f2050544654, /* 2890 */
128'h75716572206e656c0000000000000000, /* 2891 */
128'h6175746361202c5825203d2064657269, /* 2892 */
128'h000000005c2d2f7c000a7825203d206c, /* 2893 */
128'h20646564616f6c2065687420746f6f42, /* 2894 */
128'h6572646461207461206d6172676f7270, /* 2895 */
128'h000000000000000a2e2e2e7025207373, /* 2896 */
128'h445320746e756f6d206f74206c696146, /* 2897 */
128'h000000000000000a2172657669726420, /* 2898 */
128'h6e69206e69622e746f6f622064616f4c, /* 2899 */
128'h0000000000000a79726f6d656d206f74, /* 2900 */
128'h00000000000000006e69622e746f6f62, /* 2901 */
128'h62206e65706f206f742064656c696146, /* 2902 */
128'h206f74206c6961660000000a21746f6f, /* 2903 */
128'h000000000021656c69662065736f6c63, /* 2904 */
128'h6420746e756f6d75206f74206c696166, /* 2905 */
128'h20746f6f622d750a00000000216b7369, /* 2906 */
128'h67617473207473726966206465736162, /* 2907 */
128'h00000a726564616f6c20746f6f622065, /* 2908 */
128'h696166207325206e6f69747265737361, /* 2909 */
128'h696c202c732520656c6966202c64656c, /* 2910 */
128'h206e6f6974636e7566202c642520656e, /* 2911 */
128'h3a4552554c49414600000000000a7325, /* 2912 */
128'h74612078257830203d21207825783020, /* 2913 */
128'h00000a2e782578302074657366666f20, /* 2914 */
128'h7025203d203270202c7025203d203170, /* 2915 */
128'h2020202020202020000000000000000a, /* 2916 */
128'h08080808080808080000000000202020, /* 2917 */
128'h20676e69747465730000000000080808, /* 2918 */
128'h20676e69747365740000000000007525, /* 2919 */
128'h3a4552554c4941460000000000007525, /* 2920 */
128'h64612064616220656c626973736f7020, /* 2921 */
128'h666f20746120656e696c207373657264, /* 2922 */
128'h00000000000a2e782578302074657366, /* 2923 */
128'h7478656e206f7420676e697070696b53, /* 2924 */
128'h000000000000000a2e2e2e7473657420, /* 2925 */
128'h20202020200808080808080808080808, /* 2926 */
128'h08080808080808080808202020202020, /* 2927 */
128'h00000000000820080000000000000008, /* 2928 */
128'h78302073692065676e61722074736574, /* 2929 */
128'h00000000000a70257830206f74207025, /* 2930 */
128'h000000000075252f00752520706f6f4c, /* 2931 */
128'h6441206b637574530000000000000a3a, /* 2932 */
128'h0000203a732520200000007373657264, /* 2933 */
128'h00000a2e656e6f4400000000000a6b6f, /* 2934 */
128'h4d415244206c6174656d20657261420a, /* 2935 */
128'h65747365746d656d00000a7473657420, /* 2936 */
128'h20302e332e34206e6f69737265762072, /* 2937 */
128'h000000000000000a297469622d642528, /* 2938 */
128'h30322029432820746867697279706f43, /* 2939 */
128'h2073656c7261684320323130322d3130, /* 2940 */
128'h000000000000000a2e6e6f62617a6143, /* 2941 */
128'h74207265646e75206465736e6563694c, /* 2942 */
128'h50206c6172656e654720554e47206568, /* 2943 */
128'h65762065736e6563694c2063696c6275, /* 2944 */
128'h0a2e29796c6e6f282032206e6f697372, /* 2945 */
128'h5f676e696b726f770000000000000000, /* 2946 */
128'h20646c25202c424b6425203d20746573, /* 2947 */
128'h6c25202c736e6f697463757274736e69, /* 2948 */
128'h203d20495043202c73656c6379632064, /* 2949 */
128'h00000000000000000a646c252e646c25, /* 2950 */
128'h46454443424139383736353433323130, /* 2951 */
128'h6f57206f6c6c65480000000000000000, /* 2952 */
128'h205d64255b70777300000a0d21646c72, /* 2953 */
128'h73206863746977530000000a5825203d, /* 2954 */
128'h000a58252c5825203d20676e69747465, /* 2955 */
128'h5825203d2064656573206d6f646e6152, /* 2956 */
128'h0a746f6f62204453000000000000000a, /* 2957 */
128'h6f6f6220495053510000000000000000, /* 2958 */
128'h736574204d4152440000000000000a74, /* 2959 */
128'h6f6f6220505446540000000000000a74, /* 2960 */
128'h65742065686361430000000000000a74, /* 2961 */
128'h00000a0d7061727400000000000a7473, /* 2962 */
128'h00000002464c457fcccccccccccccccd, /* 2963 */
128'h1032547698badcfeefcdab8967452301, /* 2964 */
128'h5851f42d4c957f2d1000000020000000, /* 2965 */
128'haaaaaaaaaaaaaaaa5555555555555555, /* 2966 */
128'h00000000000000000000000000000000, /* 2967 */
128'h00000000000000000000000000000000, /* 2968 */
128'h00000000000000000000000000000000, /* 2969 */
128'h00000000000000000000000000000000, /* 2970 */
128'h00000000000000000000000000000000, /* 2971 */
128'h00000000000000000000000000000000, /* 2972 */
128'h00000000000000000000000000000000, /* 2973 */
128'h00000000000000000000000000000000, /* 2974 */
128'h00000000000000000000000000000000, /* 2975 */
128'h00004b4d47545045000000030f060301, /* 2976 */
128'h000000003000000000000000004b4d47, /* 2977 */
128'h00000000ffffffff0000000000000000, /* 2978 */
128'h0000646d635f6473000000000c000000, /* 2979 */
128'h00000000ffffffff00006772615f6473, /* 2980 */
128'h000000002f7c5c2d0000000087feb1f8, /* 2981 */
128'h000000060000000087feb3b0cc33aa55, /* 2982 */
128'h87fe70460000000000000000ffffffff, /* 2983 */
128'h00000000000000000000000000000000, /* 2984 */
128'h00000000000000000000000000000000, /* 2985 */
128'h00000000000000000000000000000000, /* 2986 */
128'h00000000000000000000000000000000, /* 2987 */
128'h00000000000000000000000000000000, /* 2988 */
128'h00000000000000000000000000000000, /* 2989 */
128'h00000000000000000000000000000000, /* 2990 */
128'h00000000000000000000000000000000, /* 2991 */
128'h00000000000000000000000000000000, /* 2992 */
128'h00000000000000000000000000000000, /* 2993 */
128'h00000000000000000000000000000000, /* 2994 */
128'h00000000000000000000000000000000, /* 2995 */
128'h00000000000000000000000000000000, /* 2996 */
128'h00000000000000000000000000000000, /* 2997 */
128'h00000000000000000000000000000000, /* 2998 */
128'h00000000000000000000000000000000, /* 2999 */
128'h00000000000000000000000000000000, /* 3000 */
128'h00000000000000000000000000000000, /* 3001 */
128'h00000000000000000000000000000000, /* 3002 */
128'h00000000000000000000000000000000, /* 3003 */
128'h00000000000000000000000000000000, /* 3004 */
128'h00000000000000000000000000000000, /* 3005 */
128'h00000000000000000000000000000000, /* 3006 */
128'h00000000000000000000000000000000, /* 3007 */
128'h00000000000000000000000000000000, /* 3008 */
128'h00000000000000000000000000000000, /* 3009 */
128'h00000000000000000000000000000000, /* 3010 */
128'h00000000000000000000000000000000, /* 3011 */
128'h00000000000000000000000000000000, /* 3012 */
128'h00000000000000000000000000000000, /* 3013 */
128'h00000000000000000000000000000000, /* 3014 */
128'h00000000000000000000000000000000, /* 3015 */
128'h00000000000000000000000000000000, /* 3016 */
128'h00000000000000000000000000000000, /* 3017 */
128'h00000000000000000000000000000000, /* 3018 */
128'h00000000000000000000000000000000, /* 3019 */
128'h00000000000000000000000000000000, /* 3020 */
128'h00000000000000000000000000000000, /* 3021 */
128'h00000000000000000000000000000000, /* 3022 */
128'h00000000000000000000000000000000, /* 3023 */
128'h00000000000000000000000000000000, /* 3024 */
128'h00000000000000000000000000000000, /* 3025 */
128'h00000000000000000000000000000000, /* 3026 */
128'h00000000000000000000000000000000, /* 3027 */
128'h00000000000000000000000000000000, /* 3028 */
128'h00000000000000000000000000000000, /* 3029 */
128'h00000000000000000000000000000000, /* 3030 */
128'h00000000000000000000000000000000, /* 3031 */
128'h00000000000000000000000000000000, /* 3032 */
128'h00000000000000000000000000000000, /* 3033 */
128'h00000000000000000000000000000000, /* 3034 */
128'h00000000000000000000000000000000, /* 3035 */
128'h00000000000000000000000000000000, /* 3036 */
128'h00000000000000000000000000000000, /* 3037 */
128'h00000000000000000000000000000000, /* 3038 */
128'h00000000000000000000000000000000, /* 3039 */
128'h00000000000000000000000000000000, /* 3040 */
128'h00000000000000000000000000000000, /* 3041 */
128'h00000000000000000000000000000000, /* 3042 */
128'h00000000000000000000000000000000, /* 3043 */
128'h00000000000000000000000000000000, /* 3044 */
128'h00000000000000000000000000000000, /* 3045 */
128'h00000000000000000000000000000000, /* 3046 */
128'h00000000000000000000000000000000, /* 3047 */
128'h00000000000000000000000000000000, /* 3048 */
128'h00000000000000000000000000000000, /* 3049 */
128'h00000000000000000000000000000000, /* 3050 */
128'h00000000000000000000000000000000, /* 3051 */
128'h00000000000000000000000000000000, /* 3052 */
128'h00000000000000000000000000000000, /* 3053 */
128'h00000000000000000000000000000000, /* 3054 */
128'h00000000000000000000000000000000, /* 3055 */
128'h00000000000000000000000000000000, /* 3056 */
128'h00000000000000000000000000000000, /* 3057 */
128'h00000000000000000000000000000000, /* 3058 */
128'h00000000000000000000000000000000, /* 3059 */
128'h00000000000000000000000000000000, /* 3060 */
128'h00000000000000000000000000000000, /* 3061 */
128'h00000000000000000000000000000000, /* 3062 */
128'h00000000000000000000000000000000, /* 3063 */
128'h00000000000000000000000000000000, /* 3064 */
128'h00000000000000000000000000000000, /* 3065 */
128'h00000000000000000000000000000000, /* 3066 */
128'h00000000000000000000000000000000, /* 3067 */
128'h00000000000000000000000000000000, /* 3068 */
128'h00000000000000000000000000000000, /* 3069 */
128'h00000000000000000000000000000000, /* 3070 */
128'h00000000000000000000000000000000, /* 3071 */
128'h00000000000000000000000000000000, /* 3072 */
128'h00000000000000000000000000000000, /* 3073 */
128'h00000000000000000000000000000000, /* 3074 */
128'h00000000000000000000000000000000, /* 3075 */
128'h00000000000000000000000000000000, /* 3076 */
128'h00000000000000000000000000000000, /* 3077 */
128'h00000000000000000000000000000000, /* 3078 */
128'h00000000000000000000000000000000, /* 3079 */
128'h00000000000000000000000000000000, /* 3080 */
128'h00000000000000000000000000000000, /* 3081 */
128'h00000000000000000000000000000000, /* 3082 */
128'h00000000000000000000000000000000, /* 3083 */
128'h00000000000000000000000000000000, /* 3084 */
128'h00000000000000000000000000000000, /* 3085 */
128'h00000000000000000000000000000000, /* 3086 */
128'h00000000000000000000000000000000, /* 3087 */
128'h00000000000000000000000000000000, /* 3088 */
128'h00000000000000000000000000000000, /* 3089 */
128'h00000000000000000000000000000000, /* 3090 */
128'h00000000000000000000000000000000, /* 3091 */
128'h00000000000000000000000000000000, /* 3092 */
128'h00000000000000000000000000000000, /* 3093 */
128'h00000000000000000000000000000000, /* 3094 */
128'h00000000000000000000000000000000, /* 3095 */
128'h00000000000000000000000000000000, /* 3096 */
128'h00000000000000000000000000000000, /* 3097 */
128'h00000000000000000000000000000000, /* 3098 */
128'h00000000000000000000000000000000, /* 3099 */
128'h00000000000000000000000000000000, /* 3100 */
128'h00000000000000000000000000000000, /* 3101 */
128'h00000000000000000000000000000000, /* 3102 */
128'h00000000000000000000000000000000, /* 3103 */
128'h00000000000000000000000000000000, /* 3104 */
128'h00000000000000000000000000000000, /* 3105 */
128'h00000000000000000000000000000000, /* 3106 */
128'h00000000000000000000000000000000, /* 3107 */
128'h00000000000000000000000000000000, /* 3108 */
128'h00000000000000000000000000000000, /* 3109 */
128'h00000000000000000000000000000000, /* 3110 */
128'h00000000000000000000000000000000, /* 3111 */
128'h00000000000000000000000000000000, /* 3112 */
128'h00000000000000000000000000000000, /* 3113 */
128'h00000000000000000000000000000000, /* 3114 */
128'h00000000000000000000000000000000, /* 3115 */
128'h00000000000000000000000000000000, /* 3116 */
128'h00000000000000000000000000000000, /* 3117 */
128'h00000000000000000000000000000000, /* 3118 */
128'h00000000000000000000000000000000, /* 3119 */
128'h00000000000000000000000000000000, /* 3120 */
128'h00000000000000000000000000000000, /* 3121 */
128'h00000000000000000000000000000000, /* 3122 */
128'h00000000000000000000000000000000, /* 3123 */
128'h00000000000000000000000000000000, /* 3124 */
128'h00000000000000000000000000000000, /* 3125 */
128'h00000000000000000000000000000000, /* 3126 */
128'h00000000000000000000000000000000, /* 3127 */
128'h00000000000000000000000000000000, /* 3128 */
128'h00000000000000000000000000000000, /* 3129 */
128'h00000000000000000000000000000000, /* 3130 */
128'h00000000000000000000000000000000, /* 3131 */
128'h00000000000000000000000000000000, /* 3132 */
128'h00000000000000000000000000000000, /* 3133 */
128'h00000000000000000000000000000000, /* 3134 */
128'h00000000000000000000000000000000, /* 3135 */
128'h00000000000000000000000000000000, /* 3136 */
128'h00000000000000000000000000000000, /* 3137 */
128'h00000000000000000000000000000000, /* 3138 */
128'h00000000000000000000000000000000, /* 3139 */
128'h00000000000000000000000000000000, /* 3140 */
128'h00000000000000000000000000000000, /* 3141 */
128'h00000000000000000000000000000000, /* 3142 */
128'h00000000000000000000000000000000, /* 3143 */
128'h00000000000000000000000000000000, /* 3144 */
128'h00000000000000000000000000000000, /* 3145 */
128'h00000000000000000000000000000000, /* 3146 */
128'h00000000000000000000000000000000, /* 3147 */
128'h00000000000000000000000000000000, /* 3148 */
128'h00000000000000000000000000000000, /* 3149 */
128'h00000000000000000000000000000000, /* 3150 */
128'h00000000000000000000000000000000, /* 3151 */
128'h00000000000000000000000000000000, /* 3152 */
128'h00000000000000000000000000000000, /* 3153 */
128'h00000000000000000000000000000000, /* 3154 */
128'h00000000000000000000000000000000, /* 3155 */
128'h00000000000000000000000000000000, /* 3156 */
128'h00000000000000000000000000000000, /* 3157 */
128'h00000000000000000000000000000000, /* 3158 */
128'h00000000000000000000000000000000, /* 3159 */
128'h00000000000000000000000000000000, /* 3160 */
128'h00000000000000000000000000000000, /* 3161 */
128'h00000000000000000000000000000000, /* 3162 */
128'h00000000000000000000000000000000, /* 3163 */
128'h00000000000000000000000000000000, /* 3164 */
128'h00000000000000000000000000000000, /* 3165 */
128'h00000000000000000000000000000000, /* 3166 */
128'h00000000000000000000000000000000, /* 3167 */
128'h00000000000000000000000000000000, /* 3168 */
128'h00000000000000000000000000000000, /* 3169 */
128'h00000000000000000000000000000000, /* 3170 */
128'h00000000000000000000000000000000, /* 3171 */
128'h00000000000000000000000000000000, /* 3172 */
128'h00000000000000000000000000000000, /* 3173 */
128'h00000000000000000000000000000000, /* 3174 */
128'h00000000000000000000000000000000, /* 3175 */
128'h00000000000000000000000000000000, /* 3176 */
128'h00000000000000000000000000000000, /* 3177 */
128'h00000000000000000000000000000000, /* 3178 */
128'h00000000000000000000000000000000, /* 3179 */
128'h00000000000000000000000000000000, /* 3180 */
128'h00000000000000000000000000000000, /* 3181 */
128'h00000000000000000000000000000000, /* 3182 */
128'h00000000000000000000000000000000, /* 3183 */
128'h00000000000000000000000000000000, /* 3184 */
128'h00000000000000000000000000000000, /* 3185 */
128'h00000000000000000000000000000000, /* 3186 */
128'h00000000000000000000000000000000, /* 3187 */
128'h00000000000000000000000000000000, /* 3188 */
128'h00000000000000000000000000000000, /* 3189 */
128'h00000000000000000000000000000000, /* 3190 */
128'h00000000000000000000000000000000, /* 3191 */
128'h00000000000000000000000000000000, /* 3192 */
128'h00000000000000000000000000000000, /* 3193 */
128'h00000000000000000000000000000000, /* 3194 */
128'h00000000000000000000000000000000, /* 3195 */
128'h00000000000000000000000000000000, /* 3196 */
128'h00000000000000000000000000000000, /* 3197 */
128'h00000000000000000000000000000000, /* 3198 */
128'h00000000000000000000000000000000, /* 3199 */
128'h00000000000000000000000000000000, /* 3200 */
128'h00000000000000000000000000000000, /* 3201 */
128'h00000000000000000000000000000000, /* 3202 */
128'h00000000000000000000000000000000, /* 3203 */
128'h00000000000000000000000000000000, /* 3204 */
128'h00000000000000000000000000000000, /* 3205 */
128'h00000000000000000000000000000000, /* 3206 */
128'h00000000000000000000000000000000, /* 3207 */
128'h00000000000000000000000000000000, /* 3208 */
128'h00000000000000000000000000000000, /* 3209 */
128'h00000000000000000000000000000000, /* 3210 */
128'h00000000000000000000000000000000, /* 3211 */
128'h00000000000000000000000000000000, /* 3212 */
128'h00000000000000000000000000000000, /* 3213 */
128'h00000000000000000000000000000000, /* 3214 */
128'h00000000000000000000000000000000, /* 3215 */
128'h00000000000000000000000000000000, /* 3216 */
128'h00000000000000000000000000000000, /* 3217 */
128'h00000000000000000000000000000000, /* 3218 */
128'h00000000000000000000000000000000, /* 3219 */
128'h00000000000000000000000000000000, /* 3220 */
128'h00000000000000000000000000000000, /* 3221 */
128'h00000000000000000000000000000000, /* 3222 */
128'h00000000000000000000000000000000, /* 3223 */
128'h00000000000000000000000000000000, /* 3224 */
128'h00000000000000000000000000000000, /* 3225 */
128'h00000000000000000000000000000000, /* 3226 */
128'h00000000000000000000000000000000, /* 3227 */
128'h00000000000000000000000000000000, /* 3228 */
128'h00000000000000000000000000000000, /* 3229 */
128'h00000000000000000000000000000000, /* 3230 */
128'h00000000000000000000000000000000, /* 3231 */
128'h00000000000000000000000000000000, /* 3232 */
128'h00000000000000000000000000000000, /* 3233 */
128'h00000000000000000000000000000000, /* 3234 */
128'h00000000000000000000000000000000, /* 3235 */
128'h00000000000000000000000000000000, /* 3236 */
128'h00000000000000000000000000000000, /* 3237 */
128'h00000000000000000000000000000000, /* 3238 */
128'h00000000000000000000000000000000, /* 3239 */
128'h00000000000000000000000000000000, /* 3240 */
128'h00000000000000000000000000000000, /* 3241 */
128'h00000000000000000000000000000000, /* 3242 */
128'h00000000000000000000000000000000, /* 3243 */
128'h00000000000000000000000000000000, /* 3244 */
128'h00000000000000000000000000000000, /* 3245 */
128'h00000000000000000000000000000000, /* 3246 */
128'h00000000000000000000000000000000, /* 3247 */
128'h00000000000000000000000000000000, /* 3248 */
128'h00000000000000000000000000000000, /* 3249 */
128'h00000000000000000000000000000000, /* 3250 */
128'h00000000000000000000000000000000, /* 3251 */
128'h00000000000000000000000000000000, /* 3252 */
128'h00000000000000000000000000000000, /* 3253 */
128'h00000000000000000000000000000000, /* 3254 */
128'h00000000000000000000000000000000, /* 3255 */
128'h00000000000000000000000000000000, /* 3256 */
128'h00000000000000000000000000000000, /* 3257 */
128'h00000000000000000000000000000000, /* 3258 */
128'h00000000000000000000000000000000, /* 3259 */
128'h00000000000000000000000000000000, /* 3260 */
128'h00000000000000000000000000000000, /* 3261 */
128'h00000000000000000000000000000000, /* 3262 */
128'h00000000000000000000000000000000, /* 3263 */
128'h00000000000000000000000000000000, /* 3264 */
128'h00000000000000000000000000000000, /* 3265 */
128'h00000000000000000000000000000000, /* 3266 */
128'h00000000000000000000000000000000, /* 3267 */
128'h00000000000000000000000000000000, /* 3268 */
128'h00000000000000000000000000000000, /* 3269 */
128'h00000000000000000000000000000000, /* 3270 */
128'h00000000000000000000000000000000, /* 3271 */
128'h00000000000000000000000000000000, /* 3272 */
128'h00000000000000000000000000000000, /* 3273 */
128'h00000000000000000000000000000000, /* 3274 */
128'h00000000000000000000000000000000, /* 3275 */
128'h00000000000000000000000000000000, /* 3276 */
128'h00000000000000000000000000000000, /* 3277 */
128'h00000000000000000000000000000000, /* 3278 */
128'h00000000000000000000000000000000, /* 3279 */
128'h00000000000000000000000000000000, /* 3280 */
128'h00000000000000000000000000000000, /* 3281 */
128'h00000000000000000000000000000000, /* 3282 */
128'h00000000000000000000000000000000, /* 3283 */
128'h00000000000000000000000000000000, /* 3284 */
128'h00000000000000000000000000000000, /* 3285 */
128'h00000000000000000000000000000000, /* 3286 */
128'h00000000000000000000000000000000, /* 3287 */
128'h00000000000000000000000000000000, /* 3288 */
128'h00000000000000000000000000000000, /* 3289 */
128'h00000000000000000000000000000000, /* 3290 */
128'h00000000000000000000000000000000, /* 3291 */
128'h00000000000000000000000000000000, /* 3292 */
128'h00000000000000000000000000000000, /* 3293 */
128'h00000000000000000000000000000000, /* 3294 */
128'h00000000000000000000000000000000, /* 3295 */
128'h00000000000000000000000000000000, /* 3296 */
128'h00000000000000000000000000000000, /* 3297 */
128'h00000000000000000000000000000000, /* 3298 */
128'h00000000000000000000000000000000, /* 3299 */
128'h00000000000000000000000000000000, /* 3300 */
128'h00000000000000000000000000000000, /* 3301 */
128'h00000000000000000000000000000000, /* 3302 */
128'h00000000000000000000000000000000, /* 3303 */
128'h00000000000000000000000000000000, /* 3304 */
128'h00000000000000000000000000000000, /* 3305 */
128'h00000000000000000000000000000000, /* 3306 */
128'h00000000000000000000000000000000, /* 3307 */
128'h00000000000000000000000000000000, /* 3308 */
128'h00000000000000000000000000000000, /* 3309 */
128'h00000000000000000000000000000000, /* 3310 */
128'h00000000000000000000000000000000, /* 3311 */
128'h00000000000000000000000000000000, /* 3312 */
128'h00000000000000000000000000000000, /* 3313 */
128'h00000000000000000000000000000000, /* 3314 */
128'h00000000000000000000000000000000, /* 3315 */
128'h00000000000000000000000000000000, /* 3316 */
128'h00000000000000000000000000000000, /* 3317 */
128'h00000000000000000000000000000000, /* 3318 */
128'h00000000000000000000000000000000, /* 3319 */
128'h00000000000000000000000000000000, /* 3320 */
128'h00000000000000000000000000000000, /* 3321 */
128'h00000000000000000000000000000000, /* 3322 */
128'h00000000000000000000000000000000, /* 3323 */
128'h00000000000000000000000000000000, /* 3324 */
128'h00000000000000000000000000000000, /* 3325 */
128'h00000000000000000000000000000000, /* 3326 */
128'h00000000000000000000000000000000, /* 3327 */
128'h00000000000000000000000000000000, /* 3328 */
128'h00000000000000000000000000000000, /* 3329 */
128'h00000000000000000000000000000000, /* 3330 */
128'h00000000000000000000000000000000, /* 3331 */
128'h00000000000000000000000000000000, /* 3332 */
128'h00000000000000000000000000000000, /* 3333 */
128'h00000000000000000000000000000000, /* 3334 */
128'h00000000000000000000000000000000, /* 3335 */
128'h00000000000000000000000000000000, /* 3336 */
128'h00000000000000000000000000000000, /* 3337 */
128'h00000000000000000000000000000000, /* 3338 */
128'h00000000000000000000000000000000, /* 3339 */
128'h00000000000000000000000000000000, /* 3340 */
128'h00000000000000000000000000000000, /* 3341 */
128'h00000000000000000000000000000000, /* 3342 */
128'h00000000000000000000000000000000, /* 3343 */
128'h00000000000000000000000000000000, /* 3344 */
128'h00000000000000000000000000000000, /* 3345 */
128'h00000000000000000000000000000000, /* 3346 */
128'h00000000000000000000000000000000, /* 3347 */
128'h00000000000000000000000000000000, /* 3348 */
128'h00000000000000000000000000000000, /* 3349 */
128'h00000000000000000000000000000000, /* 3350 */
128'h00000000000000000000000000000000, /* 3351 */
128'h00000000000000000000000000000000, /* 3352 */
128'h00000000000000000000000000000000, /* 3353 */
128'h00000000000000000000000000000000, /* 3354 */
128'h00000000000000000000000000000000, /* 3355 */
128'h00000000000000000000000000000000, /* 3356 */
128'h00000000000000000000000000000000, /* 3357 */
128'h00000000000000000000000000000000, /* 3358 */
128'h00000000000000000000000000000000, /* 3359 */
128'h00000000000000000000000000000000, /* 3360 */
128'h00000000000000000000000000000000, /* 3361 */
128'h00000000000000000000000000000000, /* 3362 */
128'h00000000000000000000000000000000, /* 3363 */
128'h00000000000000000000000000000000, /* 3364 */
128'h00000000000000000000000000000000, /* 3365 */
128'h00000000000000000000000000000000, /* 3366 */
128'h00000000000000000000000000000000, /* 3367 */
128'h00000000000000000000000000000000, /* 3368 */
128'h00000000000000000000000000000000, /* 3369 */
128'h00000000000000000000000000000000, /* 3370 */
128'h00000000000000000000000000000000, /* 3371 */
128'h00000000000000000000000000000000, /* 3372 */
128'h00000000000000000000000000000000, /* 3373 */
128'h00000000000000000000000000000000, /* 3374 */
128'h00000000000000000000000000000000, /* 3375 */
128'h00000000000000000000000000000000, /* 3376 */
128'h00000000000000000000000000000000, /* 3377 */
128'h00000000000000000000000000000000, /* 3378 */
128'h00000000000000000000000000000000, /* 3379 */
128'h00000000000000000000000000000000, /* 3380 */
128'h00000000000000000000000000000000, /* 3381 */
128'h00000000000000000000000000000000, /* 3382 */
128'h00000000000000000000000000000000, /* 3383 */
128'h00000000000000000000000000000000, /* 3384 */
128'h00000000000000000000000000000000, /* 3385 */
128'h00000000000000000000000000000000, /* 3386 */
128'h00000000000000000000000000000000, /* 3387 */
128'h00000000000000000000000000000000, /* 3388 */
128'h00000000000000000000000000000000, /* 3389 */
128'h00000000000000000000000000000000, /* 3390 */
128'h00000000000000000000000000000000, /* 3391 */
128'h00000000000000000000000000000000, /* 3392 */
128'h00000000000000000000000000000000, /* 3393 */
128'h00000000000000000000000000000000, /* 3394 */
128'h00000000000000000000000000000000, /* 3395 */
128'h00000000000000000000000000000000, /* 3396 */
128'h00000000000000000000000000000000, /* 3397 */
128'h00000000000000000000000000000000, /* 3398 */
128'h00000000000000000000000000000000, /* 3399 */
128'h00000000000000000000000000000000, /* 3400 */
128'h00000000000000000000000000000000, /* 3401 */
128'h00000000000000000000000000000000, /* 3402 */
128'h00000000000000000000000000000000, /* 3403 */
128'h00000000000000000000000000000000, /* 3404 */
128'h00000000000000000000000000000000, /* 3405 */
128'h00000000000000000000000000000000, /* 3406 */
128'h00000000000000000000000000000000, /* 3407 */
128'h00000000000000000000000000000000, /* 3408 */
128'h00000000000000000000000000000000, /* 3409 */
128'h00000000000000000000000000000000, /* 3410 */
128'h00000000000000000000000000000000, /* 3411 */
128'h00000000000000000000000000000000, /* 3412 */
128'h00000000000000000000000000000000, /* 3413 */
128'h00000000000000000000000000000000, /* 3414 */
128'h00000000000000000000000000000000, /* 3415 */
128'h00000000000000000000000000000000, /* 3416 */
128'h00000000000000000000000000000000, /* 3417 */
128'h00000000000000000000000000000000, /* 3418 */
128'h00000000000000000000000000000000, /* 3419 */
128'h00000000000000000000000000000000, /* 3420 */
128'h00000000000000000000000000000000, /* 3421 */
128'h00000000000000000000000000000000, /* 3422 */
128'h00000000000000000000000000000000, /* 3423 */
128'h00000000000000000000000000000000, /* 3424 */
128'h00000000000000000000000000000000, /* 3425 */
128'h00000000000000000000000000000000, /* 3426 */
128'h00000000000000000000000000000000, /* 3427 */
128'h00000000000000000000000000000000, /* 3428 */
128'h00000000000000000000000000000000, /* 3429 */
128'h00000000000000000000000000000000, /* 3430 */
128'h00000000000000000000000000000000, /* 3431 */
128'h00000000000000000000000000000000, /* 3432 */
128'h00000000000000000000000000000000, /* 3433 */
128'h00000000000000000000000000000000, /* 3434 */
128'h00000000000000000000000000000000, /* 3435 */
128'h00000000000000000000000000000000, /* 3436 */
128'h00000000000000000000000000000000, /* 3437 */
128'h00000000000000000000000000000000, /* 3438 */
128'h00000000000000000000000000000000, /* 3439 */
128'h00000000000000000000000000000000, /* 3440 */
128'h00000000000000000000000000000000, /* 3441 */
128'h00000000000000000000000000000000, /* 3442 */
128'h00000000000000000000000000000000, /* 3443 */
128'h00000000000000000000000000000000, /* 3444 */
128'h00000000000000000000000000000000, /* 3445 */
128'h00000000000000000000000000000000, /* 3446 */
128'h00000000000000000000000000000000, /* 3447 */
128'h00000000000000000000000000000000, /* 3448 */
128'h00000000000000000000000000000000, /* 3449 */
128'h00000000000000000000000000000000, /* 3450 */
128'h00000000000000000000000000000000, /* 3451 */
128'h00000000000000000000000000000000, /* 3452 */
128'h00000000000000000000000000000000, /* 3453 */
128'h00000000000000000000000000000000, /* 3454 */
128'h00000000000000000000000000000000, /* 3455 */
128'h00000000000000000000000000000000, /* 3456 */
128'h00000000000000000000000000000000, /* 3457 */
128'h00000000000000000000000000000000, /* 3458 */
128'h00000000000000000000000000000000, /* 3459 */
128'h00000000000000000000000000000000, /* 3460 */
128'h00000000000000000000000000000000, /* 3461 */
128'h00000000000000000000000000000000, /* 3462 */
128'h00000000000000000000000000000000, /* 3463 */
128'h00000000000000000000000000000000, /* 3464 */
128'h00000000000000000000000000000000, /* 3465 */
128'h00000000000000000000000000000000, /* 3466 */
128'h00000000000000000000000000000000, /* 3467 */
128'h00000000000000000000000000000000, /* 3468 */
128'h00000000000000000000000000000000, /* 3469 */
128'h00000000000000000000000000000000, /* 3470 */
128'h00000000000000000000000000000000, /* 3471 */
128'h00000000000000000000000000000000, /* 3472 */
128'h00000000000000000000000000000000, /* 3473 */
128'h00000000000000000000000000000000, /* 3474 */
128'h00000000000000000000000000000000, /* 3475 */
128'h00000000000000000000000000000000, /* 3476 */
128'h00000000000000000000000000000000, /* 3477 */
128'h00000000000000000000000000000000, /* 3478 */
128'h00000000000000000000000000000000, /* 3479 */
128'h00000000000000000000000000000000, /* 3480 */
128'h00000000000000000000000000000000, /* 3481 */
128'h00000000000000000000000000000000, /* 3482 */
128'h00000000000000000000000000000000, /* 3483 */
128'h00000000000000000000000000000000, /* 3484 */
128'h00000000000000000000000000000000, /* 3485 */
128'h00000000000000000000000000000000, /* 3486 */
128'h00000000000000000000000000000000, /* 3487 */
128'h00000000000000000000000000000000, /* 3488 */
128'h00000000000000000000000000000000, /* 3489 */
128'h00000000000000000000000000000000, /* 3490 */
128'h00000000000000000000000000000000, /* 3491 */
128'h00000000000000000000000000000000, /* 3492 */
128'h00000000000000000000000000000000, /* 3493 */
128'h00000000000000000000000000000000, /* 3494 */
128'h00000000000000000000000000000000, /* 3495 */
128'h00000000000000000000000000000000, /* 3496 */
128'h00000000000000000000000000000000, /* 3497 */
128'h00000000000000000000000000000000, /* 3498 */
128'h00000000000000000000000000000000, /* 3499 */
128'h00000000000000000000000000000000, /* 3500 */
128'h00000000000000000000000000000000, /* 3501 */
128'h00000000000000000000000000000000, /* 3502 */
128'h00000000000000000000000000000000, /* 3503 */
128'h00000000000000000000000000000000, /* 3504 */
128'h00000000000000000000000000000000, /* 3505 */
128'h00000000000000000000000000000000, /* 3506 */
128'h00000000000000000000000000000000, /* 3507 */
128'h00000000000000000000000000000000, /* 3508 */
128'h00000000000000000000000000000000, /* 3509 */
128'h00000000000000000000000000000000, /* 3510 */
128'h00000000000000000000000000000000, /* 3511 */
128'h00000000000000000000000000000000, /* 3512 */
128'h00000000000000000000000000000000, /* 3513 */
128'h00000000000000000000000000000000, /* 3514 */
128'h00000000000000000000000000000000, /* 3515 */
128'h00000000000000000000000000000000, /* 3516 */
128'h00000000000000000000000000000000, /* 3517 */
128'h00000000000000000000000000000000, /* 3518 */
128'h00000000000000000000000000000000, /* 3519 */
128'h00000000000000000000000000000000, /* 3520 */
128'h00000000000000000000000000000000, /* 3521 */
128'h00000000000000000000000000000000, /* 3522 */
128'h00000000000000000000000000000000, /* 3523 */
128'h00000000000000000000000000000000, /* 3524 */
128'h00000000000000000000000000000000, /* 3525 */
128'h00000000000000000000000000000000, /* 3526 */
128'h00000000000000000000000000000000, /* 3527 */
128'h00000000000000000000000000000000, /* 3528 */
128'h00000000000000000000000000000000, /* 3529 */
128'h00000000000000000000000000000000, /* 3530 */
128'h00000000000000000000000000000000, /* 3531 */
128'h00000000000000000000000000000000, /* 3532 */
128'h00000000000000000000000000000000, /* 3533 */
128'h00000000000000000000000000000000, /* 3534 */
128'h00000000000000000000000000000000, /* 3535 */
128'h00000000000000000000000000000000, /* 3536 */
128'h00000000000000000000000000000000, /* 3537 */
128'h00000000000000000000000000000000, /* 3538 */
128'h00000000000000000000000000000000, /* 3539 */
128'h00000000000000000000000000000000, /* 3540 */
128'h00000000000000000000000000000000, /* 3541 */
128'h00000000000000000000000000000000, /* 3542 */
128'h00000000000000000000000000000000, /* 3543 */
128'h00000000000000000000000000000000, /* 3544 */
128'h00000000000000000000000000000000, /* 3545 */
128'h00000000000000000000000000000000, /* 3546 */
128'h00000000000000000000000000000000, /* 3547 */
128'h00000000000000000000000000000000, /* 3548 */
128'h00000000000000000000000000000000, /* 3549 */
128'h00000000000000000000000000000000, /* 3550 */
128'h00000000000000000000000000000000, /* 3551 */
128'h00000000000000000000000000000000, /* 3552 */
128'h00000000000000000000000000000000, /* 3553 */
128'h00000000000000000000000000000000, /* 3554 */
128'h00000000000000000000000000000000, /* 3555 */
128'h00000000000000000000000000000000, /* 3556 */
128'h00000000000000000000000000000000, /* 3557 */
128'h00000000000000000000000000000000, /* 3558 */
128'h00000000000000000000000000000000, /* 3559 */
128'h00000000000000000000000000000000, /* 3560 */
128'h00000000000000000000000000000000, /* 3561 */
128'h00000000000000000000000000000000, /* 3562 */
128'h00000000000000000000000000000000, /* 3563 */
128'h00000000000000000000000000000000, /* 3564 */
128'h00000000000000000000000000000000, /* 3565 */
128'h00000000000000000000000000000000, /* 3566 */
128'h00000000000000000000000000000000, /* 3567 */
128'h00000000000000000000000000000000, /* 3568 */
128'h00000000000000000000000000000000, /* 3569 */
128'h00000000000000000000000000000000, /* 3570 */
128'h00000000000000000000000000000000, /* 3571 */
128'h00000000000000000000000000000000, /* 3572 */
128'h00000000000000000000000000000000, /* 3573 */
128'h00000000000000000000000000000000, /* 3574 */
128'h00000000000000000000000000000000, /* 3575 */
128'h00000000000000000000000000000000, /* 3576 */
128'h00000000000000000000000000000000, /* 3577 */
128'h00000000000000000000000000000000, /* 3578 */
128'h00000000000000000000000000000000, /* 3579 */
128'h00000000000000000000000000000000, /* 3580 */
128'h00000000000000000000000000000000, /* 3581 */
128'h00000000000000000000000000000000, /* 3582 */
128'h00000000000000000000000000000000, /* 3583 */
128'h00000000000000000000000000000000, /* 3584 */
128'h00000000000000000000000000000000, /* 3585 */
128'h00000000000000000000000000000000, /* 3586 */
128'h00000000000000000000000000000000, /* 3587 */
128'h00000000000000000000000000000000, /* 3588 */
128'h00000000000000000000000000000000, /* 3589 */
128'h00000000000000000000000000000000, /* 3590 */
128'h00000000000000000000000000000000, /* 3591 */
128'h00000000000000000000000000000000, /* 3592 */
128'h00000000000000000000000000000000, /* 3593 */
128'h00000000000000000000000000000000, /* 3594 */
128'h00000000000000000000000000000000, /* 3595 */
128'h00000000000000000000000000000000, /* 3596 */
128'h00000000000000000000000000000000, /* 3597 */
128'h00000000000000000000000000000000, /* 3598 */
128'h00000000000000000000000000000000, /* 3599 */
128'h00000000000000000000000000000000, /* 3600 */
128'h00000000000000000000000000000000, /* 3601 */
128'h00000000000000000000000000000000, /* 3602 */
128'h00000000000000000000000000000000, /* 3603 */
128'h00000000000000000000000000000000, /* 3604 */
128'h00000000000000000000000000000000, /* 3605 */
128'h00000000000000000000000000000000, /* 3606 */
128'h00000000000000000000000000000000, /* 3607 */
128'h00000000000000000000000000000000, /* 3608 */
128'h00000000000000000000000000000000, /* 3609 */
128'h00000000000000000000000000000000, /* 3610 */
128'h00000000000000000000000000000000, /* 3611 */
128'h00000000000000000000000000000000, /* 3612 */
128'h00000000000000000000000000000000, /* 3613 */
128'h00000000000000000000000000000000, /* 3614 */
128'h00000000000000000000000000000000, /* 3615 */
128'h00000000000000000000000000000000, /* 3616 */
128'h00000000000000000000000000000000, /* 3617 */
128'h00000000000000000000000000000000, /* 3618 */
128'h00000000000000000000000000000000, /* 3619 */
128'h00000000000000000000000000000000, /* 3620 */
128'h00000000000000000000000000000000, /* 3621 */
128'h00000000000000000000000000000000, /* 3622 */
128'h00000000000000000000000000000000, /* 3623 */
128'h00000000000000000000000000000000, /* 3624 */
128'h00000000000000000000000000000000, /* 3625 */
128'h00000000000000000000000000000000, /* 3626 */
128'h00000000000000000000000000000000, /* 3627 */
128'h00000000000000000000000000000000, /* 3628 */
128'h00000000000000000000000000000000, /* 3629 */
128'h00000000000000000000000000000000, /* 3630 */
128'h00000000000000000000000000000000, /* 3631 */
128'h00000000000000000000000000000000, /* 3632 */
128'h00000000000000000000000000000000, /* 3633 */
128'h00000000000000000000000000000000, /* 3634 */
128'h00000000000000000000000000000000, /* 3635 */
128'h00000000000000000000000000000000, /* 3636 */
128'h00000000000000000000000000000000, /* 3637 */
128'h00000000000000000000000000000000, /* 3638 */
128'h00000000000000000000000000000000, /* 3639 */
128'h00000000000000000000000000000000, /* 3640 */
128'h00000000000000000000000000000000, /* 3641 */
128'h00000000000000000000000000000000, /* 3642 */
128'h00000000000000000000000000000000, /* 3643 */
128'h00000000000000000000000000000000, /* 3644 */
128'h00000000000000000000000000000000, /* 3645 */
128'h00000000000000000000000000000000, /* 3646 */
128'h00000000000000000000000000000000, /* 3647 */
128'h00000000000000000000000000000000, /* 3648 */
128'h00000000000000000000000000000000, /* 3649 */
128'h00000000000000000000000000000000, /* 3650 */
128'h00000000000000000000000000000000, /* 3651 */
128'h00000000000000000000000000000000, /* 3652 */
128'h00000000000000000000000000000000, /* 3653 */
128'h00000000000000000000000000000000, /* 3654 */
128'h00000000000000000000000000000000, /* 3655 */
128'h00000000000000000000000000000000, /* 3656 */
128'h00000000000000000000000000000000, /* 3657 */
128'h00000000000000000000000000000000, /* 3658 */
128'h00000000000000000000000000000000, /* 3659 */
128'h00000000000000000000000000000000, /* 3660 */
128'h00000000000000000000000000000000, /* 3661 */
128'h00000000000000000000000000000000, /* 3662 */
128'h00000000000000000000000000000000, /* 3663 */
128'h00000000000000000000000000000000, /* 3664 */
128'h00000000000000000000000000000000, /* 3665 */
128'h00000000000000000000000000000000, /* 3666 */
128'h00000000000000000000000000000000, /* 3667 */
128'h00000000000000000000000000000000, /* 3668 */
128'h00000000000000000000000000000000, /* 3669 */
128'h00000000000000000000000000000000, /* 3670 */
128'h00000000000000000000000000000000, /* 3671 */
128'h00000000000000000000000000000000, /* 3672 */
128'h00000000000000000000000000000000, /* 3673 */
128'h00000000000000000000000000000000, /* 3674 */
128'h00000000000000000000000000000000, /* 3675 */
128'h00000000000000000000000000000000, /* 3676 */
128'h00000000000000000000000000000000, /* 3677 */
128'h00000000000000000000000000000000, /* 3678 */
128'h00000000000000000000000000000000, /* 3679 */
128'h00000000000000000000000000000000, /* 3680 */
128'h00000000000000000000000000000000, /* 3681 */
128'h00000000000000000000000000000000, /* 3682 */
128'h00000000000000000000000000000000, /* 3683 */
128'h00000000000000000000000000000000, /* 3684 */
128'h00000000000000000000000000000000, /* 3685 */
128'h00000000000000000000000000000000, /* 3686 */
128'h00000000000000000000000000000000, /* 3687 */
128'h00000000000000000000000000000000, /* 3688 */
128'h00000000000000000000000000000000, /* 3689 */
128'h00000000000000000000000000000000, /* 3690 */
128'h00000000000000000000000000000000, /* 3691 */
128'h00000000000000000000000000000000, /* 3692 */
128'h00000000000000000000000000000000, /* 3693 */
128'h00000000000000000000000000000000, /* 3694 */
128'h00000000000000000000000000000000, /* 3695 */
128'h00000000000000000000000000000000, /* 3696 */
128'h00000000000000000000000000000000, /* 3697 */
128'h00000000000000000000000000000000, /* 3698 */
128'h00000000000000000000000000000000, /* 3699 */
128'h00000000000000000000000000000000, /* 3700 */
128'h00000000000000000000000000000000, /* 3701 */
128'h00000000000000000000000000000000, /* 3702 */
128'h00000000000000000000000000000000, /* 3703 */
128'h00000000000000000000000000000000, /* 3704 */
128'h00000000000000000000000000000000, /* 3705 */
128'h00000000000000000000000000000000, /* 3706 */
128'h00000000000000000000000000000000, /* 3707 */
128'h00000000000000000000000000000000, /* 3708 */
128'h00000000000000000000000000000000, /* 3709 */
128'h00000000000000000000000000000000, /* 3710 */
128'h00000000000000000000000000000000, /* 3711 */
128'h00000000000000000000000000000000, /* 3712 */
128'h00000000000000000000000000000000, /* 3713 */
128'h00000000000000000000000000000000, /* 3714 */
128'h00000000000000000000000000000000, /* 3715 */
128'h00000000000000000000000000000000, /* 3716 */
128'h00000000000000000000000000000000, /* 3717 */
128'h00000000000000000000000000000000, /* 3718 */
128'h00000000000000000000000000000000, /* 3719 */
128'h00000000000000000000000000000000, /* 3720 */
128'h00000000000000000000000000000000, /* 3721 */
128'h00000000000000000000000000000000, /* 3722 */
128'h00000000000000000000000000000000, /* 3723 */
128'h00000000000000000000000000000000, /* 3724 */
128'h00000000000000000000000000000000, /* 3725 */
128'h00000000000000000000000000000000, /* 3726 */
128'h00000000000000000000000000000000, /* 3727 */
128'h00000000000000000000000000000000, /* 3728 */
128'h00000000000000000000000000000000, /* 3729 */
128'h00000000000000000000000000000000, /* 3730 */
128'h00000000000000000000000000000000, /* 3731 */
128'h00000000000000000000000000000000, /* 3732 */
128'h00000000000000000000000000000000, /* 3733 */
128'h00000000000000000000000000000000, /* 3734 */
128'h00000000000000000000000000000000, /* 3735 */
128'h00000000000000000000000000000000, /* 3736 */
128'h00000000000000000000000000000000, /* 3737 */
128'h00000000000000000000000000000000, /* 3738 */
128'h00000000000000000000000000000000, /* 3739 */
128'h00000000000000000000000000000000, /* 3740 */
128'h00000000000000000000000000000000, /* 3741 */
128'h00000000000000000000000000000000, /* 3742 */
128'h00000000000000000000000000000000, /* 3743 */
128'h00000000000000000000000000000000, /* 3744 */
128'h00000000000000000000000000000000, /* 3745 */
128'h00000000000000000000000000000000, /* 3746 */
128'h00000000000000000000000000000000, /* 3747 */
128'h00000000000000000000000000000000, /* 3748 */
128'h00000000000000000000000000000000, /* 3749 */
128'h00000000000000000000000000000000, /* 3750 */
128'h00000000000000000000000000000000, /* 3751 */
128'h00000000000000000000000000000000, /* 3752 */
128'h00000000000000000000000000000000, /* 3753 */
128'h00000000000000000000000000000000, /* 3754 */
128'h00000000000000000000000000000000, /* 3755 */
128'h00000000000000000000000000000000, /* 3756 */
128'h00000000000000000000000000000000, /* 3757 */
128'h00000000000000000000000000000000, /* 3758 */
128'h00000000000000000000000000000000, /* 3759 */
128'h00000000000000000000000000000000, /* 3760 */
128'h00000000000000000000000000000000, /* 3761 */
128'h00000000000000000000000000000000, /* 3762 */
128'h00000000000000000000000000000000, /* 3763 */
128'h00000000000000000000000000000000, /* 3764 */
128'h00000000000000000000000000000000, /* 3765 */
128'h00000000000000000000000000000000, /* 3766 */
128'h00000000000000000000000000000000, /* 3767 */
128'h00000000000000000000000000000000, /* 3768 */
128'h00000000000000000000000000000000, /* 3769 */
128'h00000000000000000000000000000000, /* 3770 */
128'h00000000000000000000000000000000, /* 3771 */
128'h00000000000000000000000000000000, /* 3772 */
128'h00000000000000000000000000000000, /* 3773 */
128'h00000000000000000000000000000000, /* 3774 */
128'h00000000000000000000000000000000, /* 3775 */
128'h00000000000000000000000000000000, /* 3776 */
128'h00000000000000000000000000000000, /* 3777 */
128'h00000000000000000000000000000000, /* 3778 */
128'h00000000000000000000000000000000, /* 3779 */
128'h00000000000000000000000000000000, /* 3780 */
128'h00000000000000000000000000000000, /* 3781 */
128'h00000000000000000000000000000000, /* 3782 */
128'h00000000000000000000000000000000, /* 3783 */
128'h00000000000000000000000000000000, /* 3784 */
128'h00000000000000000000000000000000, /* 3785 */
128'h00000000000000000000000000000000, /* 3786 */
128'h00000000000000000000000000000000, /* 3787 */
128'h00000000000000000000000000000000, /* 3788 */
128'h00000000000000000000000000000000, /* 3789 */
128'h00000000000000000000000000000000, /* 3790 */
128'h00000000000000000000000000000000, /* 3791 */
128'h00000000000000000000000000000000, /* 3792 */
128'h00000000000000000000000000000000, /* 3793 */
128'h00000000000000000000000000000000, /* 3794 */
128'h00000000000000000000000000000000, /* 3795 */
128'h00000000000000000000000000000000, /* 3796 */
128'h00000000000000000000000000000000, /* 3797 */
128'h00000000000000000000000000000000, /* 3798 */
128'h00000000000000000000000000000000, /* 3799 */
128'h00000000000000000000000000000000, /* 3800 */
128'h00000000000000000000000000000000, /* 3801 */
128'h00000000000000000000000000000000, /* 3802 */
128'h00000000000000000000000000000000, /* 3803 */
128'h00000000000000000000000000000000, /* 3804 */
128'h00000000000000000000000000000000, /* 3805 */
128'h00000000000000000000000000000000, /* 3806 */
128'h00000000000000000000000000000000, /* 3807 */
128'h00000000000000000000000000000000, /* 3808 */
128'h00000000000000000000000000000000, /* 3809 */
128'h00000000000000000000000000000000, /* 3810 */
128'h00000000000000000000000000000000, /* 3811 */
128'h00000000000000000000000000000000, /* 3812 */
128'h00000000000000000000000000000000, /* 3813 */
128'h00000000000000000000000000000000, /* 3814 */
128'h00000000000000000000000000000000, /* 3815 */
128'h00000000000000000000000000000000, /* 3816 */
128'h00000000000000000000000000000000, /* 3817 */
128'h00000000000000000000000000000000, /* 3818 */
128'h00000000000000000000000000000000, /* 3819 */
128'h00000000000000000000000000000000, /* 3820 */
128'h00000000000000000000000000000000, /* 3821 */
128'h00000000000000000000000000000000, /* 3822 */
128'h00000000000000000000000000000000, /* 3823 */
128'h00000000000000000000000000000000, /* 3824 */
128'h00000000000000000000000000000000, /* 3825 */
128'h00000000000000000000000000000000, /* 3826 */
128'h00000000000000000000000000000000, /* 3827 */
128'h00000000000000000000000000000000, /* 3828 */
128'h00000000000000000000000000000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00000000000000000000000000000000, /* 3840 */
128'h00000000000000000000000000000000, /* 3841 */
128'h00000000000000000000000000000000, /* 3842 */
128'h00000000000000000000000000000000, /* 3843 */
128'h00000000000000000000000000000000, /* 3844 */
128'h00000000000000000000000000000000, /* 3845 */
128'h00000000000000000000000000000000, /* 3846 */
128'h00000000000000000000000000000000, /* 3847 */
128'h00000000000000000000000000000000, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule

