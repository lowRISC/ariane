/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'h01111113fff1011b0000613711249463, /*    1 */
128'h00008297000280e70f62829300008297, /*    2 */
128'h000280e7130505130000051711c28293, /*    3 */
128'hac5606130000c617fc05859300000597, /*    4 */
128'h000f4eb701169693fff6869b000066b7, /*    5 */
128'h0085b703fffe8e930005b703240e8e9b, /*    6 */
128'hff81011301b111130110011bfe0e9ae3, /*    7 */
128'h0085b70300e6b0230005b7030006b703, /*    8 */
128'h0185b70300e6b8230105b70300e6b423, /*    9 */
128'hfcc5cce3020686930205859300e6bc23, /*   10 */
128'h40b787b300d787b30147879300000797, /*   11 */
128'h30579073090787930000079700078067, /*   12 */
128'h090606130000c617b30585930000c597, /*   13 */
128'h0005bc230005b8230005b4230005b023, /*   14 */
128'h020004b765a090effec5c6e302058593, /*   15 */
128'h02000937004484930124a02300100913, /*   16 */
128'h3440297310500073ff24c6e34009091b, /*   17 */
128'hf1402973020004b7fe090ae300897913, /*   18 */
128'h0004a903000920230099093300291913, /*   19 */
128'h4009091b0200093700448493fe091ee3, /*   20 */
128'h1050007334102373342022f3ff24c6e3, /*   21 */
128'h41206d6f7266206f6c6c6548ffdff06f, /*   22 */
128'h617720657361656c502021656e616972, /*   23 */
128'h000a2e2e2e746e656d6f6d2061207469, /*   24 */
128'h00000000000000000000000000000000, /*   25 */
128'h00000000000000000000000000000000, /*   26 */
128'h00000000000000000000000000000000, /*   27 */
128'h00000000000000000000000000000000, /*   28 */
128'h00000000000000000000000000000000, /*   29 */
128'h00000000000000000000000000000000, /*   30 */
128'h00000000000000000000000000000000, /*   31 */
128'hd963454c0005cc635735c28587ae6914, /*   32 */
128'he21c97b6470102a787b30a00051300b7, /*   33 */
128'h853e85b200030563018533038082853a, /*   34 */
128'h768686930000b697b7edfda007138302, /*   35 */
128'h87930000c79762948d0707130000c717, /*   36 */
128'h87b30280069302d787bb878d8f998c67, /*   37 */
128'h47148082853a470100e7956397ba02d7, /*   38 */
128'hf0efe4061141b7f502870713fea68de3, /*   39 */
128'hbfe545018082014160a26108c509fbbf, /*   40 */
128'hf0efe852ec4ef04af426f822fc067139, /*   41 */
128'h0000ba17440144814985892acd31f9bf, /*   42 */
128'he091450100f44d6300c92783264a0a13, /*   43 */
128'h61216a4269e2790274a2744270e25535, /*   44 */
128'h67a2ed19f29ff0ef854a85a200308082, /*   45 */
128'h50ef8552000995632485cb990087c783, /*   46 */
128'h0513bf65240521a080ef4981652250e0, /*   47 */
128'hf2dff0efe42ef406f0227179b7c1fda0, /*   48 */
128'h842aee7ff0ef083065a2c105fda00413, /*   49 */
128'h00f7096300c547030ff007936562e911, /*   50 */
128'h547980826145740270a285221e0080ef, /*   51 */
128'hf0efec4ef04af426f822fc067139bfd5, /*   52 */
128'h0000a9970ff00913440184aacd01eebf, /*   53 */
128'h74a2744270e200f4496344dc3a498993, /*   54 */
128'hf0ef852685a200308082612169e27902, /*   55 */
128'h85a20127896300c7c78367a2ed09e83f, /*   56 */
128'hb7d9240517a080ef652246a050ef854e, /*   57 */
128'he8dff0ef892eec26f406e84af0227179, /*   58 */
128'he45ff0ef84aa85ca0030c11dfda00413, /*   59 */
128'h348505130000a517864a608ced01842a, /*   60 */
128'h740270a2852213c080ef652242c050ef, /*   61 */
128'hf406ec26f022717980826145694264e2, /*   62 */
128'h85a6842ac11dfda00413e47ff0ef84ae, /*   63 */
128'hcf63445c3f4050ef320505130000a517, /*   64 */
128'h5435102080ef31e505130000a51700f4, /*   65 */
128'h003085228082614564e2740270a28522, /*   66 */
128'h0d6080ef6522f565842adcfff0ef85a6, /*   67 */
128'h5479fcf71be30ff0079300c7c70367a2, /*   68 */
128'he50965a2de1ff0eff406e42e7179bfc1, /*   69 */
128'hf96dd97ff0ef08308082614570a24501, /*   70 */
128'he42eec064108842ae8221101bfc56562, /*   71 */
128'h852200030e6302053303c919db9ff0ef, /*   72 */
128'h60e2fda005138302610560e265a26442, /*   73 */
128'h0000b7977139bfdd4501808261056442, /*   74 */
128'h04130000b417f426f822639c4f478793, /*   75 */
128'h043b840d8c0564e484930000b4976564, /*   76 */
128'h892afc06e852ec4ef04a0280079302f4, /*   77 */
128'h942602f4043325ea0a130000aa1789ae, /*   78 */
128'h69e2790274a2744270e2450100849b63, /*   79 */
128'h2f0050ef855285ca6090808261216a42, /*   80 */
128'hbfc902848493c50171d060ef854a608c, /*   81 */
128'hb7e16522f569cdbff0ef852685ce0030, /*   82 */
128'h84b68432e42efc06f04af426f8227139, /*   83 */
128'hcb5ff0ef083065a2c115cf7ff0ef893a, /*   84 */
128'h70e2978285a2615c862686ca6562e519, /*   85 */
128'hbfc5fda0051380826121790274a27442, /*   86 */
128'h84b68432e42efc06f04af426f8227139, /*   87 */
128'hc75ff0ef083065a2c115cb7ff0ef893a, /*   88 */
128'h70e2978285a2655c862686ca6562e519, /*   89 */
128'hbfc5fda0051380826121790274a27442, /*   90 */
128'hc7dff0ef84b2e42ef822fc06f4267139, /*   91 */
128'h701ce509c39ff0ef842a083065a2c105, /*   92 */
128'h8082612174a2744270e2978285a66562, /*   93 */
128'h2785c3190017f713419cbfcdfda00513, /*   94 */
128'hd71b8e5927a106220086571b419cc19c, /*   95 */
128'h0ff77713c19c0087d7138ed906a20086, /*   96 */
128'h122300d5112300c510238fd90087979b, /*   97 */
128'hf022f4067179419c80820005132300f5, /*   98 */
128'h419c00f510230457879b6785c19c27d1, /*   99 */
128'h0087979b0ff777130087d713c632842a, /*  100 */
128'hc4360509084c57fd460900f11a238fd9, /*  101 */
128'h0513016105934609006070ef00f11b23, /*  102 */
128'h00041323082c462147c17f9060ef0044, /*  103 */
128'h00f404a347c57e5060efec3e00840513, /*  104 */
128'h7cf060ef00c4051300041523006c4611, /*  105 */
128'h014406937c3060ef01040513002c4611, /*  106 */
128'hfed79ce39f31ffe7d6030789470187a2, /*  107 */
128'h9fb94107d71b9fb9934117424107579b, /*  108 */
128'h80826145740270a200f41523fff7c793, /*  109 */
128'h97b6472167856394310787930000b797, /*  110 */
128'hc7bb27850077e793fff6079b8007bc23, /*  111 */
128'h678500f747630005071b6805450102e7, /*  112 */
128'h00e588b300351713808280c6b82396be, /*  113 */
128'hbfe1050501173023973697420008b883, /*  114 */
128'he406450185aa86220005841be0221141, /*  115 */
128'h717980820141640260a28522fa1ff0ef, /*  116 */
128'he436f4064619051984b2842aec26f022, /*  117 */
128'h6ff060ef85b64619852266a270b060ef, /*  118 */
128'h00e4859b70a27402852200f4162347a1, /*  119 */
128'h6785737dc5010113fadff06f614564e2, /*  120 */
128'h38913c233a113423392138233a813023, /*  121 */
128'h3761382337513c233941302339313423, /*  122 */
128'h35a1382335913c233781302337713423, /*  123 */
128'hd00007b7943e747d978a911a35078793, /*  124 */
128'hf0040023e0040023ca040b23ce042023, /*  125 */
128'h00e7ea63892a5800073797aad0040023, /*  126 */
128'ha001002050eff5e505130000a51785aa, /*  127 */
128'h871374fd678524f71d63478900054703, /*  128 */
128'h970a350787139abacd848a93970a3507, /*  129 */
128'h49818a368cb28baed0048c13cb848b13, /*  130 */
128'hcd03013907b395ca0f0985939c3a9b3a, /*  131 */
128'h89bb058902a0071329890f07c7830015, /*  132 */
128'h22e78f63471904f76b6326e78b6301a9, /*  133 */
128'hcc848513470d2ae78963470502f76263, /*  134 */
128'h40ef062505130000a51785be22e78763, /*  135 */
128'hfee794e3473d22e783634731bf4d77f0, /*  136 */
128'h953e866ae0048513978a350787936785, /*  137 */
128'h03600713b769e00d00235c9060ef9d22, /*  138 */
128'h20e78e630330071300f76e6322e78163, /*  139 */
128'haac94605cb648513fae798e303500713, /*  140 */
128'hf8e79ce30ff0071324e7856303800713, /*  141 */
128'h8363479924f58363747d479500614583, /*  142 */
128'h16079263000ca7833af59f63478938f5, /*  143 */
128'h0593ce4405134985978a350a87936a85, /*  144 */
128'h8793551060ef013ca023953e46110109, /*  145 */
128'h953e461101490593ce840513978a350a, /*  146 */
128'h54e25a52e3c505130000a51753b060ef, /*  147 */
128'hcf840913978a350a87936bb040efde02, /*  148 */
128'h03a3478d4c5060ef854a55fd4619993e, /*  149 */
128'h978a350a879346f115231350079300f1, /*  150 */
128'h46c1051385a6460594becb740493c2a6, /*  151 */
128'h879346f106a3032007934e9060efc0d2, /*  152 */
128'h051346114a1195becf040593978a350a, /*  153 */
128'h09a3036007934c5060ef4741072346f1, /*  154 */
128'h461195becf440593978a350a879346f1, /*  155 */
128'h460557fd4a3060ef47410a2347510513, /*  156 */
128'h0d23000103a346f10ca347b1051385a6, /*  157 */
128'h45810f00061310200793489060ef4731, /*  158 */
128'h1d2310100793427060efde3e37a10513, /*  159 */
128'h36f10e233961051385de4799464136f1, /*  160 */
128'h679946f113232637879377e145b060ef, /*  161 */
128'h0413978a350a879346f1142335378793, /*  162 */
128'h051385a20440061304300693943ecec4, /*  163 */
128'h35e1051385a2460156fdba5ff0ef3721, /*  164 */
128'hcf3ff0ef0e8885de86ca5672bd9ff0ef, /*  165 */
128'h398134833a0134033a813083911a6305, /*  166 */
128'h37813a8338013a033881398339013903, /*  167 */
128'h35813c8336013c0336813b8337013b03, /*  168 */
128'h4611cd04851380823b01011335013d03, /*  169 */
128'h87936785a00d953e978a350787936785, /*  170 */
128'h60ef9d22953e866af0048513978a3507, /*  171 */
128'h39f060ef85564611b3bdf00d00233ad0, /*  172 */
128'h978a350787936785bfdd855a4611b395, /*  173 */
128'hce045783383060ef4611953ece048513, /*  174 */
128'h578300f411238fd90087979b0087d71b, /*  175 */
128'h00f410238fd90087979b0087d71bce24, /*  176 */
128'h866ab749cc048513bb39cef42023401c, /*  177 */
128'h2783b321d00d0023347060ef9d228562, /*  178 */
128'h0000a51700fa2023478512079a63000a, /*  179 */
128'h0e880109059346114b9040efc4c50513, /*  180 */
128'hcb840513978a35048793648531b060ef, /*  181 */
128'h35314703303060ef014905934611953e, /*  182 */
128'h0000a517350145833511460335214683, /*  183 */
128'h00a1468335015783479040efc1c50513, /*  184 */
128'h352157830cf71e230000b71700914603, /*  185 */
128'h0000b717c1c505130000a51700814583, /*  186 */
128'h01b14703445040ef00b147030cf71323, /*  187 */
128'h0000a517018145830191460301a14683, /*  188 */
128'h0121468301314703429040efc1c50513, /*  189 */
128'hc20505130000a5170101458301114603, /*  190 */
128'h05130000a51755c20101578340d040ef, /*  191 */
128'hb7170121578306f713230000b717c2e5, /*  192 */
128'hf6bb02f5d63b03c0079304f71e230000, /*  193 */
128'h02f5d5bbe107879b678502f6763b02f5, /*  194 */
128'h95bee0040593978a350487933cd040ef, /*  195 */
128'h350487933b5040efc08505130000a517, /*  196 */
128'hc00505130000a51795be978af0040593, /*  197 */
128'h40efc0a505130000a517bbf539d040ef, /*  198 */
128'h20234785de0794e3000a2783b3fd38f0, /*  199 */
128'ha517373040efbfe505130000a51700fa, /*  200 */
128'h350787936785367040efc02505130000, /*  201 */
128'hc08505130000a51795be978ad0040593, /*  202 */
128'hb34d343040efc0e505130000a517bf45, /*  203 */
128'hf852fc4ee0cae4a6e8a2ec86711d737d, /*  204 */
128'h6a85c22505130000a517911a89aaf456, /*  205 */
128'h0493978a020a8793747d31b040efca02, /*  206 */
128'hb797123060ef852655fd461994beff84, /*  207 */
128'hc83e4a05fef40913439ccda787930000, /*  208 */
128'h993e978a020a879312f11d2313500793, /*  209 */
128'h0793141060ef014107a31a68460585ca, /*  210 */
128'h020a879312f10f23479112f10ea30370, /*  211 */
128'h60ef13f10513461195beff040593978a, /*  212 */
128'h14f101a314510513460585ca57fd11d0, /*  213 */
128'h0fc00793103060ef000107a315410223, /*  214 */
128'h0a1060efca3e04a1051345810f000613, /*  215 */
128'h05134641479985ce04f1152310100793, /*  216 */
128'h2637879377e10d5060ef04f106230661, /*  217 */
128'h879312f11c2335378793679912f11b23, /*  218 */
128'h06930421051385a2943e1451978a020a, /*  219 */
128'h02e1051385a2821ff0ef044006130430, /*  220 */
128'h85ce86a610084652855ff0ef460156fd, /*  221 */
128'h64a66446450160e6911a630596fff0ef, /*  222 */
128'ha51785aa808261257aa27a4279e26906, /*  223 */
128'hf0a2f48671591f70406fb12505130000, /*  224 */
128'h05a1051384aa81010113e4cee8caeca6, /*  225 */
128'h60efd602e83eec3ae442893689b2e046, /*  226 */
128'h6762747d97ba810787931018678503d0, /*  227 */
128'h0521051385a2864a86ba943e7fc40413, /*  228 */
128'h863e86c285a267c26822f94ff0efd64e, /*  229 */
128'h85a6180856326882fc4ff0ef03e10513, /*  230 */
128'h7406450170a67f0101138ddff0ef86c6, /*  231 */
128'he222e606716d8082616569a6694664e6, /*  232 */
128'h00254703003547830045480300554883, /*  233 */
128'h85930000a597842a0005460300154683, /*  234 */
128'h8522143040efa76505130000a517a765, /*  235 */
128'h85930000a597860ac10d842ae01ff0ef, /*  236 */
128'h8522123040efa7e505130000a517a565, /*  237 */
128'ha98505130000a51780826151641260b2, /*  238 */
128'h7159b7cd105040efd007a8230000b797, /*  239 */
128'hec66f062f45ef85afc56e0d2e4ceeca6, /*  240 */
128'h44818aae89aae46ee8caf0a2f486e86a, /*  241 */
128'ha70b0b130000ab177a0a0a130000aa17, /*  242 */
128'h0000ac97a7cc0c130000ac1706000b93, /*  243 */
128'h035441630004841bfff58d1ba6cc8c93, /*  244 */
128'h7b427ae26a0669a6694664e6740670a6, /*  245 */
128'hc01d808261656da26d426ce27c027ba2, /*  246 */
128'hff048913085040ef855ae39d00f47793, /*  247 */
128'h588505130000a51702879d630009079b, /*  248 */
128'hc583009987b3067040ef855206d040ef, /*  249 */
128'h1263053040efa16505130000a5170007, /*  250 */
128'h87b3a80500f979134d81fffd4913068d, /*  251 */
128'he7630ff7f793fe05879b0007c5830129, /*  252 */
128'h40ef8562b75d0905029040ef856600fb, /*  253 */
128'hff2dcce32d85017040ef8552bfdd01f0, /*  254 */
128'h079b4124093b007040ef00f4f913855a, /*  255 */
128'h40ef50a505130000a51700f45a630009, /*  256 */
128'h879b0007c583012987b3bf1504857ee0, /*  257 */
128'h7d0040ef856600fbe7630ff7f793fe05, /*  258 */
128'hec267179bfdd7c6040ef8562b7f10905, /*  259 */
128'ha697893289ae84b6f022f406e44ee84a, /*  260 */
128'h968686930000a697c509222686930000, /*  261 */
128'h960606130000a617e187071300009717, /*  262 */
128'h5d6300098f63842a748040ef854a85a6, /*  263 */
128'h948606130000a61786ce40a485bb0095, /*  264 */
128'h00f44463ffe4879b9c2972a040ef954a, /*  265 */
128'h918585930000a59700890533ffd4841b, /*  266 */
128'h69a2694264e2854a740270a2306060ef, /*  267 */
128'h7115f73ff06f4581862e86b280826145, /*  268 */
128'h002cfebff0efed8645050c800613002c, /*  269 */
128'h450160ee714040ef900505130000a517, /*  270 */
128'h6963862e9ff787133b9ad7b78082612d, /*  271 */
128'h079304a7676323f78713000f47b704a7, /*  272 */
128'h0000b7173e80079346890ca7fc633e70, /*  273 */
128'hec0600074903e04a973611018cc70713, /*  274 */
128'h690264a260e2644202091663e426e822, /*  275 */
128'h6b00406f61058a6505130000a51785aa, /*  276 */
128'hbf7d240787934685b7d9a00787934681, /*  277 */
128'h47293e800793c81502f555b302f57433, /*  278 */
128'h0713cf3902f4773346a547a90687e263, /*  279 */
128'h743302f457b30640071300877d630630, /*  280 */
128'h0000a517943e001444130324341302e4, /*  281 */
128'ha51785a2c801656040ef84b285c50513, /*  282 */
128'h862660e26442646040ef852505130000, /*  283 */
128'h6105842505130000a517690264a285ca, /*  284 */
128'hf46302f45733bf6102e4543362c0406f, /*  285 */
128'h0000951785aabf554401bf51843a0086, /*  286 */
128'h86bb459958d94701862ebfa17fc50513, /*  287 */
128'h1702cf8500f557b3883e03c6879b02e8, /*  288 */
128'he426972e11017ce585930000a5979301, /*  289 */
128'h60e26442e495e04ae822ec0600074483, /*  290 */
128'h61057da505130000951785aa690264a2, /*  291 */
128'h0000951785aafab71ce327055bc0406f, /*  292 */
128'hfff7471301071733577db7f57c450513, /*  293 */
128'h03b6869b02e505334729c10d44018d79, /*  294 */
128'h746301045433942a472500d414334405, /*  295 */
128'h770505130000951785be078514590087, /*  296 */
128'h05130000951785a2c80156a040ef8932, /*  297 */
128'h690285a6864a60e2644255a040ef7665, /*  298 */
128'h5400406f610576e505130000951764a2, /*  299 */
128'hf54ef94ae1a202c7073b8cbafce67155, /*  300 */
128'he162e55ee95aed56f152fd26e586f8ea, /*  301 */
128'hf66384368d3289ae892a04000793f4ee, /*  302 */
128'h4cc1000c956302ccdcbb04000c9300e7, /*  303 */
128'h001a849b020d1a13001d1a9b03acdcbb, /*  304 */
128'h00009b9771cb0b1300009b17020a5a13, /*  305 */
128'h4501e00d5dcc0c1300008c17684b8b93, /*  306 */
128'h6b4a6aea7a0a79aa794a74ea640e60ae, /*  307 */
128'h85ca808261697da67d467ce66c0a6baa, /*  308 */
128'h00040d9b4a4040ef6d85051300009517, /*  309 */
128'h482146914781874e000c8d9b008cf463, /*  310 */
128'h9381020d979305b66b630007861b4889, /*  311 */
128'h083803bd06bb0d9de56399be034787b3, /*  312 */
128'h0b079c630006881b02e0089385ba4781, /*  313 */
128'h8c23e036694505130000951797ba1098, /*  314 */
128'h9281168241b4043b668244a040effa07, /*  315 */
128'h02dd1963b79d557dd13d0b0070ef9936, /*  316 */
128'h1602c19095aa26010828002795934310, /*  317 */
128'h6702412040efe03ae43e855a85d69201, /*  318 */
128'h1963bf9d4691482107859752488967a2, /*  319 */
128'hbfd1e19095aa0828003795936310010d, /*  320 */
128'h164208280017959300075603011d1d63, /*  321 */
128'h082c00074603bf6d00c5902395aa9241, /*  322 */
128'he03e855eb76500c580230ff6761395be, /*  323 */
128'hbf253cfdfe97eae3278567820dc070ef, /*  324 */
128'h0005450300cc053300074603bfdd4781, /*  325 */
128'h54634186561b0186161bc51909757513, /*  326 */
128'h87aa1582b70d07052785011700230006, /*  327 */
128'h8f8d25058082e21c00b7f46345019181, /*  328 */
128'h47370005668312b7f46304000793bfd5, /*  329 */
128'h0045468310e69c63478957f70713464c, /*  330 */
128'h7159038007930385570310e697634709, /*  331 */
128'hf48602059a93fc567100f0a202f70733, /*  332 */
128'hec66f062f45ef85ae0d2e4cee8caeca6, /*  333 */
128'h06eae663478d9722020ada93e46ee86a, /*  334 */
128'h8b9300009b974b054a01942a84aa892e, /*  335 */
128'h8c9300009c97586c0c1300009c17546b, /*  336 */
128'h401ca835478100fa64630384d783566c, /*  337 */
128'h2d0040ef855e85d2cbc1741c09679b63, /*  338 */
128'h8db301843d03640c04098d6302043983, /*  339 */
128'h051300009517864a02bafa6395ce00b4, /*  340 */
128'h694664e6740670a6478d2aa040ef5065, /*  341 */
128'h6d426ce27c027ba27b427ae26a0669a6, /*  342 */
128'h856686ce85ea866e80826165853e6da2, /*  343 */
128'h39830e0060ef856a85ee864e27c040ef, /*  344 */
128'h40f989b301843d030337f163701c0284, /*  345 */
128'h4581864e254040ef856285ea9d3e864e, /*  346 */
128'h4785bf99038404132a0506a060ef856a, /*  347 */
128'h8082400005378082057e45058082853e, /*  348 */
128'h00756513157d631c658707130000a717, /*  349 */
128'h450597aa20000537e308953600178693, /*  350 */
128'h0ce507638207871367858082953e057e, /*  351 */
128'h0513000095178087871308a74463862a, /*  352 */
128'h95178006079b04c7496306e60b634a65, /*  353 */
128'h951787f787936785c3ad482505130000, /*  354 */
128'h7c07879b77fd04c7c963502505130000, /*  355 */
128'h0000a5174f458593000095979e3d1141, /*  356 */
128'h0000a51760a2182040efe4065bc50513, /*  357 */
128'h0000951781078713808201415ac50513, /*  358 */
128'h000095178187879300e60a6345450513, /*  359 */
128'h9517830787138082faf612e345450513, /*  360 */
128'h879300c74963fee609e3472505130000, /*  361 */
128'h83878713bfe944e50513000095178287, /*  362 */
128'h84078793fce608e34605051300009517, /*  363 */
128'h051300009517bf754605051300009517, /*  364 */
128'h84aaf406e84aec26f022717980824165, /*  365 */
128'h551302f04463409907bb00a5893b4401, /*  366 */
128'h70a2952201045513942a904114420104, /*  367 */
128'h61459141694264e21542fff545137402, /*  368 */
128'h00c15783753050ef0068460985a68082, /*  369 */
128'h00f117238fd90087979b0087d71b0489, /*  370 */
128'he486e0a26785715dbf45943e93c117c2, /*  371 */
128'h3cf50463842e80678793f44ef84afc26, /*  372 */
128'h99638005079b0af50e636dd7879367a1, /*  373 */
128'h0913701050ef4611082884b205e94407, /*  374 */
128'h50ef4aa505130000a517461985ca0064, /*  375 */
128'he76332f5886302e00793017445836ed0, /*  376 */
128'h8263479104b7e5631cf5816347b108b7, /*  377 */
128'h9517478910f58463478502b7e3631af5, /*  378 */
128'h05130000951702f5836339a505130000, /*  379 */
128'h47a118f581634799a41503a040ef5365, /*  380 */
128'h020040effef591e33a05051300009517, /*  381 */
128'h896347c500b7ed632cf5816347f5a429, /*  382 */
128'hfef580e33bc505130000951747d916f5, /*  383 */
128'h96e3029007932af5856302100793bf6d, /*  384 */
128'h06200793b7c93d65051300009517faf5, /*  385 */
128'h2af581630330079304b7e2632cf58163, /*  386 */
128'h0320079328f5866302f0079300b7ef63, /*  387 */
128'h0793b7bdf8f58ae33d85051300009517, /*  388 */
128'h05130000951705e0079328f5836305c0, /*  389 */
128'h28f5856308400793bf91f6f58de33ee5, /*  390 */
128'h06c0079326f58a630670079300b7ef63, /*  391 */
128'h0793b73df4f58ae34005051300009517, /*  392 */
128'h079326f588630ff0079326f587630890, /*  393 */
128'hb73d40a5051300009517f0f59ce30880, /*  394 */
128'h0000a9973bc7d7830000a79701e45703, /*  395 */
128'h0000a7970204570312f713633b498993, /*  396 */
128'h50ef852285ca461910f71b633a67d783, /*  397 */
128'h50ef854a374585930000a597461958d0, /*  398 */
128'h1f23020412230204012301a4578357d0, /*  399 */
128'h102302240513fde4859b01c4578300f4, /*  400 */
128'h1e230029d78300f41d230009d78302f4, /*  401 */
128'h1e238d5d05220085579bdb3ff0ef00f4, /*  402 */
128'hda5fe0ef450185a2862602a4122300a1, /*  403 */
128'h00009517bd4920e5051300009517a06d, /*  404 */
128'hbdbd22a5051300009517b56121c50513, /*  405 */
128'h0254478300f10ea30264470302444783, /*  406 */
128'h0274470300e10ea301c1178300f10e23, /*  407 */
128'h0ea301c119030224470300e10e232781, /*  408 */
128'h56830450071300e10e230234470300e1, /*  409 */
128'h47e228d79b230000a79704e79b6301c1, /*  410 */
128'h05130000a51726e585930000a5974619, /*  411 */
128'h49f050efe43626f72b230000a7172765, /*  412 */
128'hff89061b24c787930000a79766a24762, /*  413 */
128'h74e2640660a6590060ef450102a40593, /*  414 */
128'h04e69463043007138082616179a27942, /*  415 */
128'h87930000a79722f72b230000a71747e2, /*  416 */
128'h439c22a787930000a797c799439c23a7, /*  417 */
128'h06130000a61721e686930000a697f7e9, /*  418 */
128'he0ef02a4051321e585930000a59721a6, /*  419 */
128'h0000951702e798634d200713b765d4bf, /*  420 */
128'hca2ff0ef852285a65a9030ef14450513, /*  421 */
128'h051385ca595030ef1405051300009517, /*  422 */
128'hf6e787e35fe00713bf95c8cff0ef02a4, /*  423 */
128'h02045703f6f701e317fd67c101e45703, /*  424 */
128'h08681da585930000a5974611f4f70de3, /*  425 */
128'hb33d11a5051300009517b7993cb050ef, /*  426 */
128'h051300009517b3151205051300009517, /*  427 */
128'h9517bb011445051300009517bb291365, /*  428 */
128'h1605051300009517b31915a505130000, /*  429 */
128'h00009517b9cd17e5051300009517b9f5, /*  430 */
128'hb9f91a25051300009517b1e518c50513, /*  431 */
128'h051300009517b9d11c85051300009517, /*  432 */
128'h1587d7830000a7970265d703b1e91d65, /*  433 */
128'h0285d703ecf711e3150484930000a497, /*  434 */
128'h20000793eaf719e31427d7830000a797, /*  435 */
128'h85ce461900f59a230165899302058913, /*  436 */
128'h100585930000a5974619319050ef854a, /*  437 */
128'h0f0585930000a5974619309050ef854e, /*  438 */
128'h50ef852285ca46192f7050ef00640513, /*  439 */
128'h578302f4132302a0061301c457832ed0, /*  440 */
128'hd78300f41e230004d78302f4142301e4, /*  441 */
128'hb36900f416236080079300f41f230024, /*  442 */
128'h4601443030ef15e505130000951785aa, /*  443 */
128'h30239f0101138307b603300017b7bba5, /*  444 */
128'h179b66858387b70300f6741326016081, /*  445 */
128'h300005b79fad8406879b0387f5930034, /*  446 */
128'h881b2781601134235e913c23639c97ae, /*  447 */
128'h8a1d09056c63ffc7849b5f200513fee7, /*  448 */
128'h27018f71fff7471300c5163b10100513, /*  449 */
128'h171beb3d4318026707130000a717c349, /*  450 */
128'h95ba070e9f318006871b700776130084, /*  451 */
128'hd69b0106d69b0106969b00d100a345d4, /*  452 */
128'hc6918005069b0001550300d100230086, /*  453 */
128'h0077e79337ed02d51e63806686936685, /*  454 */
128'h85b246814037d79b30000837860a2785, /*  455 */
128'h0621068500083803983a003698139742, /*  456 */
128'hf0ef8626fef845e30006881bff063c23, /*  457 */
128'h608130838287b823300017b70405a9bf, /*  458 */
128'h8082610101135f813483852660013403, /*  459 */
128'h2401ec06e42643c0e8220c2007b71101, /*  460 */
128'hc163033716938304b703300014b74781, /*  461 */
128'h311030ef0445051300009517e7990206, /*  462 */
128'h8082610564a2644260e2c3c00c2007b7, /*  463 */
128'h8432ec26f0227179bfc14785ec3ff0ef, /*  464 */
128'hf4060068f5c585930000a597461184ae, /*  465 */
128'h0007a803f14787930000a79714b050ef, /*  466 */
128'ha717efa888930000a89785a6862247b2, /*  467 */
128'h05130000a51704500693efe757030000, /*  468 */
128'h614564e2740270a285228b8ff0eff065, /*  469 */
128'h8082914115428d5d05220085579b8082, /*  470 */
128'hf00686938fd966c10185579b0185171b, /*  471 */
128'h00ff07370085151b8fd98f750085571b, /*  472 */
128'h879b070007b7715d808225018d5d8d79, /*  473 */
128'he0a2e48604b005134585460100740207, /*  474 */
128'h017070efc63eec56f052f44ef84afc26, /*  475 */
128'h4401233030eff7e50513000095178a2a, /*  476 */
128'h091300009917e7e989930000a9975ae1, /*  477 */
128'h0004059b013407b3028a863b4499f769, /*  478 */
128'h0ff6761300ca56330286061b0405854a, /*  479 */
128'ha5974611fc941ee31f9030ef00c78023, /*  480 */
128'ha5974609053050ef0048e44585930000, /*  481 */
128'hf0ef4512043050ef0028e32585930000, /*  482 */
128'h0087179bf0060613010006374722f43f, /*  483 */
128'h300016b78fd915020ff777138ff18321, /*  484 */
128'hb78380f6b42393c180a6b02317c29101, /*  485 */
128'h82f6b42347a1640660a68086b7838006, /*  486 */
128'h17b7808261616ae27a0279a2794274e2, /*  487 */
128'h0080073771398087b5838007b6033000, /*  488 */
128'hec4ef04af426f822fc068f4d91c115c2, /*  489 */
128'h05130000951780e7b423e05ae456e852, /*  490 */
128'ha797d9d747030000a71714b030efebe5, /*  491 */
128'ha697d8f848030000a817d967c7830000, /*  492 */
128'ha597d7b646030000a617d846c6830000, /*  493 */
128'h30efe925051300009517d725c5830000, /*  494 */
128'h448100044783d5e404130000a41710f0, /*  495 */
128'hd4f708230000a717d38989930000a997, /*  496 */
128'ha7176a89d2ca0a130000aa1700144783, /*  497 */
128'h193700262b3700244783d2f70da30000, /*  498 */
128'ha71700344783d2f704230000a7173000, /*  499 */
128'h09230000a71700444783d0f70ea30000, /*  500 */
128'ha797d0f703a30000a71700544783d0f7, /*  501 */
128'ha797cc07a9230000a797cc079f230000, /*  502 */
128'ha797cc07a7230000a797cc07ad230000, /*  503 */
128'h8522e78d0009a783e4a9cc07a1230000, /*  504 */
128'h03379713830937835a0b0493efbfe0ef, /*  505 */
128'hfc075de3033797138309378302074563, /*  506 */
128'h4501dff154fd000a2783bfc5c13ff0ef, /*  507 */
128'hb7e9bf9ff0efbfc1710a849300a060ef, /*  508 */
128'hff8006b78087b703300017b7b7d914fd, /*  509 */
128'h0713670580e7b4238f75e40616fd1141, /*  510 */
128'h0513000095178307b58382e7b823f007, /*  511 */
128'h30efdca50513000095177fa030efdae5, /*  512 */
128'h90738fd9880707136709300027f37ee0, /*  513 */
128'h0513000095173417907307fe47853007, /*  514 */
128'h00730ff0000f0000100f7ca030efdc65, /*  515 */
128'h00054703001547838082014160a23020, /*  516 */
128'h8fd907c200354503002547838f5d07a2, /*  517 */
128'h13630007871b4781808225018d5d0562, /*  518 */
128'h00f507330007468300f58733808200e6, /*  519 */
128'h13630005079b9e29b7d500d700230785, /*  520 */
128'h1101495cbfc5feb50fa30505808200f6, /*  521 */
128'h3903cfb500958413e04ae426ec06e822, /*  522 */
128'h02e00893482145150200061347810185, /*  523 */
128'h146302c700630007470300f9073346ad, /*  524 */
128'h0023010315630007831b0e50071300a7, /*  525 */
128'hfcd79be30785040500e4002304050114, /*  526 */
128'hf0ef00f5842384ae01c9051300b94783, /*  527 */
128'h0087979b0189470301994783c088f4bf, /*  528 */
128'h979b016947030179478300f492238fd9, /*  529 */
128'h644260e20004002300f493238fd90087, /*  530 */
128'h0593cf99873e611c80826105690264a2, /*  531 */
128'h986302d5fc630007468303a006130200, /*  532 */
128'h0705a00d577d00d706630017869300c6, /*  533 */
128'hf593fd06869b577d46050007c683b7dd, /*  534 */
128'h853ae11c0006871b078900b666630ff6, /*  535 */
128'h611cc915bfd5b06747030000a7178082, /*  536 */
128'h008557030067d683c70d0007c703cb85, /*  537 */
128'h35e060ef0017c503e406114102e69063, /*  538 */
128'h8082014160a24525c391450100157793, /*  539 */
128'h979b470d01a5c68301b5c78380824525, /*  540 */
128'h0155c70300e51d630006879b8edd0087, /*  541 */
128'h8fd50107979b8fd10087179b0145c603, /*  542 */
128'h5904e44eec26f02271798082853e2781, /*  543 */
128'h00154503842a03450993e052e84af406, /*  544 */
128'h505ce13125012ec060ef85ce86264685, /*  545 */
128'h450100e7eb6340f487bb000402234c58, /*  546 */
128'h808261456a0269a2694264e2740270a2, /*  547 */
128'h001445034c5cff2a74e34a0500344903, /*  548 */
128'hb7e5397d2aa060ef85ce86269cbd4685, /*  549 */
128'h4501f8dff06fc39900454783b7f94505, /*  550 */
128'h4401e04ae426ec06e8221101591c8082, /*  551 */
128'h0005041bfddff0ef892e84aa02b78763, /*  552 */
128'h60ef03448593864a46850014c503ec19, /*  553 */
128'h85220324a823597d4405c11925012320, /*  554 */
128'he822110180826105690264a2644260e2, /*  555 */
128'h842ad91c0005022357fde04ae426ec06, /*  556 */
128'h2324470323344783e52d2501fa3ff0ef, /*  557 */
128'hd79b776d0107979b8fd90087979b4509, /*  558 */
128'hf0ef06a4051302e79f63a55707134107, /*  559 */
128'h4537fff50913010005370005079bd4bf, /*  560 */
128'h00978c6345010127f7b3146504930054, /*  561 */
128'h8d05012575332501d25ff0ef08640513, /*  562 */
128'h80826105690264a2644260e200a03533, /*  563 */
128'hfc26e0a2e486f44ef84a715dbfcd450d, /*  564 */
128'hf0ef8932852e89aa00053023ec56f052, /*  565 */
128'h0000a7970035171302054e6347adddbf, /*  566 */
128'hb023c01547b184aa638097ba90c78793, /*  567 */
128'h17e060ef00144503c79d000447830089, /*  568 */
128'h47a9c111891100090563e38500157793, /*  569 */
128'h853e6ae27a0279a2794274e2640660a6, /*  570 */
128'h00a400a3000400230ff4f51380826161, /*  571 */
128'h00090463fb79478d00157713092060ef, /*  572 */
128'h1a634785ee5ff0ef85224581f5718911, /*  573 */
128'h478389a623a40a131fa40913848a04f5, /*  574 */
128'ha0232501c51ff0ef854ac7894501ffc9, /*  575 */
128'haa0301048913ff2a14e30991094100a9, /*  576 */
128'hea1ff0ef852285d2000a076345090004, /*  577 */
128'h00e519634785470dfe9915e30491c10d, /*  578 */
128'h47b5c1194a01f6e505e34785470dbf85, /*  579 */
128'h8fd90087979b03f4470304044783b785, /*  580 */
128'hfee791e3200007134107d79b0107979b, /*  581 */
128'h00f9e9b30089999b04a4478304b44983, /*  582 */
128'h470501342e230444448329811a098763, /*  583 */
128'hfaf769e30ff7f793009401a3fff4879b, /*  584 */
128'h079b2901fa0903e30124012304144903, /*  585 */
128'h0454478304644a83ffc100f977b3fff9, /*  586 */
128'h00faf7930154142300faeab3008a9a9b, /*  587 */
128'h8d5d0085151b0474478304844503ffbd, /*  588 */
128'h979b2501042447030434478314050e63, /*  589 */
128'h004ad71b2781033486bbdfa98fd90087, /*  590 */
128'h40c5063bf4c563e3873200d7063b9f3d, /*  591 */
128'h490516556605f3266ce384ae032655bb, /*  592 */
128'h073b090900b939331955694100b67763, /*  593 */
128'h03442023cc04d458014787bb24890147, /*  594 */
128'h06040513f00a93e310e91163470dd05c, /*  595 */
128'hd49b1ff4849b0024949bd408b09ff0ef, /*  596 */
128'hf8000793c45cc81c57fdee99e6e30094, /*  597 */
128'h47030654478308f91963478d00f402a3, /*  598 */
128'h4107d79b0107979b8fd90087979b0644, /*  599 */
128'hce7ff0ef8522001a059b06e79b634705, /*  600 */
128'h000402a32324470323344783e13d2501, /*  601 */
128'h4107d79b776d0107979b8fd90087979b, /*  602 */
128'ha8dff0ef0344051304e79263a5570713, /*  603 */
128'h051302f51763252787932501416157b7, /*  604 */
128'h272787932501614177b7a77ff0ef2184, /*  605 */
128'h0513c808a61ff0ef21c4051300f51c63, /*  606 */
128'h6927d78300009797c448a57ff0ef2204, /*  607 */
128'h132368f712230000971793c117c22785, /*  608 */
128'h0513b351478100042a230124002300f4, /*  609 */
128'h05440513b5b10005099ba27ff0ef0584, /*  610 */
128'h4789d41c9fb5e00a84e3b545a19ff0ef, /*  611 */
128'h029787bb478db7090014949b00f91563, /*  612 */
128'hec06e8221101bdcd9cbd0017d79b8885, /*  613 */
128'h00044703ed692501c01ff0ef842ae426, /*  614 */
128'h0af71b634785005447030cf71063478d, /*  615 */
128'h9fdff0ef852645812000061303440493, /*  616 */
128'h22f409a3faa0079322f4092305500793, /*  617 */
128'h0610079302f40aa302f40a2305200793, /*  618 */
128'h0ba304100713481c20f40da302f40b23, /*  619 */
128'h571b0107571b0107971b20e40d2302e4, /*  620 */
128'hd79b0107d71b20e40ea320f40e230087, /*  621 */
128'h971b501020e40f23445c20f40fa30187, /*  622 */
128'h0693001445030087571b0107571b0107, /*  623 */
128'h0107d71b260522e400a322f400230720, /*  624 */
128'h22e4012320d40ca320d40c230187d79b, /*  625 */
128'h02a35d9050ef85a64685d81022f401a3, /*  626 */
128'h25015cd050ef45814601001445030004, /*  627 */
128'h4d188082610564a2644260e200a03533, /*  628 */
128'h0025478300e7f963377985beffe5879b, /*  629 */
128'h47858082450180829d3d02b787bb5548, /*  630 */
128'hec26f022f406e84a71794d180eb7f563, /*  631 */
128'h842e46890005470302e5f963892ae44e, /*  632 */
128'hd49b00f71e6308d70d63468d06d70b63, /*  633 */
128'hac7ff0ef9dbd0094d59b9cad515c0015, /*  634 */
128'h69a2694264e2740270a257fdc9112501, /*  635 */
128'hd59b0014899b0249278380826145853e, /*  636 */
128'h0344c483854a9dbd94ca1ff4f4930099, /*  637 */
128'h4783994e1ff9f993f5792501a93ff0ef, /*  638 */
128'hbf658391c0198fc50087979b88050349, /*  639 */
128'hf0ef9dbd0085d59b515cbf4d93d117d2, /*  640 */
128'h99221fe474130014141bf1452501a65f, /*  641 */
128'hb7618fc90087979b0349450303594783, /*  642 */
128'hf93d2501a3bff0ef9dbd0075d59b515c, /*  643 */
128'hf0ef954a034505131fc575130024151b, /*  644 */
128'h8082853e4785bfb9024557931512ffaf, /*  645 */
128'he852ec4ef822fc06f04a4544f4267139, /*  646 */
128'h450900f49c63892a478500b51523e456, /*  647 */
128'h61216aa26a4269e2790274a2744270e2, /*  648 */
128'hc683e0a9842efee4f4e34f98611c8082, /*  649 */
128'h0087d703eb0d579800e69463470d0007, /*  650 */
128'h0044579bd171009928235788fce477e3, /*  651 */
128'h87930416883d0009378300f92a239fa9, /*  652 */
128'hc98384bab75d450100893c23943e0347, /*  653 */
128'h766385a60009350309924a855a7d0027, /*  654 */
128'h049be75ff0efbf7d2501e5dff0ef0134, /*  655 */
128'h4f9c00093783f69afce301448c630005, /*  656 */
128'h5583b7954505bfc14134043bf6f4f7e3, /*  657 */
128'hf35ff0ef842aec06e426e822110100a5, /*  658 */
128'h049b939ff0ef6008484ce4950005049b, /*  659 */
128'hf3cff0ef4581020006136c08ec990005, /*  660 */
128'h00e782234705601c00e7802357156c1c, /*  661 */
128'hec4e71398082610564a28526644260e2, /*  662 */
128'h4a094985e456f04af426f822fc06e852, /*  663 */
128'h47830af5f0634a0984aa4d1c0ab9f563, /*  664 */
128'h8863470d0ae78f63842e893247090005, /*  665 */
128'h00b989bb515c0015d99b093794630ee7, /*  666 */
128'h166300050a1b8bdff0ef9dbd0099d59b, /*  667 */
128'h1ff9f9930ff9779300198a9b8805060a, /*  668 */
128'hf71316c166850347c783013487b3cc19, /*  669 */
128'h99a60ff7f7938fd98ff50049179b00f7, /*  670 */
128'h009ad59b50dc00f48223478502f98a23, /*  671 */
128'h000a1f6300050a1b86fff0ef9dbd8526, /*  672 */
128'h9aa60ff979130049591bc40d1ffafa93, /*  673 */
128'h8552744270e200f482234785032a8a23, /*  674 */
128'h87b3808261216aa26a4269e2790274a2, /*  675 */
128'h9bc100f979130089591b0347c7830154, /*  676 */
128'hf0ef9dbd0085d59b515cb7e90127e933, /*  677 */
128'h74130014141bfc0a12e300050a1b815f, /*  678 */
128'h0109591b0109191b03240a2394261fe4, /*  679 */
128'h515cbf790134822303240aa30089591b, /*  680 */
128'h16e300050a1bfdcff0ef9dbd0075d59b, /*  681 */
128'h9aa603440a931fc474130024141bf80a, /*  682 */
128'h69338d71f00006372501d96ff0ef8556, /*  683 */
128'h0a230107d79b94260109179b29010125, /*  684 */
128'h591b0109579b00fa80a30087d79b0324, /*  685 */
128'hf4267139bf79012a81a300fa81230189, /*  686 */
128'h89ae84aae456e852f04af822fc06ec4e, /*  687 */
128'h02f96d634d1c0009056300c52903e991, /*  688 */
128'hed6347850005041bc5bff0efa8154905, /*  689 */
128'h69e2790274a2744270e2852244050087, /*  690 */
128'h4c9c08f4026357fd808261216aa26a42, /*  691 */
128'h24054c9c5afd4a05844afef461e3894e, /*  692 */
128'h85a24409b7e94401012a646300f46763, /*  693 */
128'h0ae305550a63c9012501c0dff0ef8526, /*  694 */
128'h85a2167d10000637b7cdfd241de3fb45, /*  695 */
128'h489c02099063e9052501debff0ef8526, /*  696 */
128'h0054c783c89c37fdf8e788e3577dc4c0, /*  697 */
128'h852685ce8622bfb500f482a30017e793, /*  698 */
128'h547df6f514e34785dd612501dbdff0ef, /*  699 */
128'h2905f822fc0600a55903f04a7139b795, /*  700 */
128'heb9993c1e456e852ec4ef42603091793, /*  701 */
128'h6aa26a4269e2790274a2744270e24511, /*  702 */
128'h842a8a2e00f97993d7ed495c80826121, /*  703 */
128'h5783e18dc85c61082785480c00099d63, /*  704 */
128'h15230996601cfcf775e30009071b0085, /*  705 */
128'h4783bf5d4501ec1c97ce034787930124, /*  706 */
128'hfc0a9fe30157fab337fd00495a9b0025, /*  707 */
128'h45090097e46347850005049bb2fff0ef, /*  708 */
128'h4d1c6008b761450500f4946357fdbf49, /*  709 */
128'h049be83ff0ef480cf60a0ee306f4e063, /*  710 */
128'h8de357fdfcf48be34785d4bd451d0005, /*  711 */
128'h06136008f5792501de0ff0ef6008fcf4, /*  712 */
128'h00043a03bf0ff0ef0345051345812000, /*  713 */
128'h60084a0502aa2823aabff0ef855285a6, /*  714 */
128'hd91c415787bb591c00faed6300254783, /*  715 */
128'h0223b7b9c848a89ff0ef85a6c8046008, /*  716 */
128'h5b1c2a856018f1412501d24ff0ef0145, /*  717 */
128'hf04afc06f426f8227139b7e9db1c2785, /*  718 */
128'h02f007130005c783e05ae456e852ec4e, /*  719 */
128'h0ce7946305c0071300e78663842e84aa, /*  720 */
128'h0ce7f06347fd000447030004a6230405, /*  721 */
128'h47834b2102e0099305c00a9302f00a13, /*  722 */
128'h462d0204b9030d5784630d4786630004, /*  723 */
128'h966300044783b42ff0ef854a02000593, /*  724 */
128'h07930b37946300144783013900230d37, /*  725 */
128'h470d1d3789630024478300f900a302e0, /*  726 */
128'h458100f905a302000793943a09479b63, /*  727 */
128'h48cc492d100519632501adfff0ef8526, /*  728 */
128'h47836c98100511632501ce0ff0ef6088, /*  729 */
128'h708cef898ba100b74783120780630007, /*  730 */
128'h46030006c68300f58633078500f706b3, /*  731 */
128'h2501df9ff0ef852645810cd60a63fff6, /*  732 */
128'h85264581bf35c55c4bdc611ca0e1dd5d, /*  733 */
128'h74a2744270e20004bc232501a81ff0ef, /*  734 */
128'h0405808261216b026aa26a4269e27902, /*  735 */
128'he76302000693f75787e3b7b54709b73d, /*  736 */
128'h45a147014681b78d02400793943a12f6, /*  737 */
128'he793a2110505a8c948e5020003134781, /*  738 */
128'h268500e50023954a9101020695130027, /*  739 */
128'h7363461194320200051392011602a865, /*  740 */
128'h95630e50071300094683c6e5460100e5, /*  741 */
128'h0027979b01659f6300e90023471500e6, /*  742 */
128'h0086661300e7946347118bb10ff7f793, /*  743 */
128'hfed714e346850037f713bded00c905a3, /*  744 */
128'h00b7c783709cf1279de3b7c501066613, /*  745 */
128'h0207f7930047f713f4e513e34711c515, /*  746 */
128'h4501e6070ae30004bc230004a623cb99, /*  747 */
128'hfbe58b91b7054515f315bfd94511b72d, /*  748 */
128'h0007c503609cdbe58bc100b5c7836c8c, /*  749 */
128'h0027979b05659a63b5a1c4c8ae4ff0ef, /*  750 */
128'h17020017061b873245ad46a10ff7f793, /*  751 */
128'hf3470be3f2e37de30007470397229301, /*  752 */
128'h0187151b02b6f263fd370ae3f35709e3, /*  753 */
128'hee0505130000851700054c634185551b, /*  754 */
128'hb5754519ef0719e30008066300054803, /*  755 */
128'hf9f7051beea8f3e30ff57513fbf7051b, /*  756 */
128'h77130017e7933701eca8efe30ff57513, /*  757 */
128'h842ae44ee84aec26f0227179bdc10ff7, /*  758 */
128'he199484c49bd0e500913451184aef406, /*  759 */
128'h6c1ce1292501aecff0ef6008a0b1c90d, /*  760 */
128'h026303f7f79300b7c783c3210007c703, /*  761 */
128'h9a630017b79317e18bfd033780630327, /*  762 */
128'h614569a2694264e2740270a245010097, /*  763 */
128'h2a23d9452501bfdff0ef852245818082, /*  764 */
128'hec06e82245811101bfe54511b7cd0004, /*  765 */
128'h0e500493e50d250187dff0ef842ae426, /*  766 */
128'hc7836c1ced092501a7eff0ef6008484c, /*  767 */
128'hbb7ff0ef85224585cb9900978d630007, /*  768 */
128'h644260e2451d00f513634791dd792501, /*  769 */
128'h842aec06e426e82211018082610564a2, /*  770 */
128'hf0ef6008484ce49d0005049bfa9ff0ef, /*  771 */
128'h4581020006136c08e0850005049ba34f, /*  772 */
128'h601c80eff0ef462d6c08700c838ff0ef, /*  773 */
128'h610564a28526644260e200e782234705, /*  774 */
128'he84af02271794d1c08b7f06347858082, /*  775 */
128'h06f5f063892e842ae052e44eec26f406, /*  776 */
128'h0005049bed6ff0ef852285ca59fd4a05, /*  777 */
128'h6a0269a2694264e2740270a24501e891, /*  778 */
128'h85ca460103348c6303448c6380826145, /*  779 */
128'h01378a63481cfd7125018abff0ef8522, /*  780 */
128'h00f402a30017e79300544783c81c2785, /*  781 */
128'hbf5d4509bf65faf4e7e30004891b4c1c, /*  782 */
128'hfc061028ec2a713980824509bf4d4505, /*  783 */
128'h979704054263832ff0eff42ee432e82e, /*  784 */
128'h6622631800a78733050eb6a787930000, /*  785 */
128'h97aa00070023c319676200070023c319, /*  786 */
128'h080c460100f618634785cb114501e398, /*  787 */
128'h452d8082612170e22501a02ff0ef0828, /*  788 */
128'hf0d2f4cef8cafca6e122e5067175bfe5, /*  789 */
128'h84aa89320005302316050c63e42eecd6, /*  790 */
128'h65a2e91d25019ceff0ef1028002c8a79, /*  791 */
128'he11964062501b61ff0efe4be1028083c, /*  792 */
128'h10078e6301f9799301c977934519e011, /*  793 */
128'h2501e7dff0ef102800f517634791c115, /*  794 */
128'h6ae67a0679a6794674e6640a60aac905, /*  795 */
128'h7793f3fd8bc5451d00b4478380826149, /*  796 */
128'ha02108090a6300897913fff945210049, /*  797 */
128'h02100713046007937a220089e9936406, /*  798 */
128'h000407a30004072300f40ca300f408a3, /*  799 */
128'h00e40c2300040ba300040b2300e40823, /*  800 */
128'h00040f2300040ea300040e23000405a3, /*  801 */
128'h4785f9bfe0ef85a2000a450300040fa3, /*  802 */
128'h00040aa300040a2300040da300040d23, /*  803 */
128'h855285ca0209036300fa02230005091b, /*  804 */
128'h397d7522fd212501e1fff0ef030a2a83, /*  805 */
128'hf793f139250180cff0ef0125262385d6, /*  806 */
128'h0309278385a279220209e993c3990089, /*  807 */
128'h00094503000485a3d09c01348523f480, /*  808 */
128'h5783daffe0ef01c40513c8c8f35fe0ef, /*  809 */
128'h0124b0230004ae230004a623c8880069, /*  810 */
128'h00b44783ee051de3bdf5450100f49423, /*  811 */
128'h00e300297913ee0716e30107f7134511, /*  812 */
128'hbdd14525bf51ec079ee3451d8b85fa09, /*  813 */
128'hf0caf4a6fc86e4d6e8d2eccef8a27119, /*  814 */
128'h0006a023ec6ef06af466f862fc5ee0da, /*  815 */
128'h0005099be85fe0ef8ab6e4328a2e842a, /*  816 */
128'h0007899bc39d662200b4478300099863, /*  817 */
128'h6aa66a4669e6790674a6854e744670e6, /*  818 */
128'h808261096de27d027ca27c427be26b06, /*  819 */
128'h445c0104290316078c638b8500a44783, /*  820 */
128'h0b930006091b00f67463893e40f907bb, /*  821 */
128'hfa090ae35cfd03040b131ff00c132000, /*  822 */
128'h00975d1b6008120791631ff777934458, /*  823 */
128'h19630ffd7d1301a7fd3337fd00254783, /*  824 */
128'h05a3478900a7ec6347854848eb11020d, /*  825 */
128'hb7e52501bc6ff0ef4c0cbfb5498900f4, /*  826 */
128'hcc08b795498500f405a3478501951763, /*  827 */
128'hd5792501b86ff0efe43e853e4c0c601c, /*  828 */
128'h072c7a6367a28dc200a6083b000d061b, /*  829 */
128'h00e6f46300c4873b0099549b0027c683, /*  830 */
128'h50ef85d2864286a60017c50341a684bb, /*  831 */
128'hc3850407f79300a44783f94525010d20, /*  832 */
128'h15020097951b0097fc6341b507bb4c48, /*  833 */
128'h949bc3ffe0ef955285da200006139101, /*  834 */
128'h4099093b445c9a3e9381020497930094, /*  835 */
128'hbf3900faa0239fa5000aa783c45c9fa5, /*  836 */
128'hc30d0407771300a44703050601634c50, /*  837 */
128'h2501098050efe44285da46850017c503, /*  838 */
128'h00f40523fbf7f793682200a44783f131, /*  839 */
128'h044050ef85da0017c50386424685601c, /*  840 */
128'hf5930009049b444c01b42e23f10d2501, /*  841 */
128'h85930007049b0127746340bb873b1ff5, /*  842 */
128'h499dbf9dbb1fe0ef855295a286260305, /*  843 */
128'hfc86e4d6e8d2eccef0caf8a27119b585, /*  844 */
128'ha023ec6ef06af466f862fc5ee0daf4a6, /*  845 */
128'h099bca3fe0ef8ab689328a2e842a0006, /*  846 */
128'h0007899bc39d00b44783000997630005, /*  847 */
128'h6aa66a4669e6790674a6854e744670e6, /*  848 */
128'h808261096de27d027ca27c427be26b06, /*  849 */
128'h0127873b445c1a0782638b8900a44783, /*  850 */
128'h03040b131ff00c1320000b9304f76e63, /*  851 */
128'h140794631ff777930409046344585cfd, /*  852 */
128'h01a7fd3337fd0025478300975d1b6008, /*  853 */
128'hcb914581485cef01040d1a630ffd7d13, /*  854 */
128'hb749498900f405a3478902e798634705, /*  855 */
128'h4818445cf3fd0005079bd6aff0ef4c0c, /*  856 */
128'h00f405230207e79300a4478312f76b63, /*  857 */
128'hbf89498500f405a3478501979763b785, /*  858 */
128'h0407f79300a44783c85ce311cc1c4858, /*  859 */
128'h40ef85da0017c50346854c50601cc38d, /*  860 */
128'h0523fbf7f79300a44783f96925017350, /*  861 */
128'h2501964ff0efe43e853e4c0c601c00f4, /*  862 */
128'h7a6367a28db200a8063b000d081bd159, /*  863 */
128'hf4630104873b0099549b0027c683072c, /*  864 */
128'h40ef85d286a60017c50341a684bb00e6, /*  865 */
128'h0297f26341b587bb4c4cf14925016e50, /*  866 */
128'h855a95d220000613918115820097959b, /*  867 */
128'h00f40523fbf7f79300a44783a29fe0ef, /*  868 */
128'h093b445c9a3e9381020497930094949b, /*  869 */
128'h00faa0239fa5000aa783c45c9fa54099, /*  870 */
128'h00d77a634458481400c70e634c58bdc9, /*  871 */
128'hfd012501649040ef85da46850017c503, /*  872 */
128'h873b1ff575130009049b444801b42e23, /*  873 */
128'h8626030505130007049b0127746340ab, /*  874 */
128'h0407e79300a447839b5fe0ef952285d2, /*  875 */
128'h1141bd15499db5f1c81cbf4100f40523, /*  876 */
128'h4783e16d2501ab7fe0ef842ae406e022, /*  877 */
128'h601cc3950407f793cf610207f71300a4, /*  878 */
128'h607040ef030405930017c50346854c50, /*  879 */
128'h00f40523fbf7f79300a44783ed4d2501, /*  880 */
128'hc703741ce1552501b5ffe0ef6008500c, /*  881 */
128'h0107169b481800e785a30207671300b7, /*  882 */
128'h00d78ea300e78e230086d69b0106d69b, /*  883 */
128'h00e78fa300d78f230187571b0107569b, /*  884 */
128'h169b00e78d2300078ba300078b234858, /*  885 */
128'h571b0107171b00e78a230107571b0107, /*  886 */
128'h07130106d69b00e78aa30087571b0107, /*  887 */
128'h8da3046007130086d69b00e78c230210, /*  888 */
128'h4783000789a30007892300e78ca300d7, /*  889 */
128'h0223478500f40523fdf7f793600800a4, /*  890 */
128'h60a24505ea3fe06f014160a2640200f5, /*  891 */
128'hf0ef842ae406e0221141808201416402, /*  892 */
128'he11925019b5fe0ef8522e9012501f01f, /*  893 */
128'he42a110180820141640260a200043023, /*  894 */
128'h0000879700054a63945fe0efec060028, /*  895 */
128'hbfe5452d8082610560e2450148a78623, /*  896 */
128'heca6f486f0a21028002c4601e42a7159, /*  897 */
128'h1028083c65a2ec190005041bb25fe0ef, /*  898 */
128'he9916586e41d0005041bcb4ff0efe4be, /*  899 */
128'h616564e6740670a68522cbd8575277a2, /*  900 */
128'h0004c50374a2cb998bc100b5c7838082, /*  901 */
128'h4415fcf41ee34791b7c5c8c8965fe0ef, /*  902 */
128'hf4cef8cae122e506e42afca67175bfd9, /*  903 */
128'hab9fe0ef1828002c460184ae00050023, /*  904 */
128'h02f00913842677e2ecbe081ce5212501, /*  905 */
128'he50567a24501040991634996c2be4bdc, /*  906 */
128'h00e780230307071b3d87470300008717, /*  907 */
128'h02f007130e94156300e780a303a00713, /*  908 */
128'h74e6640a60aa00078023078d00e78123, /*  909 */
128'hf75fe0ef182845858082614979a67946, /*  910 */
128'hf55d2501e6cff0ef18284581fd4d2501, /*  911 */
128'h4581c2aa8bdfe0ef0007c50365c677e2, /*  912 */
128'hf0ef18284581f9512501f4ffe0ef1828, /*  913 */
128'he0ef0007c50365c677e2e1052501e46f, /*  914 */
128'ha86ff0ef1828458101350e632501897f, /*  915 */
128'hb7614509f6e512e367a24711dd612501, /*  916 */
128'h9301020797134781f48fe0ef1828100c, /*  917 */
128'h60630037871be705fc97470397361094, /*  918 */
128'h930102069713662236fd86a285be04e4, /*  919 */
128'hbf199c3d01260023fff7c793e989963a, /*  920 */
128'h930117020007059bfff5871bb7e12785, /*  921 */
128'h4545b7e900e60023fc974703972a1088, /*  922 */
128'h4703973692810204169367220789bdf5, /*  923 */
128'hb721fe9465e3fee78fa3240507850007, /*  924 */
128'he456e852ec4efc06f04af426f8227139, /*  925 */
128'h000917630005091bfa8fe0ef84ae842a, /*  926 */
128'h854a744270e20007891bcf8900b44783, /*  927 */
128'h4818808261216aa26a4269e2790274a2, /*  928 */
128'h445884bae3918b8900a4478300977763, /*  929 */
128'hc81cfcf778e34818445ce4bd00042623, /*  930 */
128'h4481bf7d00f405230207e79300a44783, /*  931 */
128'h4783fc960ee34c50d3e51ff7f793445c, /*  932 */
128'h4685601cc3850407f7930304099300a4, /*  933 */
128'h4783ed51250129d040ef0017c50385ce, /*  934 */
128'h86264685601c00f40523fbf7f79300a4, /*  935 */
128'hcc44ed35250124b040ef85ce0017c503, /*  936 */
128'h377dc7290097999b002547836008bf59, /*  937 */
128'h02c6ed630337563b0336d6bbfff4869b, /*  938 */
128'hd1c19c9dc45c27814c0c8ff9413007bb, /*  939 */
128'hf793c45c9fa5445c0499ea634a855a7d, /*  940 */
128'hd49bcd112501c79fe0ef6008d7b51ff4, /*  941 */
128'h059b802ff0efe595484cbfb19ca90094, /*  942 */
128'h490900f405a3478900f5976347850005, /*  943 */
128'h490500f405a3478500f5976357fdbded, /*  944 */
128'h8b89600800a44783b765cc0cc84cb5ed, /*  945 */
128'hbf6984cee5990005059bfcbfe0efcb81, /*  946 */
128'hfabafee3fd4588e30005059bc3ffe0ef, /*  947 */
128'h413484bbcc0c445cfaf5fae34f9c601c, /*  948 */
128'he42ef822fc067139b7bdc45c013787bb, /*  949 */
128'h2501fdafe0ef0828002c4601842ac52d, /*  950 */
128'hf0eff01c101ce01c852265a267e2e115, /*  951 */
128'h8bc100b5c783cd996c0ce5292501968f, /*  952 */
128'h0007c50367e2a02d000430234515e789, /*  953 */
128'h0067d7838522458167e2c448e24fe0ef, /*  954 */
128'hfcf50be347912501cadfe0ef00f41423, /*  955 */
128'h4791bfdd452580826121744270e2f971, /*  956 */
128'he0ef842ae406e0221141b7c1fcf501e3, /*  957 */
128'h0141640260a200043023e1192501daef, /*  958 */
128'h892e842af406e84aec26f02271798082, /*  959 */
128'h458100091f63e8890005049bd8cfe0ef, /*  960 */
128'h8526740270a20005049bc4ffe0ef8522, /*  961 */
128'h85224581022430238082614564e26942, /*  962 */
128'h00042a2302f5136347912501b34ff0ef, /*  963 */
128'hf77fe0ef85224581c58fe0ef852285ca, /*  964 */
128'hd16dbf7d00042a2300f5166347912501, /*  965 */
128'h002c460184aee42aeca67159bf6584aa, /*  966 */
128'he00d0005041becefe0eff486f0a21028, /*  967 */
128'h0005041b85eff0efe4be1028083c65a2, /*  968 */
128'hc00fe0ef102885a6c489cf816786e801, /*  969 */
128'hbfcd44198082616564e6740670a68522, /*  970 */
128'h002c46018b2ee42af85a8432f0a27159, /*  971 */
128'hf45efc56e4cee8caeca6f486e0d28522, /*  972 */
128'h000a1c6300050a1be70fe0efec66f062, /*  973 */
128'h02f76263ffec871b481c01842c836000, /*  974 */
128'h69a6694664e68552740670a600fb2023, /*  975 */
128'h808261656ce27c027ba27b427ae26a06, /*  976 */
128'h59fd4481490902fb9f63478500044b83, /*  977 */
128'h093508632501a49fe0ef852285ca4a85, /*  978 */
128'hfef963e329054c1c2485e11109550863, /*  979 */
128'h202300f402a30017e793c80400544783, /*  980 */
128'h44814981490110000ab7504cb74d009b, /*  981 */
128'he0ef0015899b852200099e631afd4c09, /*  982 */
128'h200009930344091385cee9212501d04f, /*  983 */
128'h0087979b0009470300194783038b9163, /*  984 */
128'hfc0c94e33cfd39f909092485e3918fd9, /*  985 */
128'h015575332501aa2fe0efe02e854ab745, /*  986 */
128'hb7494a05b7c539f109112485e1116582, /*  987 */
128'hec06e426e8221101bfad8a2abfbd4a09, /*  988 */
128'h4783e4910005049bbb8fe0ef842ae04a, /*  989 */
128'h69028526644260e20007849bcb9100b4, /*  990 */
128'hcf390027f71300a447838082610564a2, /*  991 */
128'h0523c8180207e793fed772e348144458, /*  992 */
128'h2a232501a5aff0ef484cef01600800f4, /*  993 */
128'he0ef4c0cbf7d84aa00a405a3c5390004, /*  994 */
128'hb7dd450502f9146357fd0005091b941f, /*  995 */
128'hf9792501b25fe0ef167d100006374c0c, /*  996 */
128'hb769449db7e12501a1eff0ef85ca6008, /*  997 */
128'hfcf96ae34d1c6008fcf900e345094785, /*  998 */
128'h46854c50601cdba50407f79300a44783, /*  999 */
128'hf55d250167a040ef030405930017c503, /* 1000 */
128'h7175b7b100f40523fbf7f79300a44783, /* 1001 */
128'hf8cafca6e122e5061008002c4605e42a, /* 1002 */
128'he0be1008081c65a2e9052501c94fe0ef, /* 1003 */
128'h00b7c78345196786e1052501e27fe0ef, /* 1004 */
128'hf79300b5c483c59975e2eb890207f793, /* 1005 */
128'h6149794674e6640a60aa451dcb810014, /* 1006 */
128'h0005041baccfe0ef0009450379028082, /* 1007 */
128'h0613fc878de301492783c89d88c1cc0d, /* 1008 */
128'hcaa200a84589952fe0ef00a8100c0280, /* 1009 */
128'h838ff0ef00a84581f1612501941fe0ef, /* 1010 */
128'h9e3fe0ef1008faf518e34791d94d2501, /* 1011 */
128'hbf612501f12fe0ef7502e411f1552501, /* 1012 */
128'h7171b7edf551250191eff0ef85a27502, /* 1013 */
128'he94aed26f506f1221028002c4605e42a, /* 1014 */
128'he8eaece6f0e2f4def8dafcd6e152e54e, /* 1015 */
128'h083c65a21c0412630005041bbc4fe0ef, /* 1016 */
128'h1c0407630005041bd53fe0efe4be1028, /* 1017 */
128'hf79300b7c783441967a61af415634791, /* 1018 */
128'h049bb33fe0ef4581752218079d630207, /* 1019 */
128'h16f48c63440975224785180480630005, /* 1020 */
128'h0005041ba8cfe0ef16f48863440557fd, /* 1021 */
128'he0ef85220104d91b85a6742216041263, /* 1022 */
128'h00050c1b45812000061303440b13f60f, /* 1023 */
128'he0ef855a02000593462d886fe0ef855a, /* 1024 */
128'h0109191b0104999b0ff97a9347c187af, /* 1025 */
128'h0109591b021007930109d99b02f40fa3, /* 1026 */
128'h046007930ff4fa1304f4062302e00b93, /* 1027 */
128'h0200061304f406a30089591b0089d99b, /* 1028 */
128'h05440723040405a30404052303740a23, /* 1029 */
128'h051385da052404a305540423053407a3, /* 1030 */
128'h4603468d05740aa37722ff7fd0ef0544, /* 1031 */
128'h478100f69363571400d6166357d20007, /* 1032 */
128'h06f404230107d79b0107969b06f40723, /* 1033 */
128'h0086d69b0107d79b0106d69b0107979b, /* 1034 */
128'h00274b8306f404a306d407a30087d79b, /* 1035 */
128'h0005041bf5ffe0ef1028040b99634c85, /* 1036 */
128'h0210071300e785a3752247416786e835, /* 1037 */
128'h00078ba300078b230460071300e78c23, /* 1038 */
128'h01578a2301378da301478d2300e78ca3, /* 1039 */
128'h041bd50fe0ef00f50223478501278aa3, /* 1040 */
128'h022303852823001c0d1b7522a82d0005, /* 1041 */
128'h20000613ec090005041b8d4fe0ef0195, /* 1042 */
128'h8c6a0ffbfb93f53fd0ef3bfd855a4581, /* 1043 */
128'h70aa8522f2bfe0ef85a67522441db749, /* 1044 */
128'h7ba67b467ae66a0a69aa694a64ea740a, /* 1045 */
128'h7159b7c544218082614d6d466ce67c06, /* 1046 */
128'h10284605002c843284aee42aeca6f0a2, /* 1047 */
128'h1028083c65a2e13125019c2fe0eff486, /* 1048 */
128'hc783451967a6e9152501b55fe0efe4be, /* 1049 */
128'h00b74783c30d6706e39d0207f79300b7, /* 1050 */
128'h008705a38c3d027474138c658cbd7522, /* 1051 */
128'h740670a62501c94fe0ef00f502234785, /* 1052 */
128'h002c4605e02ee42a71718082616564e6, /* 1053 */
128'h0005079b95cfe0efed26f122f5060088, /* 1054 */
128'hf0be083cf4be008865a2678612079563, /* 1055 */
128'hc7037786100799630005079bae7fe0ef, /* 1056 */
128'h479165e61007116302077713479900b7, /* 1057 */
128'h0613e3ffd0ef102805ad46550e058d63, /* 1058 */
128'hefdfd0ef850ae33fd0ef10a8008c0280, /* 1059 */
128'h079ba9dfe0ef10a865820c054c6347ad, /* 1060 */
128'hdcbfe0ef10a80ce792634711cbf10005, /* 1061 */
128'h851302a10593464d648aebdd0005079b, /* 1062 */
128'h0207e793640602814783df7fd0ef00d4, /* 1063 */
128'h8bc100b4c78300f40223478500f485a3, /* 1064 */
128'h85a60004450306f7076357d64736cbb5, /* 1065 */
128'h059bca4fe0ef85220005059bf25fd0ef, /* 1066 */
128'h0005079bfbbfd0ef8522c1bd47890005, /* 1067 */
128'h02f69c630557468302e007936706efa9, /* 1068 */
128'h04230107d79b06f707230107969b57d6, /* 1069 */
128'hd69b0087d79b0107d79b0107979b06f7, /* 1070 */
128'h06d707a3478506f704a30086d69b0106, /* 1071 */
128'he7910005079be18fe0ef008800f70223, /* 1072 */
128'h64ea740a70aa0005079bb48fe0ef6506, /* 1073 */
128'he42ae8a2711dbfcd47a18082614d853e, /* 1074 */
128'h250180afe0efec861028002c4605842e, /* 1075 */
128'h250199dfe0efe4be1028083c65a2e929, /* 1076 */
128'heb950207f79300b7c783451967a6e129, /* 1077 */
128'h571b00e78b23752200645703cb856786, /* 1078 */
128'h571b00e78c230044570300e78ba30087, /* 1079 */
128'hacefe0ef00f50223478500e78ca30087, /* 1080 */
128'he0cae4a6711d80826125644660e62501, /* 1081 */
128'hec86e8a208284601002c893284aee42a, /* 1082 */
128'h08284581c4b9e0510005041bf95fd0ef, /* 1083 */
128'he0ef08284585e5592501c9efe0efd202, /* 1084 */
128'hc8dfd0ef8526462d75c2e93d2501b97f, /* 1085 */
128'hce89000700230200061346ad00b48713, /* 1086 */
128'hc78397a6938117820007869bfff6879b, /* 1087 */
128'h510c656202090a63fec783e3177d0007, /* 1088 */
128'h0793470d6562e0150005041be63fd0ef, /* 1089 */
128'h87930270079300e68463000546830430, /* 1090 */
128'h60e6852200a92023c15fd0ef953e0347, /* 1091 */
128'h00f51563479180826125690664a66446, /* 1092 */
128'h4605e42a711db7d5842abf5500048023, /* 1093 */
128'h0005041beddfd0efec86e8a21028002c, /* 1094 */
128'h930102079713478100010c236522e471, /* 1095 */
128'h4581ebb102000613eb2900074703972a, /* 1096 */
128'h4585e0450005041bbccfe0efda021028, /* 1097 */
128'h01814783100515632501ac3fe0ef1028, /* 1098 */
128'h07136786bb1fd0ef082c462dc7e56506, /* 1099 */
128'h8ba300078b230460071300e78c230210, /* 1100 */
128'hb77d87bab7452785a0e900e78ca30007, /* 1101 */
128'h0006c68396aa928102071693fff7871b, /* 1102 */
128'hc58300e506b3432d48e54701fec686e3, /* 1103 */
128'hf9f6881b92c1030596930017061b0006, /* 1104 */
128'h92c116c236810108ec63030858131842, /* 1105 */
128'h959ba83100068e1b8f85859300007597, /* 1106 */
128'h60e685224419feb045e34185d59b0185, /* 1107 */
128'h000805630005c8030585808261256446, /* 1108 */
128'h070595ba082cfe6702e3b7ddffc81be3, /* 1109 */
128'h02061793f8f6e9e30007069b00d58023, /* 1110 */
128'h00d779630007869b0200061347299381, /* 1111 */
128'h0834b77df0f713e30e50079301814703, /* 1112 */
128'h00f500235795b7c5078500c6802396be, /* 1113 */
128'h0005041b8b2fe0ef00f5022347857522, /* 1114 */
128'h1028d3c10181478302f51b634791b771, /* 1115 */
128'h020006136506f8350005041ba19fe0ef, /* 1116 */
128'ha8dfd0ef082c462d6506ab7fd0ef4581, /* 1117 */
128'h2e83bf81842abdd100e785a347216786, /* 1118 */
128'h110105c528830585230305452e030505, /* 1119 */
128'h869a8646040502938f2ae44ae826ec22, /* 1120 */
128'h00c6c5b33ecf8f9300005f97887687f2, /* 1121 */
128'ha403000f2583000fa38300b647338dfd, /* 1122 */
128'h2703ff4fa3839db9007585bb0fc1008f, /* 1123 */
128'he8330198581b0078159b0105883b004f, /* 1124 */
128'h00f6c6339f3100f805bb0077073b0105, /* 1125 */
128'h561b00c6171b9e39008f23838e358e6d, /* 1126 */
128'h00d383bb00c5873b008383bb8e590146, /* 1127 */
128'h007686bb8ebd00cf24038ef900b7c6b3, /* 1128 */
128'ha4039fa100d3e6b30116969b00f6d39b, /* 1129 */
128'h007777338f2d0007061b00d703bbffcf, /* 1130 */
128'h8f5d0167171b00a7579b9f3d8f2d9fa1, /* 1131 */
128'h17e300e387bb0003869b0005881b0f41, /* 1132 */
128'h8f9300005f9742ef0f1300005f17f45f, /* 1133 */
128'h8df100d7c5b342e2829300005297366f, /* 1134 */
128'h002f4403001f4383000fa58300b6c733, /* 1135 */
128'h4318972a070a93aa038a000f47039db9, /* 1136 */
128'h159b0105883b004fa7039db9942a040a, /* 1137 */
128'h0105e8330003a70301b8581b9e390058, /* 1138 */
128'h9e398e3d8e7500b7c6339f3100f805bb, /* 1139 */
128'h40189eb90176561b0096139b008fa703, /* 1140 */
128'h0075c6b30f119f3500c583bb00c3e633, /* 1141 */
128'hffcfa7039eb90fc18eadffff44838efd, /* 1142 */
128'h40980126d69b9fb900e6941b94aa048a, /* 1143 */
128'h47338f6d0083c7339fb900d3843b8ec1, /* 1144 */
128'h881b8f5d0147171b00c7579b9f3d0077, /* 1145 */
128'h1ee300e407bb0004069b0003861b0005, /* 1146 */
128'h0000539782fe34ef8f9300005f97f25f, /* 1147 */
128'h00d7c5b30003a7030102c4032c438393, /* 1148 */
128'h0112c4839f25400000c5c4b3942a040a, /* 1149 */
128'h083b40809e2194aa048a0043a4039f21, /* 1150 */
128'h683301c8581b0048171b0122c4830107, /* 1151 */
128'h8db9048a00f8073b0083a4039e210107, /* 1152 */
128'h0132c90300b6159b40809e2d9ea194aa, /* 1153 */
128'ha4839c3500c705bb03c18e4d0156561b, /* 1154 */
128'h941b992a9ea1090a8ead00e7c6b3ffc3, /* 1155 */
128'h843b8ec1000924830106d69b9fa50106, /* 1156 */
128'h579b9f3d8f219fa58f2d0007081b00d5, /* 1157 */
128'h069b0005861b02918f5d0177171b0097, /* 1158 */
128'h829300005297f45f17e300e407bb0004, /* 1159 */
128'h0002a70300d745b38f5dfff647132462, /* 1160 */
128'h038a020fc5839f2d022fc403021fc383, /* 1161 */
128'ha5839f2d942a040a418c95aa058a93aa, /* 1162 */
128'h0003a5839e2d0068171b0107083b0042, /* 1163 */
128'hc6139db100f8073b0107683301a8581b, /* 1164 */
128'h00a6139b0082a5839e2d8e3d8e59fff6, /* 1165 */
128'h00c703bb00c3e633400c9ead0166561b, /* 1166 */
128'h02c10075e5b3fff7c593023fc4839ead, /* 1167 */
128'h94aa00f5969b048a9db5ffc2a4038db9, /* 1168 */
128'h081b00b385bb40809fa18dd50115d59b, /* 1169 */
128'h9f3d007747339fa18f4dfff747130007, /* 1170 */
128'h0003861b0f918f5d0157171b00b7579b, /* 1171 */
128'h883b6462f3ff1de300e587bb0005869b, /* 1172 */
128'h282300c8863b00d306bb00fe07bb010e, /* 1173 */
128'h80826105692264c2cd70cd34c97c0505, /* 1174 */
128'he45ee85af44ef84afc26e0a2715d653c, /* 1175 */
128'h89ae84aa97b203f7f413ec56f052e486, /* 1176 */
128'h408b07bb04000b9304000b13e53c8932, /* 1177 */
128'h00090a1b00f974639381178200078a1b, /* 1178 */
128'h86560084853385ce020ada93020a1a93, /* 1179 */
128'h176399d6415909334a7020ef0144043b, /* 1180 */
128'h640660a6b7c997824401852660bc0174, /* 1181 */
128'h61616ba26b426ae27a0279a2794274e2, /* 1182 */
128'hec26842a03f7f793f0227179653c8082, /* 1183 */
128'h97a2f800071300178513e84af406e44e, /* 1184 */
128'h091b40a9863b449d0400099300e78023, /* 1185 */
128'hf5633f3020ef95224581920116020006, /* 1186 */
128'h450197828522603cfc1c078e643c0124, /* 1187 */
128'h614569a2694264e2740270a2fd24fde3, /* 1188 */
128'h04053423639cf5678793000077978082, /* 1189 */
128'h0797ed3c639cf4e7879300007797e93c, /* 1190 */
128'h0505059311018082e13cb80787930000, /* 1191 */
128'h0000769747013e5020efec06850a4641, /* 1192 */
128'h07b34541394585930000659720468693, /* 1193 */
128'h962e0047d613070506890007c78300e1, /* 1194 */
128'hfec68f230007c78397ae000646038bbd, /* 1195 */
128'h05130000751760e2fca71de3fef68fa3, /* 1196 */
128'he5060808842ae1227175808261051c65, /* 1197 */
128'he85ff0ef080885a26622f71ff0efe42e, /* 1198 */
128'h640a60aaf83ff0ef0808f01ff0ef0808, /* 1199 */
128'h469100d70d63711c46a1595880826149, /* 1200 */
128'hac2380824501cf980200071300d71763, /* 1201 */
128'hec06e426e82211018082556dbfe50007, /* 1202 */
128'h0000569702f5026384ae842a200007b7, /* 1203 */
128'h2f8585930000659708800613ff468693, /* 1204 */
128'h60e2fc2412f030ef3085051300006517, /* 1205 */
128'he4266100e82211018082610564a26442, /* 1206 */
128'h0000569702f4026384ae200007b7ec06, /* 1207 */
128'h2b8585930000659702f00613fcc68693, /* 1208 */
128'h60e2e0040ef030ef2c85051300006517, /* 1209 */
128'he4266100e82211018082610564a26442, /* 1210 */
128'h0000569702f4026384ae200007b7ec06, /* 1211 */
128'h278585930000659703600613f9c68693, /* 1212 */
128'h60e2e4040af030ef2885051300006517, /* 1213 */
128'he8226104e42611018082610564a26442, /* 1214 */
128'h0000769702f48263842e200007b7ec06, /* 1215 */
128'h238585930000659703e00613e1c68693, /* 1216 */
128'h9001140206f030ef2485051300006517, /* 1217 */
128'he42611018082610564a2644260e2e880, /* 1218 */
128'h02f48263842e200007b7ec06e8226104, /* 1219 */
128'h0000659704500613dd06869300007697, /* 1220 */
128'h02b030ef20450513000065171f458593, /* 1221 */
128'h8082610564a2644260e2ec8090011402, /* 1222 */
128'h84ae200007b7ec06e4266100e8221101, /* 1223 */
128'h04c00613ee4686930000569702f40263, /* 1224 */
128'h1c050513000065171b05859300006597, /* 1225 */
128'h8082610564a2644260e2f0047e6030ef, /* 1226 */
128'h84ae200007b7ec06e4266100e8221101, /* 1227 */
128'h05300613eb4686930000569702f40263, /* 1228 */
128'h18050513000065171705859300006597, /* 1229 */
128'h8082610564a2644260e2f4047a6030ef, /* 1230 */
128'hfc06f04af426f82200053983ec4e7139, /* 1231 */
128'h569702f984638436893284ae200007b7, /* 1232 */
128'h85930000659705a00613e7a686930000, /* 1233 */
128'h75a030efe43a13650513000065171265, /* 1234 */
128'h79130029191b8b0588090014141b6722, /* 1235 */
128'h8c4588a1012464330034949b8c590049, /* 1236 */
128'h612169e2790274a2744270e20289b823, /* 1237 */
128'h85224605468147057100e02211418082, /* 1238 */
128'hf35ff0ef45818522f7dff0efe4064581, /* 1239 */
128'h6008f67ff0ef45814605468547058522, /* 1240 */
128'h808201414501640260a2d97ff0ef4581, /* 1241 */
128'h02053c23460546814705e022e4061141, /* 1242 */
128'h45818522f39ff0ef842a458104053023, /* 1243 */
128'hf0ef46054685470545818522ef1ff0ef, /* 1244 */
128'hd4dff06f0141458160a264026008f23f, /* 1245 */
128'h842e200007b7ec06e8226104e4261101, /* 1246 */
128'h06100613da4686930000569702f48263, /* 1247 */
128'h05050513000065170405859300006597, /* 1248 */
128'h64a2644260e2fc8090411442676030ef, /* 1249 */
128'h07b7ec06e8226104e426110180826105, /* 1250 */
128'hd70686930000569702f48263842e2000, /* 1251 */
128'h00006517ffc585930000659706800613, /* 1252 */
128'h60e2e0a090511452632030ef00c50513, /* 1253 */
128'he4266100e82211018082610564a26442, /* 1254 */
128'h0000569702f4026384ae200007b7ec06, /* 1255 */
128'hfb8585930000659706f00613d3c68693, /* 1256 */
128'h60e2e4245ee030effc85051300006517, /* 1257 */
128'h00053903e04a11018082610564a26442, /* 1258 */
128'h026384ae842a200007b7ec06e426e822, /* 1259 */
128'h659707600613d06686930000569702f9, /* 1260 */
128'h30eff825051300006517f72585930000, /* 1261 */
128'h690264a2644260e2c84404993c235a80, /* 1262 */
128'hf486e8caeca67100f0a2715980826105, /* 1263 */
128'h08a3ec66f062f45ef85afc56e0d2e4ce, /* 1264 */
128'h4611d01ce03084b2892e0005d7830204, /* 1265 */
128'h60080e049c636f6020ef00c905134581, /* 1266 */
128'h3a03200007b700043983bf7ff0ef4585, /* 1267 */
128'h0017f71344810049278316f99a630404, /* 1268 */
128'h03243c234c1c4485e391448d8b89c709, /* 1269 */
128'h160786638b85008a2783000a09638cdd, /* 1270 */
128'hf0ef852245814605468147050144e493, /* 1271 */
128'h852200892583be3ff0ef85224581d73f, /* 1272 */
128'h0a13852200095583c55ff0ef00989a37, /* 1273 */
128'h4581cc7ff0ef852285a6c8bff0ef681a, /* 1274 */
128'h85224581460546854705cffff0ef8522, /* 1275 */
128'hf0ef852224058593000f45b7d31ff0ef, /* 1276 */
128'h85220d89b583cdbff0ef85224585e9bf, /* 1277 */
128'hf0ef25810015e593c30c8c9300005c97, /* 1278 */
128'h0b1300006b17e4ea8a9300006a97ebbf, /* 1279 */
128'h69a6694664e6740670a6efe9485ce5eb, /* 1280 */
128'h616545016ce27c027ba27b427ae26a06, /* 1281 */
128'h8522488cdb9ff0efe024852244cc8082, /* 1282 */
128'h3883603cee079be38b85449cdf5ff0ef, /* 1283 */
128'h47014781458163900107e68365410004, /* 1284 */
128'hec0689e36e89f005051300ff0e374311, /* 1285 */
128'he7b301e8183b070500371f1b00064803, /* 1286 */
128'hd81bf2e50067036316fd060527810107, /* 1287 */
128'h78330087981b010767330187971b0187, /* 1288 */
128'h873b8fd98fe9010767330087d79b01c8, /* 1289 */
128'h2585e31c9746938183751782170200be, /* 1290 */
128'h0613b226869300005697b76547014781, /* 1291 */
128'h051300006517d7e58593000065971490, /* 1292 */
128'h8bd2bd6100c4e493bd853b4030efd8e5, /* 1293 */
128'h859300005597000b9d633bfd20000c37, /* 1294 */
128'hb711702000efd7e5051300006517b065, /* 1295 */
128'h85d60f20061386e60189096300043903, /* 1296 */
128'h8cfd4981485c07093483374030ef855a, /* 1297 */
128'h6f630c89378302093703140480632481, /* 1298 */
128'h85224581cc5cf9200793c7817c1c00f7, /* 1299 */
128'h0044f793b29ff0ef85224581b71ff0ef, /* 1300 */
128'h00896913ff397913852201442903c39d, /* 1301 */
128'h05130000651785cad45ff0ef85ca2901, /* 1302 */
128'h01442903c39d0084f79368a000efd1e5, /* 1303 */
128'hf0ef85ca290100496913ff3979138522, /* 1304 */
128'h660000efd1c505130000651785cad1bf, /* 1305 */
128'h8c630384390300043983cfb50014f793, /* 1306 */
128'h85d609c00613a6e68693000056970189, /* 1307 */
128'h3c2300492783cba97c1c2c4030ef855a, /* 1308 */
128'h0189871308e69f630037f693470d0204, /* 1309 */
128'hff87051363104591480d468100c90793, /* 1310 */
128'h8361ff87370301068763c3900086161b, /* 1311 */
128'h603cfeb690e30791872a2685c3988f51, /* 1312 */
128'hc85c9bf9485cc85c0027e793485ccbb5, /* 1313 */
128'h01848c63040439036004cc9d49858889, /* 1314 */
128'h855a85d60ca00613a086869300005697, /* 1315 */
128'h008927830009096304043023246030ef, /* 1316 */
128'h9bf54985485cb4bff0ef8522ef8d8b85, /* 1317 */
128'h4505d8098ce3c43ff0ef8522484cc85c, /* 1318 */
128'h26230009b783dbd98b85bd85645020ef, /* 1319 */
128'h97a667a1bf41b1bff0ef8522b77100f9, /* 1320 */
128'h639c00878913dcd50109648300093983, /* 1321 */
128'h14e109a13c2020efe43e002c4621854e, /* 1322 */
128'h04800513717908b041635535b7dd87ca, /* 1323 */
128'h30ef892e84b2e44ef406e84aec26f022, /* 1324 */
128'h05130000551785a2c41d5551842a1380, /* 1325 */
128'h00006517862285aa89aa7b3010ef9765, /* 1326 */
128'h30ef852200099d63508000efbec50513, /* 1327 */
128'h614569a2694264e2740270a2557d1520, /* 1328 */
128'hf793f40401242423e01c200007b78082, /* 1329 */
128'h45018885bfe94501c45c4789c7890024, /* 1330 */
128'h0537458146098082b7f9c45c4785d8f1, /* 1331 */
128'h638897aa200007b7050ef73ff06f2000, /* 1332 */
128'h07b7e4066380e0221141711c80822501, /* 1333 */
128'h0613912686930000569702f402632000, /* 1334 */
128'h051300006517ace585930000659734c0, /* 1335 */
128'h60a2557de3914505703c104030efade5, /* 1336 */
128'hec064501842ae8221101808201416402, /* 1337 */
128'h468560e26622644285a2501010efe42e, /* 1338 */
128'hf022f4062000051371797a00006f6105, /* 1339 */
128'h651784aa03e030efe052e44ee84aec26, /* 1340 */
128'h10ef0001b503146030efb42505130000, /* 1341 */
128'h681c224010ef842a4bf010ef45014790, /* 1342 */
128'h4583402000ef638cb285051300006517, /* 1343 */
128'h546c3f2000efb26505130000651706f4, /* 1344 */
128'h91c115c20085d59bb305051300006517, /* 1345 */
128'h05130000651706c4458358303dc000ef, /* 1346 */
128'h77130ff677930106569b0086571bb265, /* 1347 */
128'h5c0c3b2000ef0186561b0ff6f6930ff7, /* 1348 */
128'h6597545c3a4000efb185051300006517, /* 1349 */
128'ha905859300006597c789aa2585930000, /* 1350 */
128'h00006517384000efb085051300006517, /* 1351 */
128'h8593000065977448098030efb1450513, /* 1352 */
128'h00006617584c19c42783d65fb0ef0865, /* 1353 */
128'h6517dca6061300006617e789a6c60613, /* 1354 */
128'hf0ef85264581346000efaf2505130000, /* 1355 */
128'h00006997af4a0a1300006a174401ed9f, /* 1356 */
128'h0004059b01f4779320000913af498993, /* 1357 */
128'h0007c583008487b3318000ef8552e781, /* 1358 */
128'h1de3302000ef819100f5f6130405854e, /* 1359 */
128'h70a22f2000ef00e5051300006517fd24, /* 1360 */
128'h8082614545016a0269a2694264e27402, /* 1361 */
128'h40f707b30003b6830083b7830103b703, /* 1362 */
128'hb8230017079300d7fe63938117822785, /* 1363 */
128'h0007802345050103b78300a7002300f3, /* 1364 */
128'h96130103b7830083b703808245018082, /* 1365 */
128'h8e9dfff706930003b7038f9992010205, /* 1366 */
128'h0007869b47819d9dfff7059b00c6f563, /* 1367 */
128'h8082852e0007002300b6e6630103b703, /* 1368 */
128'h0006c68300f506b300d3b82300170693, /* 1369 */
128'he681000556634301bfd900d700230785, /* 1370 */
128'h04100693c21906100693430540a0053b, /* 1371 */
128'hf53b0005089b385986ba4e250ff6f813, /* 1372 */
128'h76130306061b04ae6a630ff5761302b8, /* 1373 */
128'hfcb8ffe302b8d53bfec68fa306850ff6, /* 1374 */
128'he96300a606bb0300059340e0063b8536, /* 1375 */
128'h050500f5002302d007930003076302f6, /* 1376 */
128'hfff5081b46810015559b9d1900050023, /* 1377 */
128'hbf4500c8063b808200b7ea630006879b, /* 1378 */
128'h9381178240f807bbb7d1feb50fa30505, /* 1379 */
128'h0685000648830007c30300d7063397ba, /* 1380 */
128'h011cf0ca7119b7e10117802300660023, /* 1381 */
128'he0dafc86e4d6e8d2eccef4a6f8a2597d, /* 1382 */
128'h02500993f82af02ef42afc3e843684b2, /* 1383 */
128'h77a277420209591303000a9306c00a13, /* 1384 */
128'h178276820017079bc52d8f1d0004c503, /* 1385 */
128'h0201039304850135086304d7ff639381, /* 1386 */
128'h048905450f630014c503bfe1e71ff0ef, /* 1387 */
128'hfd07879bcb9d0004c783035510634781, /* 1388 */
128'h0014c503478100f6f36346a50ff7f793, /* 1389 */
128'h069302a6eb6306d50f63064006930489, /* 1390 */
128'hf55d08f509630630079304d50f630580, /* 1391 */
128'h6b066aa66a4669e6790674a6744670e6, /* 1392 */
128'hb74d048d0024c503808261090007051b, /* 1393 */
128'h0700071300a76c6306e50e6307300713, /* 1394 */
128'ha00d46014685003800840b13f6e51ee3, /* 1395 */
128'hf6e510e30780071302e5006307500713, /* 1396 */
128'h001636134685003800840b13fa850613, /* 1397 */
128'hb693003800840b13f8b50693a81145c1, /* 1398 */
128'h0005059be31ff0ef400845a946010016, /* 1399 */
128'h00044503a809dd1ff0ef002802010393, /* 1400 */
128'hb5fd845ad89ff0ef00840b1302010393, /* 1401 */
128'h501010ef852201247433600000840b13, /* 1402 */
128'hf436715db7f18522020103930005059b, /* 1403 */
128'hf0efe436e4c6e0c2fc3ef83aec061034, /* 1404 */
128'h862ef436f032715d8082616160e2e8df, /* 1405 */
128'he4c6e0c2fc3ef83aec06100005931014, /* 1406 */
128'hf62e710d8082616160e2e69ff0efe436, /* 1407 */
128'hee060808100005931234862afe36fa32, /* 1408 */
128'he3fff0efe436eec6eac2e6bee2baea22, /* 1409 */
128'h6135645260f28522125020ef0808842a, /* 1410 */
128'h8302000303630087b303679c691c8082, /* 1411 */
128'h86930000469704b7ec63479d80824501, /* 1412 */
128'he822ec061101431c9736002597134666, /* 1413 */
128'h7540f55c08c52483795c878297b6e426, /* 1414 */
128'h64a260e2029454330e7010ef90811482, /* 1415 */
128'h617cbff17d5c8082610545016442e900, /* 1416 */
128'h557db7f1659c95aa058e05e135f1bfe1, /* 1417 */
128'hf0ef842ae406e02211418082557d8082, /* 1418 */
128'h07630207b303679c681c00055e63ff5f, /* 1419 */
128'h60a245018302014160a2640285220003, /* 1420 */
128'h00a7eb6347ad8082557d808201416402, /* 1421 */
128'h6108953e81753fe78793000047971502, /* 1422 */
128'h679c691c80826e650513000055178082, /* 1423 */
128'h47d502f1102347a1715d83020007b303, /* 1424 */
128'h07930030e83ee42e078517824785d23e, /* 1425 */
128'h60a6fd3ff0efcc3ed402e486100c2000, /* 1426 */
128'h011308e6e063400407374d1480826161, /* 1427 */
128'h342385a2980101f1041322813823dc01, /* 1428 */
128'he909fadff0ef1a05348322113c232291, /* 1429 */
128'hfb60051300f70d630a0447830a04c703, /* 1430 */
128'h24010113228134832301340323813083, /* 1431 */
128'hc703fef711e30dd447830dd4c7038082, /* 1432 */
128'h47830e04c703fcf71be30c0447830c04, /* 1433 */
128'h0d4485130d4405934611fcf715e30e04, /* 1434 */
128'h717980824501bf654501fd4559b010ef, /* 1435 */
128'h85226ea020eff4063e800513842af022, /* 1436 */
128'hf21ff0efc202c40200011023858a4601, /* 1437 */
128'h70a285226cc020ef7d000513e509842a, /* 1438 */
128'h478500f1102347857179808261457402, /* 1439 */
128'h4538691cc195842ac402c23ef406f022, /* 1440 */
128'h06b78ff58ff9f80686934bdc008006b7, /* 1441 */
128'h4601c43e8fd9400007378fd98f756000, /* 1442 */
128'h70a2c43c47b2e119ec9ff0ef8522858a, /* 1443 */
128'h47d500f1102347b5711d808261457402, /* 1444 */
128'h0107979bf852fc4ee0ca07c55783c23e, /* 1445 */
128'hec86f05ae4a6e8a26a056989fdf94937, /* 1446 */
128'h8993080909134495c43e842e8b2af456, /* 1447 */
128'he71ff0ef855a858a4601e00a0a13e009, /* 1448 */
128'h95630135f7b3c7891005f79345b2ed15, /* 1449 */
128'h5405051300005517c7950125f7b30547, /* 1450 */
128'h690664a6644660e6fba00513d4dff0ef, /* 1451 */
128'hc5e334fd808261257b027aa27a4279e2, /* 1452 */
128'h20ef3e80051300805863fff40a9bfe04, /* 1453 */
128'h5517fc8047e345018456b74d84565d60, /* 1454 */
128'hbf6df9200513d07ff0ef512505130000, /* 1455 */
128'hc42e00f1102347c17139e7a919c52783, /* 1456 */
128'hc23e842af426fc06f822858a460147d5, /* 1457 */
128'h4495cb918b891b842783c11ddddff0ef, /* 1458 */
128'hf8ed34fdc901dc7ff0ef8522858a4601, /* 1459 */
128'h4501bfd545018082612174a2744270e2, /* 1460 */
128'h892a4785e8a2ec86e0cae4a6711d8082, /* 1461 */
128'h02f1102302c9270347c906d7f66384b6, /* 1462 */
128'hcc3ee42e4755d432cf3108c927832601, /* 1463 */
128'hf0efc83eca26d23a854a100c47850030, /* 1464 */
128'h102347b10497f0634785e529842ad6ff, /* 1465 */
128'hf0efd23ed402854a100c47f5460102f1, /* 1466 */
128'hc41ff0ef46c5051300005517c11dd4ff, /* 1467 */
128'h47c580826125690664a6644660e68522, /* 1468 */
128'h4401b7d50004841bb74d02f6063bbf61, /* 1469 */
128'he852ec4ef04af426f822fc067139b7c5, /* 1470 */
128'h10ef8ab684b28a2e4148842ace05e456, /* 1471 */
128'h869fa0ef852200b44583c11d892a4a40, /* 1472 */
128'h551700b67a63014485b3681000054d63, /* 1473 */
128'h2583a0894481bd7ff0ef422505130000, /* 1474 */
128'h0109378389a6f96decdff0ef854a08c9, /* 1475 */
128'h85d6865286a2844e0089f3630207e403, /* 1476 */
128'h89b308c96783fc851ae3f01ff0ef854a, /* 1477 */
128'h70e2fc0999e39aa2028784339a224089, /* 1478 */
128'h61216aa26a4269e274a2790285267442, /* 1479 */
128'h8e55479971390106161b0086969b8082, /* 1480 */
128'hf426f82247f58e5500f11023030006b7, /* 1481 */
128'h8526858a4601440dc432c23e84aafc06, /* 1482 */
128'hd8bff0ef85263e800593e919c4dff0ef, /* 1483 */
128'hbfcdfc79347d8082612174a2744270e2, /* 1484 */
128'h9fb923213823bffc07b7db0101134d18, /* 1485 */
128'h2331342322913c232481302324113423, /* 1486 */
128'h980101f104131ce7f36349013ffc0737, /* 1487 */
128'hb7831e051a63892ac03ff0ef84aa85a2, /* 1488 */
128'h1aa4b0236ee020ef20000513e7991a04, /* 1489 */
128'h10ef85a2200006131e0505631a04b503, /* 1490 */
128'h000047171cf76d6347210c04478313d0, /* 1491 */
128'h8793400407b753b897ba078afa470713, /* 1492 */
128'h071367050d44278300e7fd63cc981ff7, /* 1493 */
128'h4783f8dc00d773630147d69307a68007, /* 1494 */
128'h0019f9938b8506f48f2309b449830a04, /* 1495 */
128'h08f480a30b344783c7890e244783e781, /* 1496 */
128'h09c44783c7898b890a04478300098a63, /* 1497 */
128'h0c848613091407130e24478306f48fa3, /* 1498 */
128'h07c6468109d405130a844783fcdc07c6, /* 1499 */
128'h959b0087979b00074583fff74783e0fc, /* 1500 */
128'h8c634685c39197aeffe745839fad0105, /* 1501 */
128'h87b30dd4478302f585b30e0445830009, /* 1502 */
128'h8f63fce514e30621070de21c07ce02b7, /* 1503 */
128'h0107979b468508d4470308e447830409, /* 1504 */
128'h0e04470397ba08c447039fb90087171b, /* 1505 */
128'hf8fc07ce02e787b30dd4478302f70733, /* 1506 */
128'h0107171b0187979b08a4470308b44783, /* 1507 */
128'h088447039fb90087171b089447039fb9, /* 1508 */
128'h0a044783f4fc07a6c319f4fc54d89fb9, /* 1509 */
128'h4685c6b5e3918bfd09c44783c7898b85, /* 1510 */
128'h4785e141e0bff0ef852645850af00613, /* 1511 */
128'h08f4aa2300a7979b0e0447830af407a3, /* 1512 */
128'hf8dc07a60d44278300098663c79954dc, /* 1513 */
128'h00a7979b02e787bb0dd447030e044783, /* 1514 */
128'h2481308308f480230a74478308f4ac23, /* 1515 */
128'h39832301390323813483854a24013403, /* 1516 */
128'hf3dd8b850af447838082250101132281, /* 1517 */
128'h27058bfd8b7d0057d79b00a7d71b50fc, /* 1518 */
128'hb503892ab75d08f4aa2302f707bb2785, /* 1519 */
128'h5951bf451a04b02354c020efdd4d1a04, /* 1520 */
128'h382322113c23dc010113b7655929b775, /* 1521 */
128'h06f58463478923213023229134232281, /* 1522 */
128'h0b900613842eed8554a9468104b7ec63, /* 1523 */
128'hffe4059be11d84aad3fff0ef892a4585, /* 1524 */
128'h854a85a2980101f10413ed91258199f5, /* 1525 */
128'hdf400493e3990b944783e9159a7ff0ef, /* 1526 */
128'h34832201390385262301340323813083, /* 1527 */
128'h54a94705ffc5879b8082240101132281, /* 1528 */
128'hec267179bfd984aab7554685fef760e3, /* 1529 */
128'h0ff5f99308154783f022f406e44ee84a, /* 1530 */
128'h45850b3006138edd892e9be10079f693, /* 1531 */
128'h00f51e63842a57b5c519cc1ff0ef84aa, /* 1532 */
128'h8526842a86dff0ef852685ca00091c63, /* 1533 */
128'h64e2740270a28522013505a317a010ef, /* 1534 */
128'h28113c23d60101138082614569a26942, /* 1535 */
128'h27313c23292130232891342328813823, /* 1536 */
128'h25713c23276130232751342327413823, /* 1537 */
128'h23b13c2325a130232591342325813823, /* 1538 */
128'hbff7879bbffc07b74d180ac7ed634789, /* 1539 */
128'h8a2e8b3284aabfe787933ffc07b79f3d, /* 1540 */
128'h07e4c68300e7eb630205051300005517, /* 1541 */
128'hf0ef0425051300005517e7b90016f793, /* 1542 */
128'h29013403298130838522f8400413f8ef, /* 1543 */
128'h27013a03278139832801390328813483, /* 1544 */
128'h25013c0325813b8326013b0326813a83, /* 1545 */
128'h2a01011323813d8324013d0324813c83, /* 1546 */
128'hdb4501a50513000055170984a7038082, /* 1547 */
128'h060a8063fe09f99302f109930045aa83, /* 1548 */
128'hcb8902ecf7bb0005ac83e79102eaf7bb, /* 1549 */
128'hb7615429f14ff0ef0185051300005517, /* 1550 */
128'h8c0a009c9c9be3994b8502eadabb54dc, /* 1551 */
128'h280343114e0547818956866200ca0513, /* 1552 */
128'h551700088d6302e878bb0017859b0005, /* 1553 */
128'h4a814c81b7c9ed6ff0ef012505130000, /* 1554 */
128'h020800630116202302e858bbb7f14b81, /* 1555 */
128'h00be17bbcb898b850107c78397d2078e, /* 1556 */
128'h061105210128893b0ffbfb9300fbebb3, /* 1557 */
128'h000055178a89000b8963fa6596e387ae, /* 1558 */
128'hf8aff0ef852685ceee068de3ff450513, /* 1559 */
128'h161b09e9c78309f9c603ee051ae3842a, /* 1560 */
128'h7a63963e09d9c7839e3d0087979b0106, /* 1561 */
128'he50ff0effec505130000551785ca0126, /* 1562 */
128'h89360017f7130a79c683008a4783b5c9, /* 1563 */
128'h47810016e913c3990fe6f9138b89c719, /* 1564 */
128'h579b4b9897d2078e0017861b45914505, /* 1565 */
128'h979b0027571b00c517bbc39d8b850017, /* 1566 */
128'h4189591b4187d79b8b050189191b0187, /* 1567 */
128'hfcb614e387b20ff979130127e933c70d, /* 1568 */
128'h00005517ef898b850a69c78302d90263, /* 1569 */
128'h7933fff7c793b5a92f8020effa450513, /* 1570 */
128'h00005517cb898b8509b9c783bfd100f9, /* 1571 */
128'he20b05e3b535547ddb8ff0effd450513, /* 1572 */
128'h45850af006134685e3958b850af9c783, /* 1573 */
128'hc7830af987a34785e579a21ff0ef8526, /* 1574 */
128'h169b4d914d0108f4aa2300a7979b0e09, /* 1575 */
128'h76130ff6f693f88d061b00dcd6bb003d, /* 1576 */
128'h2d05e9458a2a9edff0ef852645850ff6, /* 1577 */
128'h061b00dad6bb003a169b4c8dfdbd1fe3, /* 1578 */
128'hf0ef852645850ff676130ff6f693f8ca, /* 1579 */
128'h4d6108f00a13ff9a10e32a05e92d9c5f, /* 1580 */
128'h45858656000c26834c818ad209b00d93, /* 1581 */
128'he139999ff0ef85260ff6f6930196d6bb, /* 1582 */
128'h7a132a0dffac90e30ffafa932ca12a85, /* 1583 */
128'h458509c0061386defdba18e30c110ffa, /* 1584 */
128'hc783d4fb0ee34785ed19971ff0ef8526, /* 1585 */
128'h8526458509b00613468501279b630a79, /* 1586 */
128'h45850a70061386cab381842a953ff0ef, /* 1587 */
128'hb325842ab335dd79842a941ff0ef8526, /* 1588 */
128'h00055e63ffdfe0ef842ae406e0221141, /* 1589 */
128'h64028522000307630187b303679c681c, /* 1590 */
128'h80820141640260a245058302014160a2, /* 1591 */
128'h866384aa4791f04af822fc06f4267139, /* 1592 */
128'h10230370079304f592635529478500f5, /* 1593 */
128'h46010107979b4955842e07c4d78300f1, /* 1594 */
128'h4799ed19d44ff0efc43ec24a8526858a, /* 1595 */
128'hc43e478900f41f634791c24a00f11023, /* 1596 */
128'h74a2744270e2d26ff0ef8526858a4601, /* 1597 */
128'hb7cdc402fef414e34785808261217902, /* 1598 */
128'h87ae00d5f3630007869b4f5c6918e215, /* 1599 */
128'h87ba00d5f3630007069b0007859b4f18, /* 1600 */
128'h8082c18ff06f02c50823dd0c0007859b, /* 1601 */
128'hf8a2070d4b9c711910000737691c8082, /* 1602 */
128'hfc5ee0dae4d6e8d2eccef0caf4a6fc86, /* 1603 */
128'hc509f07ff0ef842ac17c8fd9f466f862, /* 1604 */
128'h0000551702042423eb8d6b9c679c681c, /* 1605 */
128'h744670e6f8500493b98ff0efdd450513, /* 1606 */
128'h7be26b066aa66a4669e674a679068526, /* 1607 */
128'hf0eff3e54481541c808261097ca27c42, /* 1608 */
128'h2c2302f4082347851af42c23478df93f, /* 1609 */
128'h409010ef7d000513b8eff0ef85220204, /* 1610 */
128'h2783f94584aa97826b9c679c8522681c, /* 1611 */
128'h478508f422231a04282318042e230884, /* 1612 */
128'hf0ef852245814601b5eff0ef8522d85c, /* 1613 */
128'h00ef8522f14984aacdaff0ef8522f13f, /* 1614 */
128'h8737681c00f1102347a1000505a346d0, /* 1615 */
128'h0aa00713e3991aa007138ff94bdc00ff, /* 1616 */
128'hbe0ff0efc23ec43a8522858a460147d5, /* 1617 */
128'h07b700f715630aa0079300c14703e911, /* 1618 */
128'h0a934a55037009933e900913cc1c8002, /* 1619 */
128'h40000cb780020c3700ff8bb74b050290, /* 1620 */
128'hf0efc402c252013110238522858a4601, /* 1621 */
128'hc25a4bdc015110234c18681ce13db9ef, /* 1622 */
128'hc43e0197e7b301871563c43e0177f7b3, /* 1623 */
128'hca6347b2ed1db76ff0ef8522858a4601, /* 1624 */
128'h319010ef3e80051306090863397d0007, /* 1625 */
128'h8001073700e68563800207374c14bf45, /* 1626 */
128'h06041e23d45c8b8541e7d79bc43ccc18, /* 1627 */
128'h02f51f63f9200793b55d18f40ca34785, /* 1628 */
128'hed09c1cff0ef85224581becff0ef8522, /* 1629 */
128'h4585bfd118f40c2347850007d663443c, /* 1630 */
128'hc505051300005517d965c04ff0ef8522, /* 1631 */
128'h551cb58584aab595fa1004939fcff0ef, /* 1632 */
128'hfed6e352e74eeb4aef26f706f3227161, /* 1633 */
128'he3b54401e6eeeaeaeee6f2e2f6defada, /* 1634 */
128'hc783c7b1199bc7831e7010ef45018baa, /* 1635 */
128'h460104f110234789e7b5180b8ca3198b, /* 1636 */
128'h842aaa2ff0efc482c2be855e008c479d, /* 1637 */
128'h46014495cf818b851b8ba78312050ae3, /* 1638 */
128'h34fd10050de3842aa88ff0ef855e008c, /* 1639 */
128'h842ad99ff0ef855ea031020ba423f4fd, /* 1640 */
128'h6a1a69ba695a64fa741a70ba8522d55d, /* 1641 */
128'h615d6db66d566cf67c167bb67b567af6, /* 1642 */
128'h855e0407c163180b8c23048ba7838082, /* 1643 */
128'h908102051493155010ef4501afeff0ef, /* 1644 */
128'hf155842ab1eff0ef855e45853e800913, /* 1645 */
128'h6fe3131010ef85260007cc63048ba783, /* 1646 */
128'h400007b7bfe91bf010ef0640051308a9, /* 1647 */
128'ha6238b8541e7d79b048ba78300fbac23, /* 1648 */
128'h071b40010737bf0506fb9e23478502fb, /* 1649 */
128'h00ebac234007071b40010737a0292007, /* 1650 */
128'h8b3d5aaa0a1300003a178a1d0036571b, /* 1651 */
128'h45050f8747031086260396529752060a, /* 1652 */
128'ha8238a0500c7d61b02c7073b018ba883, /* 1653 */
128'ha22308eba42304cba823180bae231a0b, /* 1654 */
128'h090ba62300e5183b8b3d0107d71b08eb, /* 1655 */
128'h14070f6302cba703090ba8231408dd63, /* 1656 */
128'h8fd90106d79b8f7d003f07370107979b, /* 1657 */
128'hbc23030787b300d797b32689078546a1, /* 1658 */
128'hbc230c0bb8230c0bb4230c0bb0230a0b, /* 1659 */
128'hd463200007930afbb8230e0bb0230c0b, /* 1660 */
128'hf46320000793090ba70308fba6230107, /* 1661 */
128'h8e63577d04cba783c21508fba82300e7, /* 1662 */
128'h1023855e008c46010107979b471100e7, /* 1663 */
128'h04f11023479d8f6ff0efc282c4be04e1, /* 1664 */
128'h855e008c0107979b4601495507cbd783, /* 1665 */
128'h4785e4051ce3842a8d8ff0efc4bec2ca, /* 1666 */
128'hc94ff0ef855e08fb80a357fd08fbaa23, /* 1667 */
128'h00b54583113000ef855ee40510e3842a, /* 1668 */
128'h018ba703e20515e3842aff3fe0ef855e, /* 1669 */
128'h079304fba0232789100007b754075963, /* 1670 */
128'h979b108c460107cbd78306f110230370, /* 1671 */
128'hd2caed05874ff0efd4bed2ca855e0107, /* 1672 */
128'h988102091a93033007930bf104934905, /* 1673 */
128'h108c08104b210a854991d48206f11023, /* 1674 */
128'h39fdc529844ff0efd05aec56e826855e, /* 1675 */
128'h0737bd8940020737bb75842afe0996e3, /* 1676 */
128'h89bd0165d59bbd9140040737bda94003, /* 1677 */
128'h979b17716705b54508bba82300b515bb, /* 1678 */
128'h00f6d69b17828fd901e6d71b8ff90027, /* 1679 */
128'h0187569b00ff05374098bd798a9d9381, /* 1680 */
128'h0087569b8e698fd50087161b0187179b, /* 1681 */
128'haa2327818fd58ef1f00706138fd16741, /* 1682 */
128'h159b8ecd0187169b0187559b40d804fb, /* 1683 */
128'hac238f558f718ecd0087571b8de90087, /* 1684 */
128'h4689c70109270d638b3d0187d71b04eb, /* 1685 */
128'h02d7971300ebac238001073708d70e63, /* 1686 */
128'ha0238fd920000737040ba78300075963, /* 1687 */
128'h579708f71363800107b7018ba70304fb, /* 1688 */
128'h0ff10c13040ba903639c02a787930000, /* 1689 */
128'h7c933c24849300003497044ba783f0be, /* 1690 */
128'h83f9791302079a93478500f97933fe0c, /* 1691 */
128'h278100f977b300e797bb478540980a85, /* 1692 */
128'hfef493e33a4787930000379704a1ebc5, /* 1693 */
128'hdf400413e15fe0ef8985051300005517, /* 1694 */
128'h03079713b7bda007071b80011737b949, /* 1695 */
128'hbfa980030737b7858002073700074563, /* 1696 */
128'h49959881190201000ab70ff104934905, /* 1697 */
128'h08f1102347990209886339fd09053ac5, /* 1698 */
128'hc556855e010c040007931030c33e47d5, /* 1699 */
128'h4cdce6051de3eb7fe0efdc3ef84af426, /* 1700 */
128'h969bf0070713674144dcfbe18b8583a5, /* 1701 */
128'h50e302e797138fd58ff90087d79b0087, /* 1702 */
128'hbf0104fba0230087e793040ba783f207, /* 1703 */
128'had0340dc840b0b1b06010993017d8b37, /* 1704 */
128'h12078e63278101a7f7b300f977b30009, /* 1705 */
128'h4591200007b700fd0d6345a1400007b7, /* 1706 */
128'h0015b59340bd05b3100005b700fd0863, /* 1707 */
128'h400007370e0519638daa8bfff0ef855e, /* 1708 */
128'h00ed086347912000073700ed0d6347a1, /* 1709 */
128'h02fbaa23001d379340fd0d33100007b7, /* 1710 */
128'h470d00e786634705409cd41fe0ef855e, /* 1711 */
128'hd33e47d50af1102347994d850ae79d63, /* 1712 */
128'h0110d53e00fde7b317c12d81810007b7, /* 1713 */
128'he0efc93ee556e166855e110c04000793, /* 1714 */
128'h409c09b790638bbd010cc783e541dcff, /* 1715 */
128'h0017b79317ed088ba583efd91afba823, /* 1716 */
128'h895ff0ef855e460118fbae2308bba223, /* 1717 */
128'h4601475507cbd7830af1102303700793, /* 1718 */
128'he0efd53ee03ad33a855e110c0107979b, /* 1719 */
128'h0af11023fe0c7d1347b56702ed05d7ff, /* 1720 */
128'h110c0110040007134791d5028dead33a, /* 1721 */
128'hd51fe0efe03ac93ae556e16ae43e855e, /* 1722 */
128'h017d85b74785f3f537fd670267a2c521, /* 1723 */
128'h85934601180bae23096ba2231afba823, /* 1724 */
128'hdef98be310bc099181dff0ef855e8405, /* 1725 */
128'h837902079713f6f762e34581472db575, /* 1726 */
128'h0537040d059366c1bf91118725839752, /* 1727 */
128'h0187d61b0d11000d2783f006869300ff, /* 1728 */
128'h0087d79b8e690087961b8f510187971b, /* 1729 */
128'ha703fda59ee3fefd2e238fd98ff58f51, /* 1730 */
128'ha60300f6f8638bbd00c7579b46a5008d, /* 1731 */
128'h86930000369704d61c63800306b7018b, /* 1732 */
128'hae230087171b1487a78397b6078a0966, /* 1733 */
128'h8ff90186d61b17fd67c100cda68308fb, /* 1734 */
128'hc30503f777130126d71bc78d27818fd1, /* 1735 */
128'h57bb8a8d0106d69b02e6073b3e800613, /* 1736 */
128'ha7830adba2230afba02302d606bb02f7, /* 1737 */
128'h20000793c79919cba7831afbaa231b0b, /* 1738 */
128'h15234a0000ef855e08fba82308fba623, /* 1739 */
128'hd6b7aaaab7b708cba703000506230005, /* 1740 */
128'h27818ef98ff9ccc68693aaa78793cccc, /* 1741 */
128'hf0f0f6b79fb500f037b3068600d036b3, /* 1742 */
128'h06b79fb5068a00d036b38ef90f068693, /* 1743 */
128'h9fb5068e00d036b38ef9f0068693ff01, /* 1744 */
128'h9fb9071200e037338f750207161376c1, /* 1745 */
128'hd70302c7d7b3ed1092010a8bb783d11c, /* 1746 */
128'h0000459784aa06fbc603074bd68307ab, /* 1747 */
128'ha8dfe0effef536230245051357458593, /* 1748 */
128'h0086d79b06cbc603077bc883070ba683, /* 1749 */
128'h0ff777130ff7f7930ff6f8130106d71b, /* 1750 */
128'h04d4851355458593000045970186d69b, /* 1751 */
128'h5505859300004597074ba603a59fe0ef, /* 1752 */
128'h8a3d8abd0146561b0106569b06248513, /* 1753 */
128'h02fba4234785768010ef8526a39fe0ef, /* 1754 */
128'h400407b704fba0232785100007b7b0cd, /* 1755 */
128'hecf769e3400407b700f778631a0bb603, /* 1756 */
128'hb1294c25051300004517e611b5f1e225, /* 1757 */
128'h0c46478304fba0230016879b700006b7, /* 1758 */
128'hf593cd910027f5931abba42303f7f593, /* 1759 */
128'h040ba68304dba0230216869bc58900c7, /* 1760 */
128'h040ba783d7dd8b8504dba0230106e693, /* 1761 */
128'he6f769e3400407b704fba02300c7e793, /* 1762 */
128'hf9b34601088ba583044ba783040ba983, /* 1763 */
128'h849300003497daaff0ef2981855e00f9, /* 1764 */
128'h3c974c2df44b0b1300003b174a85f2e4, /* 1765 */
128'h00f9f7b300fa97bb409cf76c8c930000, /* 1766 */
128'h051300004517ff6498e304a1eb992781, /* 1767 */
128'hf109091300003917bd2197bfe0ef3fe5, /* 1768 */
128'h17ed00494703409c10000db720000d37, /* 1769 */
128'hf7b30009270340dc04f719630017b793, /* 1770 */
128'h0b70061300894683c3a127818ff900f9, /* 1771 */
128'h4681c90ddbbfe0ef855e0fb6f6934585, /* 1772 */
128'h088ba783dabfe0ef855e45850b700613, /* 1773 */
128'h035baa2308fba223180bae231a0ba823, /* 1774 */
128'h2783bfa5fb9910e30931941fe0ef855e, /* 1775 */
128'h8663471100d789634721400006b70009, /* 1776 */
128'h855e02ebaa230017b71341b787b301a7, /* 1777 */
128'h2683f14dfeffe0ef855e408c913fe0ef, /* 1778 */
128'hef8d1afba823409ce79d0046f7930089, /* 1779 */
128'hae2308bba2230017b79317ed088ba583, /* 1780 */
128'h9d9fe0ef855ec9aff0ef855e460118fb, /* 1781 */
128'h855e45850b7006130ff6f693bb35f53d, /* 1782 */
128'h9713fcfc65e34581bfa1d171d13fe0ef, /* 1783 */
128'hfa100413bf6d11872583975283790207, /* 1784 */
128'h6ce000ef06cb851300ec4641ef2ff06f, /* 1785 */
128'h979b008c460107cbd78304f11023478d, /* 1786 */
128'h842a943fe0efc2be47d5855ec4be0107, /* 1787 */
128'h04e157830007d663018ba783ec051163, /* 1788 */
128'hd783c2be479d04f1102347a506fb9e23, /* 1789 */
128'he0efc4be855e0107979b008c460107cb, /* 1790 */
128'h45e646d647c64636e8051763842a90ff, /* 1791 */
128'h06dba22306fba02304cbae23018ba503, /* 1792 */
128'h01a6571bf0e51c634000073706bba423, /* 1793 */
128'h1702ef056863450d0007081b377d8b3d, /* 1794 */
128'h972a4318972a8379ca05051300003517, /* 1795 */
128'h8082557d8082557d80824501c56c8702, /* 1796 */
128'h439cc5e7879300005797808218b50d23, /* 1797 */
128'h00005717842ae406e02247851141ef9d, /* 1798 */
128'h5563ac0fe0ef852212a000efc4f72423, /* 1799 */
128'h13e000ef02c00513fc5ff0ef85220005, /* 1800 */
128'h4501808201414501640260a20dc000ef, /* 1801 */
128'h90636394631cc1670713000057178082, /* 1802 */
128'he406332505130000451785aa114102e7, /* 1803 */
128'ha60380820141853e478160a2f3cfe0ef, /* 1804 */
128'h41488082853ebfd187b600a604630fc7, /* 1805 */
128'h10354703c105fbdff0efe42eec061101, /* 1806 */
128'h0c630ff007930815470302b7006365a2, /* 1807 */
128'h610560e25535e97fe06f610560e200f7, /* 1808 */
128'he4261101bfcdf8400513bfe545018082, /* 1809 */
128'hf0ef842acd09f7dff0ef84aee822ec06, /* 1810 */
128'h64a2644260e2e0800f840413e501ce0f, /* 1811 */
128'h9b87879300005797bfd5553580826105, /* 1812 */
128'h80820f8505138082c3980015071b4388, /* 1813 */
128'h57971101808243889a07879300005797, /* 1814 */
128'h84beec06e4266380e822b4a787930000, /* 1815 */
128'h47838082610564a2644260e200941763, /* 1816 */
128'h5797b7d56000a8cff0ef8522c78119a4, /* 1817 */
128'hab2300005797e79ce39cb1a787930000, /* 1818 */
128'h6798b027879300005797e50880829407, /* 1819 */
128'h5497e4a6711d8082e308e518e11ce788, /* 1820 */
128'hf456f852fc4e6080e8a2aea484930000, /* 1821 */
128'h89aae0caec86e06ae466e862ec5ef05a, /* 1822 */
128'h218a8a9300004a97218a0a1300004a17, /* 1823 */
128'h218b8b9300004b97218b0b1300004b17, /* 1824 */
128'h15634d29794c8c9300003c9700050c1b, /* 1825 */
128'h7aa27a4279e2690664a660e664460294, /* 1826 */
128'h0513000045176d026ca26c426be27b02, /* 1827 */
128'h4c1cc7914901541cdb8fe06f61252d65, /* 1828 */
128'h855a0fc42603681c89560007c3638952, /* 1829 */
128'he0ef855e85ca00090663d9afe0ef638c, /* 1830 */
128'hd80fe0ef856685e200978e63601cd8ef, /* 1831 */
128'h290010ef71c505130000351701a98863, /* 1832 */
128'h4401e04ae426ec06e8221101b7716000, /* 1833 */
128'hcbad511ccbbd4d5ccfad44014d1cc141, /* 1834 */
128'h1c00059384aa892ec7ad639cc7bd651c, /* 1835 */
128'h4799c57c57fdcd21842a166010ef4505, /* 1836 */
128'h03253023e90410f502a347850ef52c23, /* 1837 */
128'h8fa78793fffff797e65ff0ef04052823, /* 1838 */
128'h18f43023224787930000179716f43c23, /* 1839 */
128'h2e23681c18f434232147879300001797, /* 1840 */
128'he99ff0ef10f400230247c78385220ea4, /* 1841 */
128'h106f80826105690264a2644260e28522, /* 1842 */
128'h65186294611c68e68693000046971220, /* 1843 */
128'h0127d713e11897360017671302d786b3, /* 1844 */
128'h17bb40f007bb00f7553b93ed836d8f3d, /* 1845 */
128'h9605051300005517808225018d5d00f7, /* 1846 */
128'h842afefff0efe022e4061141fc3ff06f, /* 1847 */
128'h2501640260a28d410105151bfe9ff0ef, /* 1848 */
128'h041bfdbff0efe022e406114180820141, /* 1849 */
128'h60a28d4115029001fd1ff0ef14020005, /* 1850 */
128'h0785fff5c703058587aa808201416402, /* 1851 */
128'h873300c78c6347818082fb75fee78fa3, /* 1852 */
128'h00e68023078500f506b30007470300f5, /* 1853 */
128'heb09001786930007c70387aa8082f76d, /* 1854 */
128'h8082fb75fee78fa30785fff5c7030585, /* 1855 */
128'h0007c70387b68082e21987aab7d587b6, /* 1856 */
128'h0785fff5c7030585963efb7d00178693, /* 1857 */
128'h808200078023fec799e3d375fee78fa3, /* 1858 */
128'h979b40f707bbfff5c783000547030585, /* 1859 */
128'h8082853ef37d0505e3994187d79b0187, /* 1860 */
128'hc68300e507b3a015478100e614634701, /* 1861 */
128'h979b40f687bb0007c78300e587b30007, /* 1862 */
128'h8082853efee10705e3994187d79b0187, /* 1863 */
128'hc399808200b79363000547830ff5f593, /* 1864 */
128'h000547830ff5f59380824501bfcd0505, /* 1865 */
128'hc70387aabfcd0505dffd808200b79363, /* 1866 */
128'h1101bfcd0785808240a78533e7010007, /* 1867 */
128'h952265a2fe5ff0efec06842ae42ee822, /* 1868 */
128'h7be3157d00b78663000547830ff5f593, /* 1869 */
128'h87aa95aa80826105644260e24501fe85, /* 1870 */
128'h808240a78533e7010007c70300b78563, /* 1871 */
128'hea990007468300f507334781b7fd0785, /* 1872 */
128'hfa7d000746030705fed60ee38082853e, /* 1873 */
128'h468300f507334781bfd5872eb7d50785, /* 1874 */
128'h4603070500d60863a021872eca890007, /* 1875 */
128'h00054703b7c507858082853efa7d0007, /* 1876 */
128'h0007c6830785fee68fe380824501eb19, /* 1877 */
128'he426e8221101bfd587aeb7e50505fafd, /* 1878 */
128'h7607879300004797e519842a84aeec06, /* 1879 */
128'h4783942afa1ff0ef85a68522cc116380, /* 1880 */
128'h852244017407b22300004797ef810004, /* 1881 */
128'hf0ef852285a68082610564a2644260e2, /* 1882 */
128'h050500050023c78100054783c519f9ff, /* 1883 */
128'h6104e4261101bfd970a7bc2300004797, /* 1884 */
128'hc501f73ff0ef8526842ac891e822ec06, /* 1885 */
128'h64a28526644260e2e008050500050023, /* 1886 */
128'hc68387aacf9900054783c11d80826105, /* 1887 */
128'h00e780238082e3110017c703ce810007, /* 1888 */
128'h0075771380824501b7e5078900d780a3, /* 1889 */
128'h8f5537fd07220ff5f69347a1eb0587aa, /* 1890 */
128'hee6340f88833469d00c508b387aaffed, /* 1891 */
128'h97aa078e02e787335761003657930106, /* 1892 */
128'hfee7bc2307a1808200c79763963e963a, /* 1893 */
128'h67b304b50463b7f5feb78fa30785bfe9, /* 1894 */
128'h86b3a811471d4781eb9d872a8b9d00b5, /* 1895 */
128'h0106b02307a100f506b30006b80300f5, /* 1896 */
128'h8733576100365793fed765e340f606b3, /* 1897 */
128'h1363478100f50733963a95be078e02e7, /* 1898 */
128'h00f706b30006c80300f586b3808200f6, /* 1899 */
128'h852e842af0227179b7e5010680230785, /* 1900 */
128'h6622dd3ff0efe02ee84af406e432ec26, /* 1901 */
128'hfff6091300c564636582892ace1184aa, /* 1902 */
128'h70a200040023f75ff0ef944a864a8522, /* 1903 */
128'he02211418082614564e2694285267402, /* 1904 */
128'h60a28522f53ff0ef00a5e963842ae406, /* 1905 */
128'h4781fff6461386ae8832808201416402, /* 1906 */
128'hc58300e685b300f80733fef605e317fd, /* 1907 */
128'h00e614634701b7e500b7002397220005, /* 1908 */
128'h0007c78300e586b300e507b3a8214781, /* 1909 */
128'h962a8082853ed3f59f9507050006c683, /* 1910 */
128'h0505feb78de300054783808200c51363, /* 1911 */
128'hf406e84aec26852e842af0227179bfc5, /* 1912 */
128'h8522c8990005049bd19ff0ef892ee44e, /* 1913 */
128'h0097db63408987bb008509bbd0dff0ef, /* 1914 */
128'h614569a2694264e2740270a285224401, /* 1915 */
128'h0405d17df83ff0ef852285ca86268082, /* 1916 */
128'h8082450100c514630ff5f593962abfe1, /* 1917 */
128'hb7ed853efeb70be30015079300054703, /* 1918 */
128'he60187aa260100c7ef630ff5f59347c1, /* 1919 */
128'h0785feb71ce30007c7038082853e4781, /* 1920 */
128'h083b9f1d4721c39d00757793b7f5367d, /* 1921 */
128'h869b0785fcb69de30007c68387aa00a7, /* 1922 */
128'h97938e19953a93011702fed819e30007, /* 1923 */
128'h020796938fd90107179300b7e7330085, /* 1924 */
128'hd24d8a1deb1187aa27018edd00365713, /* 1925 */
128'hb803bfcd367d0785f8b71fe30007c703, /* 1926 */
128'h12e30007c70300d80a63008785130007, /* 1927 */
128'hb7f1377d87aabfa5fef51be30785f8b7, /* 1928 */
128'h06f71e630300079300054703e7c9419c, /* 1929 */
128'h00e786b305c787930000279700154703, /* 1930 */
128'h0ff777130207071bc6898a850006c683, /* 1931 */
128'hc78397ba0025470304d7176307800693, /* 1932 */
128'h00054703c19c47c1cf950447f7930007, /* 1933 */
128'h000027170015478302f71f6303000793, /* 1934 */
128'h879bc7098b0500074703973e01470713, /* 1935 */
128'h050900e79c63078007130ff7f7930207, /* 1936 */
128'h8fe34741bfed47a98082c19c47a1a809, /* 1937 */
128'hc632ec06006c842ee82211018082fae7, /* 1938 */
128'h081300002817468100c16583f61ff0ef, /* 1939 */
128'h460300f806330007079b00054703fc68, /* 1940 */
128'h644260e2ec0500089863044678930006, /* 1941 */
128'h879b00088b6300467893808261058536, /* 1942 */
128'hb7d196be050502d586b3feb7f4e3fd07, /* 1943 */
128'hfc97879b0ff7f793fe07079bc6098a09, /* 1944 */
128'hf04afc06f426f8227139b7e1e008b7cd, /* 1945 */
128'h65a2b03ff0ef84b2842ae42e00063023, /* 1946 */
128'h80826121790274a2744270e25529e901, /* 1947 */
128'h82e367e2f5dff0ef8522082c892a862e, /* 1948 */
128'hfd279be307858f81cb010007c703fe87, /* 1949 */
128'h00054683b7e94501e088fcf718e347a9, /* 1950 */
128'h05051141f2dff06f00e6846302d00713, /* 1951 */
128'h8082014140a0053360a2f23ff0efe406, /* 1952 */
128'h0693601cf0dff0ef842ee406e0221141, /* 1953 */
128'h069300e6ea6302d704630007c70304b0, /* 1954 */
128'h069380820141640260a202d70e630470, /* 1955 */
128'hc683fed716e306b0069302d7076304d0, /* 1956 */
128'h0027c683fce69fe3052a069007130017, /* 1957 */
128'h052ab7e9e01c078d00e6986304200713, /* 1958 */
128'h006c842ee8221101bfd50789bff1052a, /* 1959 */
128'h2817468100c16583e0dff0efc632ec06, /* 1960 */
128'h06330007079b00054703e72808130000, /* 1961 */
128'hec0500089863044678930006460300f8, /* 1962 */
128'h8b6300467893808261058536644260e2, /* 1963 */
128'h050502d586b3feb7f4e3fd07879b0008, /* 1964 */
128'h0ff7f793fe07079bc6098a09b7d196be, /* 1965 */
128'he406e0221141b7e1e008b7cdfc97879b, /* 1966 */
128'h0007c70304b00693601cf87ff0ef842e, /* 1967 */
128'h02d70e630470069300e6ea6302d70463, /* 1968 */
128'h02d7076304d0069380820141640260a2, /* 1969 */
128'h069007130017c683fed716e306b00693, /* 1970 */
128'h9863042007130027c683fce69fe3052a, /* 1971 */
128'h0789bff1052a052ab7e9e01c078d00e6, /* 1972 */
128'h951ff0efe589842ae406e0221141bfd5, /* 1973 */
128'hd987879300002797fff5c70300a405b3, /* 1974 */
128'h60a2e7198b1100074703973efff58513, /* 1975 */
128'h4703fea47ae3157d80820141557d6402, /* 1976 */
128'h60a26402f77d8b1100074703973e0005, /* 1977 */
128'hf06f4581d7dff06f0141050545814629, /* 1978 */
128'h9141154211418d5d05220085579bfa5f, /* 1979 */
128'he31900054703462946a5478180820141, /* 1980 */
128'h07bb00b6e763fd07059b27018082853e, /* 1981 */
128'he0221141b7c50505fd07879b9fb902f6, /* 1982 */
128'h45a900b7f86347a500a04563842ee406, /* 1983 */
128'h02a4753b4529fe7ff0ef357d02b455bb, /* 1984 */
128'h47854e80006f03050513014160a26402, /* 1985 */
128'h3723000047172cf737230000471707fe, /* 1986 */
128'h2c04041300004417e822110180822cf7, /* 1987 */
128'ha1fff0efec06600885aa84ae862ee426, /* 1988 */
128'h8082610564a26442e00c95a660e2600c, /* 1989 */
128'h000044972947879300004797e4261101, /* 1990 */
128'h35170004b9036380e04ae82228448493, /* 1991 */
128'hd0ef85a24124043bec067b2505130000, /* 1992 */
128'h862286aa608ce41fc0ef85a26088b6ff, /* 1993 */
128'h0000100fb55fd0ef7a85051300003517, /* 1994 */
128'h834a64a260e26442f14025730ff0000f, /* 1995 */
128'h8302610525011fe58593000025976902, /* 1996 */
128'h00850363830fa0ef8432e406e0221141, /* 1997 */
128'h8082450180820141640260a28522547d, /* 1998 */
128'hf606852289aae64e01258413f2227169, /* 1999 */
128'h00a404b30505fa6ff0ef892eea4aee26, /* 2000 */
128'h071beabff0ef95260505f9aff0ef8526, /* 2001 */
128'haf230000479704e7ee631ff00793fff5, /* 2002 */
128'h05130000351784aaf78ff0ef85221aa7, /* 2003 */
128'h04a7f2630ff007939526f6aff0ef5365, /* 2004 */
128'h5185051300003517842af5aff0ef8522, /* 2005 */
128'h6f8505130000351700a405b3f4cff0ef, /* 2006 */
128'h615569b2695264f2741270b2a8dfd0ef, /* 2007 */
128'hb75516f7212300004717200007938082, /* 2008 */
128'h00003597885ff0ef850a458110000613, /* 2009 */
128'h079301294703e10ff0ef850a4d458593, /* 2010 */
128'h850a6ca585930000359700f7096302f0, /* 2011 */
128'h00004797e1cff0ef850a85a2e24ff0ef, /* 2012 */
128'h6b05051300003517858a439011c78793, /* 2013 */
128'h00004717451101f417934405a1dfd0ef, /* 2014 */
128'hdb7ff0ef10f732230000471710f73223, /* 2015 */
128'h4797da9ff0ef4501eea7902300004797, /* 2016 */
128'hec858593000045974611eca79a230000, /* 2017 */
128'hb7990c87932300004797eafff0ef854e, /* 2018 */
128'hdf638432478de04ae426ec06e8221101, /* 2019 */
128'h0004d783d6bff0ef84ae450d892a08c7, /* 2020 */
128'hf0ef096555030000451708a795632501, /* 2021 */
128'hffc4059b06a79a6325010024d783d55f, /* 2022 */
128'h4797d39ff0ef4511dc1ff0ef00448513, /* 2023 */
128'hf0ef0665550300004517e6a791230000, /* 2024 */
128'h00004597e4a79723000047974611d25f, /* 2025 */
128'h256000ef4535e2bff0ef854ae4458593, /* 2026 */
128'h0513d33ff0ef451503c5d58300004597, /* 2027 */
128'hd7830267879300004797240000ef0200, /* 2028 */
128'h0000479700f71c230000471727850007, /* 2029 */
128'h000035170087cf63278d439c00c78793, /* 2030 */
128'h690264a260e26442909fd0ef5bc50513, /* 2031 */
128'h6105690264a2644260e2d5fff06f6105, /* 2032 */
128'h0fa346890105c703f022f40671798082, /* 2033 */
128'h0e6301e1570300e10f230115c70300e1, /* 2034 */
128'h0000351770a2740202f70a63478d00d7, /* 2035 */
128'h00003517842a8b7fd06f614559c50513, /* 2036 */
128'h65a2740285228a7fd0efe42e57450513, /* 2037 */
128'h05c170a241907402d8dff06f614570a2, /* 2038 */
128'h342322813823dc010113ebfff06f6145, /* 2039 */
128'h06134581893284ae842a232130232291, /* 2040 */
128'h061385a6e84ff0ef22113c2300282180, /* 2041 */
128'h8522002cec2ff0efe802c44a08282040, /* 2042 */
128'h228134832301340323813083f63ff0ef, /* 2043 */
128'hd7830000479780822401011322013903, /* 2044 */
128'hf06fd0a58593000045974611cb81f227, /* 2045 */
128'h1041e703492000efe40611418082cf3f, /* 2046 */
128'h10e1a02327051001a70300e57763878e, /* 2047 */
128'h91011782150260a21007e78310a7a223, /* 2048 */
128'he822ec06110180824501808201418d5d, /* 2049 */
128'h07933ce000ef842afc1ff0ef84aae426, /* 2050 */
128'hd533644260e29101150202f407b33e80, /* 2051 */
128'he022e40611418082610564a28d0502a7, /* 2052 */
128'h8793000f47b73a2000ef842af95ff0ef, /* 2053 */
128'h014191011502640260a202f407b32407, /* 2054 */
128'he04ae426e822ec061101808202a7d533, /* 2055 */
128'h02a48533370000ef892af63ff0ef84aa, /* 2056 */
128'h0405944a0285543324040413000f4437, /* 2057 */
128'h690264a2644260e2fe856ee3f45ff0ef, /* 2058 */
128'hec06e822009894b7e426110180826105, /* 2059 */
128'h89260084f363892268048493842ae04a, /* 2060 */
128'h644260e2f47dfa1ff0ef41240433854a, /* 2061 */
128'h4503808200b5002380826105690264a2, /* 2062 */
128'h020575130147c503100007b780820005, /* 2063 */
128'hdfe50207f79301474783100007378082, /* 2064 */
128'h071300078223100007b7808200a70023, /* 2065 */
128'h0007822300e78023476d00e78623f800, /* 2066 */
128'h071300e78423fc70071300e78623470d, /* 2067 */
128'h842ae406e0221141808200e788230200, /* 2068 */
128'hf0ef80820141640260a2e50900044503, /* 2069 */
128'h7713d027879300002797b7f50405fa5f, /* 2070 */
128'h0007c7830007470397aa973e811100f5, /* 2071 */
128'h002ce8221101808200f5802300e580a3, /* 2072 */
128'hf0ef00814503fd1ff0efec068121842a, /* 2073 */
128'h0ff47513002cf5dff0ef00914503f65f, /* 2074 */
128'h00914503f4bff0ef00814503fb7ff0ef, /* 2075 */
128'hf022717980826105644260e2f43ff0ef, /* 2076 */
128'h0089553b54e14461892af406e84aec26, /* 2077 */
128'h346100814503f81ff0ef0ff57513002c, /* 2078 */
128'hfe9410e3f0bff0ef00914503f13ff0ef, /* 2079 */
128'hf022717980826145694264e2740270a2, /* 2080 */
128'h553354e103800413892af406e84aec26, /* 2081 */
128'h00814503f3fff0ef0ff57513002c0089, /* 2082 */
128'h10e3ec9ff0ef00914503ed1ff0ef3461, /* 2083 */
128'h110180826145694264e2740270a2fe94, /* 2084 */
128'hea7ff0ef00814503f13ff0efec06002c, /* 2085 */
128'h100f8082610560e2e9fff0ef00914503, /* 2086 */
128'h000025974305f14025730ff0000f0000, /* 2087 */
128'h35974605d90101138302037ec4458593, /* 2088 */
128'h3423c725051300004517fe2585930000, /* 2089 */
128'h34232521382324913c23268130232611, /* 2090 */
128'h3517c5152501e43fa0ef254130232531, /* 2091 */
128'h340326813083d36fd0ef23a505130000, /* 2092 */
128'h3a032481398325013903258134832601, /* 2093 */
128'h23050513000035178082270101132401, /* 2094 */
128'h080824258593000035974605d0cfd0ef, /* 2095 */
128'h09620bf00913e12d44812501e53fa0ef, /* 2096 */
128'h0074918102049593300a0a1300003a17, /* 2097 */
128'hd41be5052501fbbfa0ef080895ca6605, /* 2098 */
128'h9452dc9ff0ef880d45210004099b00c4, /* 2099 */
128'h47b225a010ef854edbfff0ef00044503, /* 2100 */
128'hc9192501c6efb0ef54020808f3f99cbd, /* 2101 */
128'h051300003517bfb92005051300003517, /* 2102 */
128'h4501efa58593000035974605bf911de5, /* 2103 */
128'h1f05051300003517c5112501d79fa0ef, /* 2104 */
128'h351785a20184961386a20bf00493bf1d, /* 2105 */
128'h051300003517c56fd0ef1f2505130000, /* 2106 */
128'h8d6f90ef0184951385a2c4afd0ef22e5, /* 2107 */
128'h2285051300003517c981c62e0005059b, /* 2108 */
128'hd0ef9fa5051300003517bdddc2cfd0ef, /* 2109 */
128'h25011141900200000023e8dff0efc1ef, /* 2110 */
128'h24050513000f4537a001ddbff0efe406, /* 2111 */
128'h631cafa7071300004717808245018082, /* 2112 */
128'h0513e30895360017869300756513157d, /* 2113 */
128'he822110102b506338082953e055e10d0, /* 2114 */
128'h6622c509842afd1ff0efe4328532ec06, /* 2115 */
128'h80826105644260e285229daff0ef4581, /* 2116 */
128'hd0efe4061c4505130000351711418082, /* 2117 */
128'h0141450160a2f51fc0ef20000537b9ef, /* 2118 */
128'h47a9b000257380824501808245018082, /* 2119 */
128'h85aa862e86b287361141808202f55533, /* 2120 */
128'h4505b62fd0efe4061b05051300003517, /* 2121 */
128'he406952e842ae0221141a001d2dff0ef, /* 2122 */
128'h8d7d640260a29522408007b3f57ff0ef, /* 2123 */
128'h80824505808245058082450580820141, /* 2124 */
128'h186300c684bb842ef406ec26f0227179, /* 2125 */
128'h85b280826145450164e2740270a20096, /* 2126 */
128'h2605200404136622ea3fc0efe4328522, /* 2127 */
128'h8082808245098082450980824509bff9, /* 2128 */
128'hc2dff06f808245018082450180828082, /* 2129 */
128'h84b3003796934781e426e822ec061101, /* 2130 */
128'h64a2644260e200c7986300d5043300d5, /* 2131 */
128'h02e80363609800043803808261054501, /* 2132 */
128'haa0fd0ef12450513000035176090600c, /* 2133 */
128'ha90fd0ef13c505130000351785a28626, /* 2134 */
128'h0000351784aafc26715dbf5d0785a001, /* 2135 */
128'he85aec56f052f44ef84ae0a213c50513, /* 2136 */
128'h00003997a64fd0ef4401892ee45ee486, /* 2137 */
128'h00003b17134a8a9300003a9712c98993, /* 2138 */
128'h00040b9ba44fd0ef854e4a4113cb0b13, /* 2139 */
128'h03271863470187a6a38fd0ef855685de, /* 2140 */
128'h87a6a22fd0ef855a85dea2afd0ef854e, /* 2141 */
128'h00003517fd4417e30405032599634581, /* 2142 */
128'h008706b3a0a94501a08fd0ef16450513, /* 2143 */
128'h07056394e390fff7c613c299863e8a85, /* 2144 */
128'hc31986be8b05639000858733bf6d07a1, /* 2145 */
128'h051300003517058e02d60b63fff7c693, /* 2146 */
128'hd0ef0fa50513000035179cafd0ef0ce5, /* 2147 */
128'h7a0279a2794274e2640660a6557d9bef, /* 2148 */
128'hb75107a10585808261616ba26b426ae2, /* 2149 */
128'heca6020005138aaa6a05fc56e0d27159, /* 2150 */
128'hec66e8caf0a2f486f062f45ef85ae4ce, /* 2151 */
128'h4981bc5ff0ef44818bb28b2ee46ee86a, /* 2152 */
128'h00349793474c0c1300003c179c4a0a13, /* 2153 */
128'h0000351703749b6300fb0cb300fa8db3, /* 2154 */
128'h69a6694670a67406948fd0ef0cc50513, /* 2155 */
128'h85da86266da26d426ce27c027ba26a06, /* 2156 */
128'he0efe47ff06f61657ae285567b4264e6, /* 2157 */
128'h892ac7ffe0ef8d2ac85fe0ef842ac8bf, /* 2158 */
128'h010d1d1b0105151b0344f7b3c79fe0ef, /* 2159 */
128'h8d4191011402150201a4643300a96533, /* 2160 */
128'hb33ff0ef4521ef8100adb02300acb023, /* 2161 */
128'hb23ff0ef0007c50397e20039f7930985, /* 2162 */
128'hf426f822fc06e032e42e7139b7ad0485, /* 2163 */
128'hc1dfe0ef842ac23fe0ef89aaec4ef04a, /* 2164 */
128'h0105151bc11fe0ef84aac17fe0ef892a, /* 2165 */
128'h178265a2660215028fc18d450109179b, /* 2166 */
128'h974e00e588330037971347818d5d9101, /* 2167 */
128'h69e2854e790274a270e2744200c79c63, /* 2168 */
128'he3148ea907856314d8dff06f6121863e, /* 2169 */
128'he42e7139b7f100e830238f2900083703, /* 2170 */
128'he0ef89aaec4ef04af426f822fc06e032, /* 2171 */
128'h84aab9ffe0ef892aba5fe0ef842ababf, /* 2172 */
128'h8fc18d450109179b0105151bb99fe0ef, /* 2173 */
128'h971347818d5d9101178265a266021502, /* 2174 */
128'h70e2744200c79c63974e00e588330037, /* 2175 */
128'hd15ff06f6121863e69e2854e790274a2, /* 2176 */
128'h30238f0900083703e3148e8907856314, /* 2177 */
128'hf426f822fc06e032e42e7139b7f100e8, /* 2178 */
128'hb2dfe0ef842ab33fe0ef89aaec4ef04a, /* 2179 */
128'h0105151bb21fe0ef84aab27fe0ef892a, /* 2180 */
128'h178265a2660215028fc18d450109179b, /* 2181 */
128'h974e00e588330037971347818d5d9101, /* 2182 */
128'h69e2854e790274a270e2744200c79c63, /* 2183 */
128'h02a686b307856314c9dff06f6121863e, /* 2184 */
128'hb7e100e8302302a7073300083703e314, /* 2185 */
128'hec4ef04af426f822fc06e032e42e7139, /* 2186 */
128'he0ef892aab1fe0ef842aab7fe0ef89aa, /* 2187 */
128'h0109179b0105151baa5fe0ef84aaaabf, /* 2188 */
128'h8d5d9101178265a2660215028fc18d45, /* 2189 */
128'h00c79c63974e00e58833003797134781, /* 2190 */
128'h6121863e69e2854e790274a270e27442, /* 2191 */
128'h02a6d6b3078563144505e111c21ff06f, /* 2192 */
128'hb7d100e8302302a7573300083703e314, /* 2193 */
128'hec4ef04af426f822fc06e032e42e7139, /* 2194 */
128'he0ef892aa31fe0ef842aa37fe0ef89aa, /* 2195 */
128'h0109179b0105151ba25fe0ef84aaa2bf, /* 2196 */
128'h8d5d9101178265a2660215028fc18d45, /* 2197 */
128'h00c79c63974e00e58833003797134781, /* 2198 */
128'h6121863e69e2854e790274a270e27442, /* 2199 */
128'h00083703e3148ec907856314ba1ff06f, /* 2200 */
128'hfc06e032e42e7139b7f100e830238f49, /* 2201 */
128'h842a9bffe0ef89aaec4ef04af426f822, /* 2202 */
128'h9adfe0ef84aa9b3fe0ef892a9b9fe0ef, /* 2203 */
128'h660215028fc18d450109179b0105151b, /* 2204 */
128'h88330037971347818d5d9101178265a2, /* 2205 */
128'h790274a270e2744200c79c63974e00e5, /* 2206 */
128'h07856314b29ff06f6121863e69e2854e, /* 2207 */
128'hb7f100e830238f6900083703e3148ee9, /* 2208 */
128'hec4ef04af426f822fc06e032e42e7139, /* 2209 */
128'he0ef892a941fe0ef842a947fe0ef89aa, /* 2210 */
128'h0109179b0105151b935fe0ef84aa93bf, /* 2211 */
128'h8fc59081178265a2660214828fc18cc9, /* 2212 */
128'h00c71c6396ae00d98833003716934701, /* 2213 */
128'h6121863a69e2854e790274a270e27442, /* 2214 */
128'h070500a83023e28800f70533ab1ff06f, /* 2215 */
128'hc305051300003517892ae8ca7159bfc9, /* 2216 */
128'hf486f062f45ef85afc56e0d2e4cef0a2, /* 2217 */
128'h3a17d53fc0ef44018b3289aeec66eca6, /* 2218 */
128'h3c17c22b8b9300003b97c1aa0a130000, /* 2219 */
128'hd31fc0ef855204000a93c2ac0c130000, /* 2220 */
128'h0cb3d23fc0ef8885855e85a2fff44493, /* 2221 */
128'h97ce00f905b30036179314fd46014090, /* 2222 */
128'h856285a2d05fc0efe432855205661863, /* 2223 */
128'h84aaa17ff0ef854a85ce6622cfdfc0ef, /* 2224 */
128'hc385051300003517fb541be32405e129, /* 2225 */
128'h69a664e669468526740670a6cddfc0ef, /* 2226 */
128'h808261656ce27c027ba27b427ae26a06, /* 2227 */
128'h0605e198e3988726c291876600167693, /* 2228 */
128'h0000351784aaeca67159bfc154fdbf59, /* 2229 */
128'hf85afc56e0d2e4cee8caf0a2b5c50513, /* 2230 */
128'h44018ab2892ee86af486ec66f062f45e, /* 2231 */
128'h00003b17b449899300003997c7dfc0ef, /* 2232 */
128'h00003c17e3cb8b9300003b97e3cb0b13, /* 2233 */
128'h04000a13b44c8c9300003c97b3cc0c13, /* 2234 */
128'h000bbd03cba500147793c4bfc0ef854e, /* 2235 */
128'h1793fffd45134601c39fc0ef856285a2, /* 2236 */
128'he432854e05561c6397ca00f485b30036, /* 2237 */
128'h85ca6622c15fc0ef856685a2c1dfc0ef, /* 2238 */
128'hfb441ae32405e5298d2a92fff0ef8526, /* 2239 */
128'h740670a6bf5fc0efb505051300003517, /* 2240 */
128'h7ba27b427ae26a0669a6694664e6856a, /* 2241 */
128'hbf49000b3d03808261656d426ce27c02, /* 2242 */
128'h0605e198e398872ac291876a00167693, /* 2243 */
128'h00003517842ae8a2711db7e15d7db779, /* 2244 */
128'hec5ef05af456f852e0cae4a6a6c50513, /* 2245 */
128'hb91fc0ef4c018ab284aefc4eec86e862, /* 2246 */
128'ha60b0b1300003b17a589091300003917, /* 2247 */
128'hc0ef854a10000a13a68b8b9300003b97, /* 2248 */
128'h1713b63fc0ef855a85ce000c099bb6ff, /* 2249 */
128'h018c17130187e7b38fd9008c1793010c, /* 2250 */
128'h17138fd9028c17138fd9020c17138fd9, /* 2251 */
128'h0036171346018fd9038c17138fd9030c, /* 2252 */
128'hc0efe432854a05561763972600e406b3, /* 2253 */
128'h852285a66622b17fc0ef855e85ceb1ff, /* 2254 */
128'h3517f94c19e30c05e91d89aa831ff0ef, /* 2255 */
128'h854e644660e6af7fc0efa52505130000, /* 2256 */
128'h6c426be27b027aa27a4279e2690664a6, /* 2257 */
128'hbff159fdb74d0605e29ce31c80826125, /* 2258 */
128'hf8a2982505130000351784aaf4a67119, /* 2259 */
128'hf466f862fc5ee0dae4d6e8d2eccef0ca, /* 2260 */
128'haa1fc0ef44018b32892eec6efc86f06a, /* 2261 */
128'h970c8c9300003c97968a0a1300003a17, /* 2262 */
128'h0d1300003d1703f00c13498507f00b93, /* 2263 */
128'h856685a2a75fc0ef855208000a9396ed, /* 2264 */
128'h008995b300e99733408b873ba6dfc0ef, /* 2265 */
128'h05661a6397ca00f486b3003617934601, /* 2266 */
128'ha41fc0ef856a85a2a49fc0efe4328552, /* 2267 */
128'h2405e1398daaf5aff0ef852685ca6622, /* 2268 */
128'ha21fc0ef97c5051300003517fb541be3, /* 2269 */
128'h6aa66a4669e6790674a6856e744670e6, /* 2270 */
128'h808261096de27d027ca27c427be26b06, /* 2271 */
128'he298e398bf610605e28ce38c008c6663, /* 2272 */
128'h0000351784aaf4a67119b7f15dfdbfe5, /* 2273 */
128'he0dae4d6e8d2eccef0caf8a289c50513, /* 2274 */
128'h8b32892eec6efc86f06af466f862fc5e, /* 2275 */
128'h3c97882a0a1300003a179bbfc0ef4401, /* 2276 */
128'h03f00c13498507f00b9388ac8c930000, /* 2277 */
128'hc0ef855208000a93888d0d1300003d17, /* 2278 */
128'h97b3408b87bb987fc0ef856685a298ff, /* 2279 */
128'h4601fff6c693fff7c793008996b300f9, /* 2280 */
128'h855205661a63974a00e485b300361713, /* 2281 */
128'h6622953fc0ef856a85a295bfc0efe432, /* 2282 */
128'h17e32405e1398daae6cff0ef852685ca, /* 2283 */
128'h70e6933fc0ef88e5051300003517fb54, /* 2284 */
128'h6b066aa66a4669e6790674a6856e7446, /* 2285 */
128'h6663808261096de27d027ca27c427be2, /* 2286 */
128'hbfe5e19ce31cbf610605e194e314008c, /* 2287 */
128'h05130000251784aaf4a67119b7f15dfd, /* 2288 */
128'hfc5ee0dae4d6e8d2eccef0caf8a27ae5, /* 2289 */
128'h44018a32892eec6efc86f06af466f862, /* 2290 */
128'h00002c1779498993000029978cdfc0ef, /* 2291 */
128'h0b9308100b134d0507f00a9379cc0c13, /* 2292 */
128'h8a1fc0ef854e796c8c9300002c9703f0, /* 2293 */
128'h408b07bb408a873b899fc0ef856285a2, /* 2294 */
128'h17b30024079b8f5d00ed173300fd17b3, /* 2295 */
128'hfff7c893fff743138fd5008d16b300fd, /* 2296 */
128'h05461c6396ca00d48533003616934601, /* 2297 */
128'h851fc0ef856685a2859fc0efe432854e, /* 2298 */
128'h2405ed298daad6aff0ef852685ca6622, /* 2299 */
128'h7885051300002517f8f41be308000793, /* 2300 */
128'h69e6790674a6856e744670e682dfc0ef, /* 2301 */
128'h6de27d027ca27c427be26b066aa66a46, /* 2302 */
128'h036385be008bea630016781380826109, /* 2303 */
128'h0be385bab7610605e10ce28c85c60008, /* 2304 */
128'h892af0ca7119bf755dfdbfc5859afe08, /* 2305 */
128'hf466fc5ee8d2ecce6985051300002517, /* 2306 */
128'hf862e0dae4d6f4a6f8a2fc86ec6ef06a, /* 2307 */
128'h0a1300002a17fb6fc0ef4b81e03289ae, /* 2308 */
128'h0d1300002d17686c8c9300002c9767ea, /* 2309 */
128'h4401003b949b01779c3347854da168ed, /* 2310 */
128'hc0ef856685da00848b3bf8afc0ef8552, /* 2311 */
128'h08330036171367824601fffc4a93f7ef, /* 2312 */
128'hf60fc0efe432855206f61063974e00e9, /* 2313 */
128'hf0ef854a85ce6622f58fc0ef856a85da, /* 2314 */
128'h2b85fbb41be38c562405e9318b2ac72f, /* 2315 */
128'h6885051300002517fafb90e304000793, /* 2316 */
128'h69e6790674a6855a744670e6f2cfc0ef, /* 2317 */
128'h6de27d027ca27c427be26b066aa66a46, /* 2318 */
128'he30c85d6e11185e20016751380826109, /* 2319 */
128'hfca67175b7e95b7db749060500b83023, /* 2320 */
128'hf0d269850200051384ae892af4cef8ca, /* 2321 */
128'he122e506f86afc66e0e2e4dee8daecd6, /* 2322 */
128'h4b014a098ba6918ff0ef8acae032f46e, /* 2323 */
128'h3d179c4989934ca1018c0c1300003c17, /* 2324 */
128'h96d6003d969367824d819bad0d130000, /* 2325 */
128'h842abb6ff0ef854a85a6866e04fd9663, /* 2326 */
128'h0000251702fa18638aa68bca4785ed4d, /* 2327 */
128'h74e6640a60aa8522e78fc0ef5fc50513, /* 2328 */
128'h7ce26c066ba66b466ae67a0679a67946, /* 2329 */
128'he0efec36b7754a05808261497da27d42, /* 2330 */
128'he42a9aefe0efe82a9b4fe0ef842a9baf, /* 2331 */
128'h161b8d5d0105151b664267a29a8fe0ef, /* 2332 */
128'h37978d4166e29101140215028c510106, /* 2333 */
128'hc683018786b34781e288f6a7bd230000, /* 2334 */
128'h00d600230ff6f693078500fb86330006, /* 2335 */
128'hf0ef4521ef910ba1033df7b3ff9795e3, /* 2336 */
128'hc50397ea8b8d00078b1b001b079b840f, /* 2337 */
128'h7175bfb1547dbf050d8582cff0ef0007, /* 2338 */
128'h69850200051384ae892af4cef8cafca6, /* 2339 */
128'he506f86afc66e0e2e4dee8daecd6f0d2, /* 2340 */
128'h4a098ba6ff7fe0ef8acae032f46ee122, /* 2341 */
128'h9c4989934ca1efec0c1300003c174b01, /* 2342 */
128'h003d969367824d81898d0d1300003d17, /* 2343 */
128'ha94ff0ef854a85a6866e04fd966396d6, /* 2344 */
128'h251702fa18638aa68bca4785ed4d842a, /* 2345 */
128'h640a60aa8522d56fc0ef4da505130000, /* 2346 */
128'h6c066ba66b466ae67a0679a6794674e6, /* 2347 */
128'hec36b7754a05808261497da27d427ce2, /* 2348 */
128'h88cfe0efe82a892fe0ef842a898fe0ef, /* 2349 */
128'h8d5d0105151b664267a2886fe0efe42a, /* 2350 */
128'h8d4166e29101140215028c510106161b, /* 2351 */
128'h018786b34781e288e6a7b02300003797, /* 2352 */
128'h102392c116c2078900fb86330006d683, /* 2353 */
128'h4521ef910ba1033df7b3ff9795e300d6, /* 2354 */
128'h97ea8b8d00078b1b001b079bf1ffe0ef, /* 2355 */
128'hbfb1547dbf050d85f0bfe0ef0007c503, /* 2356 */
128'hf8a2fff5861389b2ecce711980826505, /* 2357 */
128'h05130000251785aa842a892e962af0ca, /* 2358 */
128'hf466f862fc5ee0dae4d6e8d2f4a64165, /* 2359 */
128'h00395793c74fc0efe436fc86ec6ef06a, /* 2360 */
128'h2b9740ab0b1300002b1744854a81e03e, /* 2361 */
128'h2c9740ac0c1300002c1740ab8b930000, /* 2362 */
128'h2d97412d0d1300002d1740ac8c930000, /* 2363 */
128'hf863d7aa0a1300003a17412d8d930000, /* 2364 */
128'h70e6c22fc0ef40650513000025170299, /* 2365 */
128'h6b066aa66a4669e6790674a685567446, /* 2366 */
128'h85a6808261096de27d027ca27c427be2, /* 2367 */
128'hc0ef855e85ce00098663bfafc0ef855a, /* 2368 */
128'hbe0fc0ef856a85e6be8fc0ef8562beef, /* 2369 */
128'hbd0fc0ef856ee129952ff0ef85226582, /* 2370 */
128'hc985000a358302f74c636722010a2783, /* 2371 */
128'h008a3783bb4fc0ef3885051300002517, /* 2372 */
128'h25179782852295a20049561300195593, /* 2373 */
128'h2517b7d14a89b96fc0ef372505130000, /* 2374 */
128'h7179bf890485b86fc0ef0a2505130000, /* 2375 */
128'he84aec26f022f4063605051300002517, /* 2376 */
128'h05130000251704000593cb7fe0efe44e, /* 2377 */
128'hc0ef37a5051300002517b5afc0ef35e5, /* 2378 */
128'h2517b42fc0ef39e5051300002517b4ef, /* 2379 */
128'h99934441b34fc0ef4485052505130000, /* 2380 */
128'h0135853346054685008495b3497901f4, /* 2381 */
128'h64e2740270a2ff2417e3e73ff0ef2405, /* 2382 */
128'h00c5131b460580828082614569a26942, /* 2383 */
128'h081387f245a901f61e13468148814701, /* 2384 */
128'h802397aa0007802397aa000780234000, /* 2385 */
128'hfe0813e397aa387d0007802397aa0007, /* 2386 */
128'hc00026f38e15c020267302b71d632705, /* 2387 */
128'h4000059302a68733411686b33e800513, /* 2388 */
128'h02a7473302a767b302b345bb02c74733, /* 2389 */
128'hfac710e3a94fc06f3385051300002517, /* 2390 */
128'h4501e4061141bf51c00028f3c02026f3, /* 2391 */
128'hf6fff0ef4509f75ff0ef4505f7bff0ef, /* 2392 */
128'hf0ef4541f63ff0ef4521f69ff0ef4511, /* 2393 */
128'h8082e388400007b791011502bff1f5df, /* 2394 */
128'hb823400007b7808225016388400007b7, /* 2395 */
128'h25017b88400007b7808225016b880007, /* 2396 */
128'h07b78d510106161b8d5d0085979b8082, /* 2397 */
128'h0007871b4000063747812581f7884000, /* 2398 */
128'h8b097a98400006b73e80079300b76f63, /* 2399 */
128'h971380827388400007b7ffe537fdc319, /* 2400 */
128'h1141bfc1f61807850007670397360027, /* 2401 */
128'h551b35fd00b7d763842a4785e406e022, /* 2402 */
128'h2a87879300002797883dfedff0ef0045, /* 2403 */
128'hab7fe06f014160a2640200044503943e, /* 2404 */
128'h0810049369054405e0cae4a6e8a2711d, /* 2405 */
128'h09b7047eec5ef05aec86f456f852fc4e, /* 2406 */
128'h079b04e25ae1b0000a373009091380b0, /* 2407 */
128'h87bb0187571b0087979b00f9873b0004, /* 2408 */
128'h4589460100340587e793012767330147, /* 2409 */
128'h458946010034f2dff0efc63ec43a454d, /* 2410 */
128'h00f556b3038007938722f21ff0ef454d, /* 2411 */
128'h18e30421ff579ae3070537e100d70023, /* 2412 */
128'h097e2ca989930000199744014905fa94, /* 2413 */
128'h0a3700100ab7e2eb0b1300002b174bc1, /* 2414 */
128'hc0ef854ef27ff0ef0004051b45a10100, /* 2415 */
128'h45890007c50397ca009407b344818fef, /* 2416 */
128'hff7494e38e4fc0ef854ef0dff0ef0485, /* 2417 */
128'hb43fe0effd4415e38d8fc0ef9456855a, /* 2418 */
128'h7b027aa27a4279e2690664a6644660e6, /* 2419 */
128'he06f2525051300002517808261256be2, /* 2420 */
128'he852ec4ef04af426f822fc0671399fbf, /* 2421 */
128'h19050513000025179b3fe0efe05ae456, /* 2422 */
128'h091300002917400009b744019d9fe0ef, /* 2423 */
128'h0004059b639097ce00341793449518e9, /* 2424 */
128'hdfcf80effe9416e3868fc0ef0405854a, /* 2425 */
128'h2a97400004b7286b0b1300002b174901, /* 2426 */
128'h499117aa0a1300002a1716aa8a930000, /* 2427 */
128'h608ce09c090585560007c783016907b3, /* 2428 */
128'h0004b823824fc0ef8622240125816080, /* 2429 */
128'h7413fd391be3816fc0ef25818552688c, /* 2430 */
128'h0000071702f7646347190054579b0ff4, /* 2431 */
128'h2517878297ba439c97ba078a6a470713, /* 2432 */
128'ha6dfe0ef8522fe7fb0ef13a505130000, /* 2433 */
128'h8522fd3fb0ef1365051300002517a001, /* 2434 */
128'hb0ef1325051300002517b7f5e21ff0ef, /* 2435 */
128'h1305051300002517bfe9c3dff0effbff, /* 2436 */
128'h051300002517b7e1e2af80effadfb0ef, /* 2437 */
128'h00000000bf5dd15ff0eff9bfb0ef12e5, /* 2438 */
128'h00000000000000000000000000000000, /* 2439 */
128'h00000000000000000000000000000000, /* 2440 */
128'h00000000000000000000000000000000, /* 2441 */
128'h00000000000000000000000000000000, /* 2442 */
128'h00000000000000000000000000000000, /* 2443 */
128'h00000000000000000000000000000000, /* 2444 */
128'h00000000000000000000000000000000, /* 2445 */
128'h00000000000000000000000000000000, /* 2446 */
128'h00000000000000000000000000000000, /* 2447 */
128'h08082828282828080808080808080808, /* 2448 */
128'h08080808080808080808080808080808, /* 2449 */
128'h101010101010101010101010101010a0, /* 2450 */
128'h10101010101004040404040404040404, /* 2451 */
128'h01010101010101010141414141414110, /* 2452 */
128'h10101010100101010101010101010101, /* 2453 */
128'h02020202020202020242424242424210, /* 2454 */
128'h08101010100202020202020202020202, /* 2455 */
128'h00000000000000000000000000000000, /* 2456 */
128'h00000000000000000000000000000000, /* 2457 */
128'h101010101010101010101010101010a0, /* 2458 */
128'h10101010101010101010101010101010, /* 2459 */
128'h01010101010101010101010101010101, /* 2460 */
128'h02010101010101011001010101010101, /* 2461 */
128'h02020202020202020202020202020202, /* 2462 */
128'h02020202020202021002020202020202, /* 2463 */
128'hc1bdceee242070dbe8c7b756d76aa478, /* 2464 */
128'hfd469501a83046134787c62af57c0faf, /* 2465 */
128'h895cd7beffff5bb18b44f7af698098d8, /* 2466 */
128'h49b40821a679438efd9871936b901122, /* 2467 */
128'he9b6c7aa265e5a51c040b340f61e2562, /* 2468 */
128'he7d3fbc8d8a1e68102441453d62f105d, /* 2469 */
128'h455a14edf4d50d87c33707d621e1cde6, /* 2470 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /* 2471 */
128'hfde5380c6d9d61228771f681fffa3942, /* 2472 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /* 2473 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /* 2474 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /* 2475 */
128'hfc93a039ab9423a7432aff97f4292244, /* 2476 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /* 2477 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /* 2478 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /* 2479 */
128'h0c07020d08030e09040f0a05000b0601, /* 2480 */
128'h020f0c090603000d0a0704010e0b0805, /* 2481 */
128'h09020b040d060f08010a030c050e0700, /* 2482 */
128'h6c5f7465735f64735f63736972776f6c, /* 2483 */
128'h6e67696c615f64730000000000006465, /* 2484 */
128'h645f6b6c635f64730000000000000000, /* 2485 */
128'h69747465735f64730000000000007669, /* 2486 */
128'h735f646d635f6473000000000000676e, /* 2487 */
128'h74657365725f64730000000074726174, /* 2488 */
128'h6e636b6c625f64730000000000000000, /* 2489 */
128'h69736b6c625f64730000000000000074, /* 2490 */
128'h6f656d69745f6473000000000000657a, /* 2491 */
128'h655f7172695f64730000000000007475, /* 2492 */
128'h5f63736972776f6c000000000000006e, /* 2493 */
128'h00000000646d635f74726174735f6473, /* 2494 */
128'h746e695f746961775f63736972776f6c, /* 2495 */
128'h000000000067616c665f747075727265, /* 2496 */
128'h00007172695f64735f63736972776f6c, /* 2497 */
128'h695f646d635f64735f63736972776f6c, /* 2498 */
128'h5f63736972776f6c0000000000007172, /* 2499 */
128'h007172695f646e655f617461645f6473, /* 2500 */
128'h00000000bffe9c8800000000bffeafc8, /* 2501 */
128'h004c4b40004c4b400030000020000000, /* 2502 */
128'h6d6d5f6472616f62000000020000ffff, /* 2503 */
128'h00000000bffe4ef40064637465675f63, /* 2504 */
128'h00000000bffe4d6200000000bffe4b04, /* 2505 */
128'h00000000000000000000000000000000, /* 2506 */
128'hffffbbdeffffbbdaffffbbdaffffbbb6, /* 2507 */
128'hffffbbe2ffffbbe2ffffbbe2ffffbbe2, /* 2508 */
128'hffffcc04ffffcbfeffffcbf8ffffca54, /* 2509 */
128'h00000000bffeb2f000000000bffeb2e0, /* 2510 */
128'h00000000bffeb31800000000bffeb300, /* 2511 */
128'h00000000bffeb34800000000bffeb330, /* 2512 */
128'h00000000bffeb37800000000bffeb360, /* 2513 */
128'h00000000bffeb3a800000000bffeb390, /* 2514 */
128'h00000000bffeb3d800000000bffeb3c0, /* 2515 */
128'h40040300400402004004010040040000, /* 2516 */
128'h40050000400405004004040140040400, /* 2517 */
128'h30000000000000030000000040050100, /* 2518 */
128'h60000000000000053000000000000001, /* 2519 */
128'h70000000000000027000000000000004, /* 2520 */
128'h00000001400000007000000000000000, /* 2521 */
128'h00000005000000012000000000000006, /* 2522 */
128'h20000000000000020000000040000000, /* 2523 */
128'h00000000100000000000000100000000, /* 2524 */
128'h1e19140f0d0c0a000000000000000000, /* 2525 */
128'h000186a00000271050463c37322d2823, /* 2526 */
128'h017d7840017d784000989680000f4240, /* 2527 */
128'h031975000319750002faf080018cba80, /* 2528 */
128'h02faf08005f5e10002faf080017d7840, /* 2529 */
128'h00000020000000000bebc2000c65d400, /* 2530 */
128'h00000200000001000000008000000040, /* 2531 */
128'h00002000000010000000080000000400, /* 2532 */
128'h0000c000000080000000600000004000, /* 2533 */
128'h37363534333231300002000000010000, /* 2534 */
128'h2043534952776f4c4645444342413938, /* 2535 */
128'h746f6f622d7520646573696d696e696d, /* 2536 */
128'h00000000647261432d445320726f6620, /* 2537 */
128'hfffff980fffff996fffff982fffff96e, /* 2538 */
128'h00000000fffff9bafffff980fffff9a8, /* 2539 */
128'he00600003800000039080000edfe0dd0, /* 2540 */
128'h00000000100000001100000028000000, /* 2541 */
128'h0000000000000000a806000059010000, /* 2542 */
128'h00000000010000000000000000000000, /* 2543 */
128'h02000000000000000400000003000000, /* 2544 */
128'h020000000f0000000400000003000000, /* 2545 */
128'h2c6874651b0000001400000003000000, /* 2546 */
128'h007665642d657261622d656e61697261, /* 2547 */
128'h2c687465260000001000000003000000, /* 2548 */
128'h0100000000657261622d656e61697261, /* 2549 */
128'h1a0000000300000000006e65736f6863, /* 2550 */
128'h303140747261752f636f732f2c000000, /* 2551 */
128'h0000003030323531313a303030303030, /* 2552 */
128'h00000000737570630100000002000000, /* 2553 */
128'h01000000000000000400000003000000, /* 2554 */
128'h000000000f0000000400000003000000, /* 2555 */
128'h40787d01380000000400000003000000, /* 2556 */
128'h03000000000000304075706301000000, /* 2557 */
128'h0300000080f0fa024b00000004000000, /* 2558 */
128'h03000000007570635b00000004000000, /* 2559 */
128'h03000000000000006700000004000000, /* 2560 */
128'h0000000079616b6f6b00000005000000, /* 2561 */
128'h7a6874651b0000001300000003000000, /* 2562 */
128'h0000766373697200656e61697261202c, /* 2563 */
128'h34367672720000000b00000003000000, /* 2564 */
128'h0b000000030000000000636466616d69, /* 2565 */
128'h0000393376732c76637369727c000000, /* 2566 */
128'h01000000850000000000000003000000, /* 2567 */
128'h6f72746e6f632d747075727265746e69, /* 2568 */
128'h04000000030000000000000072656c6c, /* 2569 */
128'h0000000003000000010000008f000000, /* 2570 */
128'h1b0000000f00000003000000a0000000, /* 2571 */
128'h000063746e692d7570632c7663736972, /* 2572 */
128'h01000000b50000000400000003000000, /* 2573 */
128'h01000000bb0000000400000003000000, /* 2574 */
128'h01000000020000000200000002000000, /* 2575 */
128'h0030303030303030384079726f6d656d, /* 2576 */
128'h6f6d656d5b0000000700000003000000, /* 2577 */
128'h67000000100000000300000000007972, /* 2578 */
128'h00000040000000000000008000000000, /* 2579 */
128'h0300000000636f730100000002000000, /* 2580 */
128'h03000000020000000000000004000000, /* 2581 */
128'h03000000020000000f00000004000000, /* 2582 */
128'h616972612c6874651b0000001f000000, /* 2583 */
128'h706d697300636f732d657261622d656e, /* 2584 */
128'h000000000300000000007375622d656c, /* 2585 */
128'h303240746e696c6301000000c3000000, /* 2586 */
128'h0d000000030000000000003030303030, /* 2587 */
128'h30746e696c632c76637369721b000000, /* 2588 */
128'hca000000100000000300000000000000, /* 2589 */
128'h07000000010000000300000001000000, /* 2590 */
128'h00000000670000001000000003000000, /* 2591 */
128'h0300000000000c000000000000000002, /* 2592 */
128'h006c6f72746e6f63de00000008000000, /* 2593 */
128'h7075727265746e690100000002000000, /* 2594 */
128'h3030634072656c6c6f72746e6f632d74, /* 2595 */
128'h04000000030000000000000030303030, /* 2596 */
128'h04000000030000000000000000000000, /* 2597 */
128'h0c00000003000000010000008f000000, /* 2598 */
128'h003063696c702c76637369721b000000, /* 2599 */
128'h03000000a00000000000000003000000, /* 2600 */
128'h0b00000001000000ca00000010000000, /* 2601 */
128'h10000000030000000900000001000000, /* 2602 */
128'h000000000000000c0000000067000000, /* 2603 */
128'he8000000040000000300000000000004, /* 2604 */
128'hfb000000040000000300000007000000, /* 2605 */
128'hb5000000040000000300000003000000, /* 2606 */
128'hbb000000040000000300000002000000, /* 2607 */
128'h75626564010000000200000002000000, /* 2608 */
128'h0000304072656c6c6f72746e6f632d67, /* 2609 */
128'h637369721b0000001000000003000000, /* 2610 */
128'h03000000003331302d67756265642c76, /* 2611 */
128'hffff000001000000ca00000008000000, /* 2612 */
128'h00000000670000001000000003000000, /* 2613 */
128'h03000000001000000000000000000000, /* 2614 */
128'h006c6f72746e6f63de00000008000000, /* 2615 */
128'h30303140747261750100000002000000, /* 2616 */
128'h08000000030000000000003030303030, /* 2617 */
128'h03000000003035373631736e1b000000, /* 2618 */
128'h00000010000000006700000010000000, /* 2619 */
128'h04000000030000000010000000000000, /* 2620 */
128'h040000000300000080f0fa024b000000, /* 2621 */
128'h040000000300000000c2010006010000, /* 2622 */
128'h04000000030000000200000014010000, /* 2623 */
128'h04000000030000000100000025010000, /* 2624 */
128'h04000000030000000200000030010000, /* 2625 */
128'h0100000002000000040000003a010000, /* 2626 */
128'h3030303240636d6d2d63736972776f6c, /* 2627 */
128'h10000000030000000000000030303030, /* 2628 */
128'h00000000000000200000000067000000, /* 2629 */
128'h14010000040000000300000000000100, /* 2630 */
128'h25010000040000000300000002000000, /* 2631 */
128'h1b0000000c0000000300000002000000, /* 2632 */
128'h0200000000636d6d2d63736972776f6c, /* 2633 */
128'h406874652d63736972776f6c01000000, /* 2634 */
128'h03000000000000003030303030303033, /* 2635 */
128'h2d63736972776f6c1b0000000c000000, /* 2636 */
128'h5b000000080000000300000000687465, /* 2637 */
128'h0400000003000000006b726f7774656e, /* 2638 */
128'h04000000030000000200000014010000, /* 2639 */
128'h06000000030000000300000025010000, /* 2640 */
128'h0300000000007fe3023e180047010000, /* 2641 */
128'h00000030000000006700000010000000, /* 2642 */
128'h01000000020000000080000000000000, /* 2643 */
128'h303440646e7277682d63736972776f6c, /* 2644 */
128'h0e000000030000000000303030303030, /* 2645 */
128'h6e7277682d63736972776f6c1b000000, /* 2646 */
128'h67000000100000000300000000000064, /* 2647 */
128'h00100000000000000000004000000000, /* 2648 */
128'h09000000020000000200000002000000, /* 2649 */
128'h2300736c6c65632d7373657264646123, /* 2650 */
128'h61706d6f6300736c6c65632d657a6973, /* 2651 */
128'h6f647473006c65646f6d00656c626974, /* 2652 */
128'h65736162656d697400687461702d7475, /* 2653 */
128'h6b636f6c630079636e6575716572662d, /* 2654 */
128'h63697665640079636e6575716572662d, /* 2655 */
128'h75746174730067657200657079745f65, /* 2656 */
128'h2d756d6d006173692c76637369720073, /* 2657 */
128'h230074696c70732d626c740065707974, /* 2658 */
128'h00736c6c65632d747075727265746e69, /* 2659 */
128'h6f72746e6f632d747075727265746e69, /* 2660 */
128'h646e6168702c78756e696c0072656c6c, /* 2661 */
128'h727265746e69007365676e617200656c, /* 2662 */
128'h6572006465646e657478652d73747075, /* 2663 */
128'h616d2c76637369720073656d616e2d67, /* 2664 */
128'h766373697200797469726f6972702d78, /* 2665 */
128'h70732d746e6572727563007665646e2c, /* 2666 */
128'h61702d747075727265746e6900646565, /* 2667 */
128'h0073747075727265746e6900746e6572, /* 2668 */
128'h6f692d6765720074666968732d676572, /* 2669 */
128'h63616d2d6c61636f6c0068746469772d, /* 2670 */
128'h0000000000000000737365726464612d, /* 2671 */
128'h0000000000203a642520656369766544, /* 2672 */
128'h00203a6425206563697665642073250a, /* 2673 */
128'h00000000203a6425206563697665440a, /* 2674 */
128'h000a656369766564206e776f6e6b6e75, /* 2675 */
128'h00000a2973252c73252870756b6f6f6c, /* 2676 */
128'h7265206c616e7265746e692070636864, /* 2677 */
128'h00000000000000000a7025202c726f72, /* 2678 */
128'h5145525f5043484420676e69646e6553, /* 2679 */
128'h4b434120504348440000000a54534555, /* 2680 */
128'h696c432050434844000000000000000a, /* 2681 */
128'h203a7373657264644120504920746e65, /* 2682 */
128'h0000000a64252e64252e64252e642520, /* 2683 */
128'h73657264644120504920726576726553, /* 2684 */
128'h0a64252e64252e64252e642520203a73, /* 2685 */
128'h6120726574756f520000000000000000, /* 2686 */
128'h252e64252e642520203a737365726464, /* 2687 */
128'h6b73616d2074654e0000000a64252e64, /* 2688 */
128'h64252e642520203a7373657264646120, /* 2689 */
128'h697420657361654c000a64252e64252e, /* 2690 */
128'h7364253a6d64253a686425203d20656d, /* 2691 */
128'h3d206e69616d6f44000000000000000a, /* 2692 */
128'h4820746e65696c4300000a2273252220, /* 2693 */
128'h000a22732522203d20656d616e74736f, /* 2694 */
128'h000000000a44455050494b53204b4341, /* 2695 */
128'h000000000000000a4b414e2050434844, /* 2696 */
128'h73657264646120646574736575716552, /* 2697 */
128'h0000000000000a646573756665722073, /* 2698 */
128'h000000000000000a732520726f727245, /* 2699 */
128'h6e6f6974706f2064656c646e61686e75, /* 2700 */
128'h656c646e61686e55000000000a642520, /* 2701 */
128'h64252065646f63706f20504348442064, /* 2702 */
128'h20676e69646e6553000000000000000a, /* 2703 */
128'h000a595245564f435349445f50434844, /* 2704 */
128'h00000000000a29732528726f72726570, /* 2705 */
128'h3a2043414d2073250000000030687465, /* 2706 */
128'h3a583230253a583230253a5832302520, /* 2707 */
128'h000a583230253a583230253a58323025, /* 2708 */
128'h484420646e65732074276e646c756f43, /* 2709 */
128'h206e6f20595245564f43534944205043, /* 2710 */
128'h00000a7325203a732520656369766564, /* 2711 */
128'h5043484420726f6620676e6974696157, /* 2712 */
128'h2020202020202020000a524546464f5f, /* 2713 */
128'h00000000000063250000000000000020, /* 2714 */
128'h0000005832302520000000000000002e, /* 2715 */
128'h00000000732573250000000000000a0a, /* 2716 */
128'h00000000007325203a646c697542202c, /* 2717 */
128'h73257a4820756c250000000000007325, /* 2718 */
128'h0000000000756c250000000000000000, /* 2719 */
128'h0073257a4863252000000000646c252e, /* 2720 */
128'h00000000007325736574794220756c25, /* 2721 */
128'h00003a786c3830250073254269632520, /* 2722 */
128'h000a73252020202000786c6c2a302520, /* 2723 */
128'h000000203a5d64255b6e6f6974636553, /* 2724 */
128'h25203d206465726975716572206e656c, /* 2725 */
128'h000a7825203d206c6175746361202c58, /* 2726 */
128'h302c782578302c7825287970636d656d, /* 2727 */
128'h25287465736d656d00000a3b29782578, /* 2728 */
128'h00000000000a3b29782578302c302c78, /* 2729 */
128'h0000000054455346464f5f4f4c43414d, /* 2730 */
128'h0000000054455346464f5f494843414d, /* 2731 */
128'h000000000054455346464f5f524c5054, /* 2732 */
128'h000000000054455346464f5f53434654, /* 2733 */
128'h0054455346464f5f4c5254434f49444d, /* 2734 */
128'h000000000054455346464f5f53434652, /* 2735 */
128'h00000000000054455346464f5f525352, /* 2736 */
128'h000000000054455346464f5f44414252, /* 2737 */
128'h000000000054455346464f5f524c5052, /* 2738 */
128'h46464f5f524c5052000000003f3f3f3f, /* 2739 */
128'h0000000000000047000064252b544553, /* 2740 */
128'h0a50495049203d206f746f7250205049, /* 2741 */
128'h00000000000000540000000000000000, /* 2742 */
128'h000a504745203d206f746f7250205049, /* 2743 */
128'h000a505550203d206f746f7250205049, /* 2744 */
128'h0000000a3a7265646165682074736574, /* 2745 */
128'h000a3a73746e65746e6f632074736574, /* 2746 */
128'h000a504449203d206f746f7250205049, /* 2747 */
128'h00000a5054203d206f746f7250205049, /* 2748 */
128'h0a50434344203d206f746f7250205049, /* 2749 */
128'h00000000000000360000000000000000, /* 2750 */
128'h0a50565352203d206f746f7250205049, /* 2751 */
128'h6f746f72502050490000000000000000, /* 2752 */
128'h6f746f7250205049000a455247203d20, /* 2753 */
128'h6f746f7250205049000a505345203d20, /* 2754 */
128'h6f746f725020504900000a4841203d20, /* 2755 */
128'h6f746f7250205049000a50544d203d20, /* 2756 */
128'h0000000000000a485054454542203d20, /* 2757 */
128'h5041434e45203d206f746f7250205049, /* 2758 */
128'h000000000000004d000000000000000a, /* 2759 */
128'h0a504d4f43203d206f746f7250205049, /* 2760 */
128'h6f746f72502050490000000000000000, /* 2761 */
128'h00000000000000000a50544353203d20, /* 2762 */
128'h494c504455203d206f746f7250205049, /* 2763 */
128'h6f746f725020504900000000000a4554, /* 2764 */
128'h00000000000000000a534c504d203d20, /* 2765 */
128'h000a574152203d206f746f7250205049, /* 2766 */
128'h7075736e75203d206f746f7270205049, /* 2767 */
128'h000000000a2978252820646574726f70, /* 2768 */
128'h257830203d20657079745f6f746f7270, /* 2769 */
128'h656c646e61686e750000000000000a78, /* 2770 */
128'h0000000a21747075727265746e692064, /* 2771 */
128'h000a726464612043414d207075746553, /* 2772 */
128'h25203d205d64255b4d454f2049505351, /* 2773 */
128'h6c25203d2043414d0000000000000a78, /* 2774 */
128'h726464612043414d00000a786c253a78, /* 2775 */
128'h3a783230253a78323025203d20737365, /* 2776 */
128'h253a783230253a783230253a78323025, /* 2777 */
128'h74656e72656874450000000a2e783230, /* 2778 */
128'h757461747320747075727265746e6920, /* 2779 */
128'h00000000000000000a646c25203d2073, /* 2780 */
128'h20646564616f6c2065687420746f6f42, /* 2781 */
128'h00000000000a2e2e2e6d6172676f7270, /* 2782 */
128'h207265746f6f62202c657962646f6f47, /* 2783 */
128'h3d3c3b3a2c2b2a22000000000a2e2e2e, /* 2784 */
128'h3c3b3a2e2c2b2a2200007f7c5d5b3f3e, /* 2785 */
128'h3736353433323130007f7c5d5b3f3e3d, /* 2786 */
128'h00000000000000006665646362613938, /* 2787 */
128'h2e636d6d5f63736972776f6c2f637273, /* 2788 */
128'h20657361625f64730000000000000063, /* 2789 */
128'h00726464615f657361625f6473203d3d, /* 2790 */
128'h74207325203a64735f63736972776f6c, /* 2791 */
128'h6d65722064726143000a74756f656d69, /* 2792 */
128'h676e616863206b73616d202c6465766f, /* 2793 */
128'h000000000000000a6425206f74206465, /* 2794 */
128'h6d202c6465747265736e692064726143, /* 2795 */
128'h25206f74206465676e616863206b7361, /* 2796 */
128'h6165726320636d6d0000000000000a64, /* 2797 */
128'h2074736f68202c782520746120646574, /* 2798 */
128'h00000000007365590000000a7825203d, /* 2799 */
128'h00000000524444200000000000006f4e, /* 2800 */
128'h203a656369766544002020203a434d4d, /* 2801 */
128'h74636166756e614d00000000000a7325, /* 2802 */
128'h000000000a7825203a44492072657275, /* 2803 */
128'h00000000000000000a7825203a4d454f, /* 2804 */
128'h63256325632563256325203a656d614e, /* 2805 */
128'h65657053207375420000000000000a20, /* 2806 */
128'h706143206867694800000a6425203a64, /* 2807 */
128'h0000000000000a7325203a7974696361, /* 2808 */
128'h000000000000203a7974696361706143, /* 2809 */
128'h69622d6425203a687464695720737542, /* 2810 */
128'h000000203a78250a000000000a732574, /* 2811 */
128'h5f63736972776f6c0000007825782520, /* 2812 */
128'h206e776f6e6b6e550000000000006473, /* 2813 */
128'h45207375746174530000000065646f6d, /* 2814 */
128'h0000000a583830257830203a726f7272, /* 2815 */
128'h20676e69746961772074756f656d6954, /* 2816 */
128'h00000000000a79646165722064726163, /* 2817 */
128'h646e6573206f74206c69616620636d6d, /* 2818 */
128'h0000000000000a646d6320706f747320, /* 2819 */
128'h65626d756e206b636f6c62203a434d4d, /* 2820 */
128'h207364656563786520786c2578302072, /* 2821 */
128'h00000000000a29786c2578302878616d, /* 2822 */
128'h7571657220342e34203d3e20434d4d65, /* 2823 */
128'h65636e61686e6520726f662064657269, /* 2824 */
128'h61657261206174616420726573752064, /* 2825 */
128'h656f642064726143000000000000000a, /* 2826 */
128'h61702074726f7070757320746f6e2073, /* 2827 */
128'h00000000000a676e696e6f6974697472, /* 2828 */
128'h656420746f6e2073656f642064726143, /* 2829 */
128'h70756f726720505720434820656e6966, /* 2830 */
128'h746164207265735500000a657a697320, /* 2831 */
128'h2061657261206465636e61686e652061, /* 2832 */
128'h2070756f726720505720434820746f6e, /* 2833 */
128'h0000000a64656e67696c6120657a6973, /* 2834 */
128'h6e206e6f697469747261702069255047, /* 2835 */
128'h732070756f726720505720434820746f, /* 2836 */
128'h000000000a64656e67696c6120657a69, /* 2837 */
128'h757320746f6e2073656f642064726143, /* 2838 */
128'h61206465636e61686e652074726f7070, /* 2839 */
128'h000000000000000a6574756269727474, /* 2840 */
128'h73206465636e61686e65206c61746f54, /* 2841 */
128'h6978616d207364656563786520657a69, /* 2842 */
128'h00000a297525203e20752528206d756d, /* 2843 */
128'h757320746f6e2073656f642064726143, /* 2844 */
128'h72746e6f632074736f682074726f7070, /* 2845 */
128'h206e6f697469747261702064656c6c6f, /* 2846 */
128'h74696c696261696c6572206574697277, /* 2847 */
128'h00000000000a73676e69747465732079, /* 2848 */
128'h7261702079646165726c612064726143, /* 2849 */
128'h000000000000000a64656e6f69746974, /* 2850 */
128'h6572702064726163206f6e203a434d4d, /* 2851 */
128'h64696420647261430000000a746e6573, /* 2852 */
128'h206f7420646e6f7073657220746f6e20, /* 2853 */
128'h0a217463656c657320656761746c6f76, /* 2854 */
128'h7420656c62616e750000000000000000, /* 2855 */
128'h0a65646f6d2061207463656c6573206f, /* 2856 */
128'h635f747865206f4e0000000000000000, /* 2857 */
128'h0000000000000a21646e756f66206473, /* 2858 */
128'h34302520726e532078363025206e614d, /* 2859 */
128'h63256325632563250000007834302578, /* 2860 */
128'h00000064252e64250000000063256325, /* 2861 */
128'h00000000000079636167656c20434d4d, /* 2862 */
128'h0000000000000079636167654c204453, /* 2863 */
128'h28206465657053206867694820434d4d, /* 2864 */
128'h20686769482044530000297a484d3632, /* 2865 */
128'h000000297a484d303528206465657053, /* 2866 */
128'h28206465657053206867694820434d4d, /* 2867 */
128'h3552444420434d4d0000297a484d3235, /* 2868 */
128'h00000000000000297a484d3235282032, /* 2869 */
128'h7a484d35322820323152445320534855, /* 2870 */
128'h32524453205348550000000000000029, /* 2871 */
128'h00000000000000297a484d3035282035, /* 2872 */
128'h484d3030312820303552445320534855, /* 2873 */
128'h3552444420534855000000000000297a, /* 2874 */
128'h00000000000000297a484d3035282030, /* 2875 */
128'h4d383032282034303152445320534855, /* 2876 */
128'h32282030303253480000000000297a48, /* 2877 */
128'h6976654420434d4d0000297a484d3030, /* 2878 */
128'h0a646e756f6620746f6e206425206563, /* 2879 */
128'h00000000000044530000000000000000, /* 2880 */
128'h00006425203a732500000000434d4d65, /* 2881 */
128'h0000000000636d6d0000002973252820, /* 2882 */
128'h6425203d206874676e656c20656c6946, /* 2883 */
128'h252c70252835646d000000000000000a, /* 2884 */
128'h00000000000000000a7325203d202964, /* 2885 */
128'h6f6f7420687461702074736575716552, /* 2886 */
128'h00000000000a646c25202e676e6f6c20, /* 2887 */
128'h732522203a717277000000000000002f, /* 2888 */
128'h0a64253d657a69736b636f6c62202c22, /* 2889 */
128'h20657669656365520000000000000000, /* 2890 */
128'h0000000000000a2e646e6520656c6966, /* 2891 */
128'h656c6c6163207172775f656c646e6168, /* 2892 */
128'h206c6167656c6c4900000000000a2e64, /* 2893 */
128'h0a2e6e6f6974617265706f2050544654, /* 2894 */
128'h206f74206c6961460000000000000000, /* 2895 */
128'h2172657669726420445320746e756f6d, /* 2896 */
128'h6f6f622064616f4c000000000000000a, /* 2897 */
128'h726f6d656d206f746e69206e69622e74, /* 2898 */
128'h6e69622e746f6f620000000000000a79, /* 2899 */
128'h742064656c6961460000000000000000, /* 2900 */
128'h0000000a21746f6f62206e65706f206f, /* 2901 */
128'h69662065736f6c63206f74206c696166, /* 2902 */
128'h206f74206c696166000000000021656c, /* 2903 */
128'h00000000216b73696420746e756f6d75, /* 2904 */
128'h20736574796220642520646564616f4c, /* 2905 */
128'h7365726464612079726f6d656d206f74, /* 2906 */
128'h622e746f6f62206d6f72662078252073, /* 2907 */
128'h0a2e736574796220642520666f206e69, /* 2908 */
128'h666c652064616f6c0000000000000000, /* 2909 */
128'h000a79726f6d656d20524444206f7420, /* 2910 */
128'h2064656c696166206461657220666c65, /* 2911 */
128'h0000000064252065646f632068746977, /* 2912 */
128'h20746f6f622d750a000000005c2d2f7c, /* 2913 */
128'h67617473207473726966206465736162, /* 2914 */
128'h00000a726564616f6c20746f6f622065, /* 2915 */
128'h696166207325206e6f69747265737361, /* 2916 */
128'h696c202c732520656c6966202c64656c, /* 2917 */
128'h206e6f6974636e7566202c642520656e, /* 2918 */
128'h3a4552554c49414600000000000a7325, /* 2919 */
128'h74612078257830203d21207825783020, /* 2920 */
128'h00000a2e782578302074657366666f20, /* 2921 */
128'h7025203d203270202c7025203d203170, /* 2922 */
128'h2020202020202020000000000000000a, /* 2923 */
128'h08080808080808080000000000202020, /* 2924 */
128'h20676e69747465730000000000080808, /* 2925 */
128'h20676e69747365740000000000007525, /* 2926 */
128'h3a4552554c4941460000000000007525, /* 2927 */
128'h64612064616220656c626973736f7020, /* 2928 */
128'h666f20746120656e696c207373657264, /* 2929 */
128'h00000000000a2e782578302074657366, /* 2930 */
128'h7478656e206f7420676e697070696b53, /* 2931 */
128'h000000000000000a2e2e2e7473657420, /* 2932 */
128'h20202020200808080808080808080808, /* 2933 */
128'h08080808080808080808202020202020, /* 2934 */
128'h00000000000820080000000000000008, /* 2935 */
128'h78302073692065676e61722074736574, /* 2936 */
128'h00000000000a70257830206f74207025, /* 2937 */
128'h000000000075252f00752520706f6f4c, /* 2938 */
128'h6441206b637574530000000000000a3a, /* 2939 */
128'h0000203a732520200000007373657264, /* 2940 */
128'h00000a2e656e6f4400000000000a6b6f, /* 2941 */
128'h4d415244206c6174656d20657261420a, /* 2942 */
128'h65747365746d656d00000a7473657420, /* 2943 */
128'h20302e332e34206e6f69737265762072, /* 2944 */
128'h000000000000000a297469622d642528, /* 2945 */
128'h30322029432820746867697279706f43, /* 2946 */
128'h2073656c7261684320323130322d3130, /* 2947 */
128'h000000000000000a2e6e6f62617a6143, /* 2948 */
128'h74207265646e75206465736e6563694c, /* 2949 */
128'h50206c6172656e654720554e47206568, /* 2950 */
128'h65762065736e6563694c2063696c6275, /* 2951 */
128'h0a2e29796c6e6f282032206e6f697372, /* 2952 */
128'h5f676e696b726f770000000000000000, /* 2953 */
128'h20646c25202c424b6425203d20746573, /* 2954 */
128'h6c25202c736e6f697463757274736e69, /* 2955 */
128'h203d20495043202c73656c6379632064, /* 2956 */
128'h00000000000000000a646c252e646c25, /* 2957 */
128'h46454443424139383736353433323130, /* 2958 */
128'h6f57206f6c6c65480000000000000000, /* 2959 */
128'h205d64255b70777300000a0d21646c72, /* 2960 */
128'h73206863746977530000000a5825203d, /* 2961 */
128'h000a58252c5825203d20676e69747465, /* 2962 */
128'h5825203d2064656573206d6f646e6152, /* 2963 */
128'h0a746f6f62204453000000000000000a, /* 2964 */
128'h6f6f6220495053510000000000000000, /* 2965 */
128'h736574204d4152440000000000000a74, /* 2966 */
128'h6f6f6220505446540000000000000a74, /* 2967 */
128'h65742065686361430000000000000a74, /* 2968 */
128'h00000a0d7061727400000000000a7473, /* 2969 */
128'hefcdab8967452301cccccccccccccccd, /* 2970 */
128'h10000000200000001032547698badcfe, /* 2971 */
128'h55555555555555555851f42d4c957f2d, /* 2972 */
128'h000000030f060301aaaaaaaaaaaaaaaa, /* 2973 */
128'h00000000004b4d4700004b4d47545045, /* 2974 */
128'h00000000000000000000000030000000, /* 2975 */
128'h000000000c00000000000000ffffffff, /* 2976 */
128'h00006772615f64730000646d635f6473, /* 2977 */
128'h00000000cc33aa5500000000bffeb270, /* 2978 */
128'h00000000000000000000000000000000, /* 2979 */
128'h00000000000000000000000000000000, /* 2980 */
128'h00000000000000000000000000000000, /* 2981 */
128'h00000000000000000000000000000000, /* 2982 */
128'h00000000000000000000000000000000, /* 2983 */
128'h00000000000000000000000000000000, /* 2984 */
128'h00000000000000000000000000000000, /* 2985 */
128'h00000000000000000000000000000000, /* 2986 */
128'h00000000000000000000000000000000, /* 2987 */
128'h00000000000000000000000000000000, /* 2988 */
128'h00000000000000000000000000000000, /* 2989 */
128'h00000000000000000000000000000000, /* 2990 */
128'h00000000000000000000000000000000, /* 2991 */
128'h000000002f7c5c2d00000000ffffffff, /* 2992 */
128'hffffffff0000000600000000bffeb428, /* 2993 */
128'h00000000bffe711c0000000000000000, /* 2994 */
128'h000000000000000000000000000000de, /* 2995 */
128'h00000000000000000000000000000000, /* 2996 */
128'h00000000000000000000000000000000, /* 2997 */
128'h00000000000000000000000000000000, /* 2998 */
128'h00000000000000000000000000000000, /* 2999 */
128'h00000000000000000000000000000000, /* 3000 */
128'h00000000000000000000000000000000, /* 3001 */
128'h00000000000000000000000000000000, /* 3002 */
128'h00000000000000000000000000000000, /* 3003 */
128'h00000000000000000000000000000000, /* 3004 */
128'h00000000000000000000000000000000, /* 3005 */
128'h00000000000000000000000000000000, /* 3006 */
128'h00000000000000000000000000000000, /* 3007 */
128'h00000000000000000000000000000000, /* 3008 */
128'h00000000000000000000000000000000, /* 3009 */
128'h00000000000000000000000000000000, /* 3010 */
128'h00000000000000000000000000000000, /* 3011 */
128'h00000000000000000000000000000000, /* 3012 */
128'h00000000000000000000000000000000, /* 3013 */
128'h00000000000000000000000000000000, /* 3014 */
128'h00000000000000000000000000000000, /* 3015 */
128'h00000000000000000000000000000000, /* 3016 */
128'h00000000000000000000000000000000, /* 3017 */
128'h00000000000000000000000000000000, /* 3018 */
128'h00000000000000000000000000000000, /* 3019 */
128'h00000000000000000000000000000000, /* 3020 */
128'h00000000000000000000000000000000, /* 3021 */
128'h00000000000000000000000000000000, /* 3022 */
128'h00000000000000000000000000000000, /* 3023 */
128'h00000000000000000000000000000000, /* 3024 */
128'h00000000000000000000000000000000, /* 3025 */
128'h00000000000000000000000000000000, /* 3026 */
128'h00000000000000000000000000000000, /* 3027 */
128'h00000000000000000000000000000000, /* 3028 */
128'h00000000000000000000000000000000, /* 3029 */
128'h00000000000000000000000000000000, /* 3030 */
128'h00000000000000000000000000000000, /* 3031 */
128'h00000000000000000000000000000000, /* 3032 */
128'h00000000000000000000000000000000, /* 3033 */
128'h00000000000000000000000000000000, /* 3034 */
128'h00000000000000000000000000000000, /* 3035 */
128'h00000000000000000000000000000000, /* 3036 */
128'h00000000000000000000000000000000, /* 3037 */
128'h00000000000000000000000000000000, /* 3038 */
128'h00000000000000000000000000000000, /* 3039 */
128'h00000000000000000000000000000000, /* 3040 */
128'h00000000000000000000000000000000, /* 3041 */
128'h00000000000000000000000000000000, /* 3042 */
128'h00000000000000000000000000000000, /* 3043 */
128'h00000000000000000000000000000000, /* 3044 */
128'h00000000000000000000000000000000, /* 3045 */
128'h00000000000000000000000000000000, /* 3046 */
128'h00000000000000000000000000000000, /* 3047 */
128'h00000000000000000000000000000000, /* 3048 */
128'h00000000000000000000000000000000, /* 3049 */
128'h00000000000000000000000000000000, /* 3050 */
128'h00000000000000000000000000000000, /* 3051 */
128'h00000000000000000000000000000000, /* 3052 */
128'h00000000000000000000000000000000, /* 3053 */
128'h00000000000000000000000000000000, /* 3054 */
128'h00000000000000000000000000000000, /* 3055 */
128'h00000000000000000000000000000000, /* 3056 */
128'h00000000000000000000000000000000, /* 3057 */
128'h00000000000000000000000000000000, /* 3058 */
128'h00000000000000000000000000000000, /* 3059 */
128'h00000000000000000000000000000000, /* 3060 */
128'h00000000000000000000000000000000, /* 3061 */
128'h00000000000000000000000000000000, /* 3062 */
128'h00000000000000000000000000000000, /* 3063 */
128'h00000000000000000000000000000000, /* 3064 */
128'h00000000000000000000000000000000, /* 3065 */
128'h00000000000000000000000000000000, /* 3066 */
128'h00000000000000000000000000000000, /* 3067 */
128'h00000000000000000000000000000000, /* 3068 */
128'h00000000000000000000000000000000, /* 3069 */
128'h00000000000000000000000000000000, /* 3070 */
128'h00000000000000000000000000000000, /* 3071 */
128'h00000000000000000000000000000000, /* 3072 */
128'h00000000000000000000000000000000, /* 3073 */
128'h00000000000000000000000000000000, /* 3074 */
128'h00000000000000000000000000000000, /* 3075 */
128'h00000000000000000000000000000000, /* 3076 */
128'h00000000000000000000000000000000, /* 3077 */
128'h00000000000000000000000000000000, /* 3078 */
128'h00000000000000000000000000000000, /* 3079 */
128'h00000000000000000000000000000000, /* 3080 */
128'h00000000000000000000000000000000, /* 3081 */
128'h00000000000000000000000000000000, /* 3082 */
128'h00000000000000000000000000000000, /* 3083 */
128'h00000000000000000000000000000000, /* 3084 */
128'h00000000000000000000000000000000, /* 3085 */
128'h00000000000000000000000000000000, /* 3086 */
128'h00000000000000000000000000000000, /* 3087 */
128'h00000000000000000000000000000000, /* 3088 */
128'h00000000000000000000000000000000, /* 3089 */
128'h00000000000000000000000000000000, /* 3090 */
128'h00000000000000000000000000000000, /* 3091 */
128'h00000000000000000000000000000000, /* 3092 */
128'h00000000000000000000000000000000, /* 3093 */
128'h00000000000000000000000000000000, /* 3094 */
128'h00000000000000000000000000000000, /* 3095 */
128'h00000000000000000000000000000000, /* 3096 */
128'h00000000000000000000000000000000, /* 3097 */
128'h00000000000000000000000000000000, /* 3098 */
128'h00000000000000000000000000000000, /* 3099 */
128'h00000000000000000000000000000000, /* 3100 */
128'h00000000000000000000000000000000, /* 3101 */
128'h00000000000000000000000000000000, /* 3102 */
128'h00000000000000000000000000000000, /* 3103 */
128'h00000000000000000000000000000000, /* 3104 */
128'h00000000000000000000000000000000, /* 3105 */
128'h00000000000000000000000000000000, /* 3106 */
128'h00000000000000000000000000000000, /* 3107 */
128'h00000000000000000000000000000000, /* 3108 */
128'h00000000000000000000000000000000, /* 3109 */
128'h00000000000000000000000000000000, /* 3110 */
128'h00000000000000000000000000000000, /* 3111 */
128'h00000000000000000000000000000000, /* 3112 */
128'h00000000000000000000000000000000, /* 3113 */
128'h00000000000000000000000000000000, /* 3114 */
128'h00000000000000000000000000000000, /* 3115 */
128'h00000000000000000000000000000000, /* 3116 */
128'h00000000000000000000000000000000, /* 3117 */
128'h00000000000000000000000000000000, /* 3118 */
128'h00000000000000000000000000000000, /* 3119 */
128'h00000000000000000000000000000000, /* 3120 */
128'h00000000000000000000000000000000, /* 3121 */
128'h00000000000000000000000000000000, /* 3122 */
128'h00000000000000000000000000000000, /* 3123 */
128'h00000000000000000000000000000000, /* 3124 */
128'h00000000000000000000000000000000, /* 3125 */
128'h00000000000000000000000000000000, /* 3126 */
128'h00000000000000000000000000000000, /* 3127 */
128'h00000000000000000000000000000000, /* 3128 */
128'h00000000000000000000000000000000, /* 3129 */
128'h00000000000000000000000000000000, /* 3130 */
128'h00000000000000000000000000000000, /* 3131 */
128'h00000000000000000000000000000000, /* 3132 */
128'h00000000000000000000000000000000, /* 3133 */
128'h00000000000000000000000000000000, /* 3134 */
128'h00000000000000000000000000000000, /* 3135 */
128'h00000000000000000000000000000000, /* 3136 */
128'h00000000000000000000000000000000, /* 3137 */
128'h00000000000000000000000000000000, /* 3138 */
128'h00000000000000000000000000000000, /* 3139 */
128'h00000000000000000000000000000000, /* 3140 */
128'h00000000000000000000000000000000, /* 3141 */
128'h00000000000000000000000000000000, /* 3142 */
128'h00000000000000000000000000000000, /* 3143 */
128'h00000000000000000000000000000000, /* 3144 */
128'h00000000000000000000000000000000, /* 3145 */
128'h00000000000000000000000000000000, /* 3146 */
128'h00000000000000000000000000000000, /* 3147 */
128'h00000000000000000000000000000000, /* 3148 */
128'h00000000000000000000000000000000, /* 3149 */
128'h00000000000000000000000000000000, /* 3150 */
128'h00000000000000000000000000000000, /* 3151 */
128'h00000000000000000000000000000000, /* 3152 */
128'h00000000000000000000000000000000, /* 3153 */
128'h00000000000000000000000000000000, /* 3154 */
128'h00000000000000000000000000000000, /* 3155 */
128'h00000000000000000000000000000000, /* 3156 */
128'h00000000000000000000000000000000, /* 3157 */
128'h00000000000000000000000000000000, /* 3158 */
128'h00000000000000000000000000000000, /* 3159 */
128'h00000000000000000000000000000000, /* 3160 */
128'h00000000000000000000000000000000, /* 3161 */
128'h00000000000000000000000000000000, /* 3162 */
128'h00000000000000000000000000000000, /* 3163 */
128'h00000000000000000000000000000000, /* 3164 */
128'h00000000000000000000000000000000, /* 3165 */
128'h00000000000000000000000000000000, /* 3166 */
128'h00000000000000000000000000000000, /* 3167 */
128'h00000000000000000000000000000000, /* 3168 */
128'h00000000000000000000000000000000, /* 3169 */
128'h00000000000000000000000000000000, /* 3170 */
128'h00000000000000000000000000000000, /* 3171 */
128'h00000000000000000000000000000000, /* 3172 */
128'h00000000000000000000000000000000, /* 3173 */
128'h00000000000000000000000000000000, /* 3174 */
128'h00000000000000000000000000000000, /* 3175 */
128'h00000000000000000000000000000000, /* 3176 */
128'h00000000000000000000000000000000, /* 3177 */
128'h00000000000000000000000000000000, /* 3178 */
128'h00000000000000000000000000000000, /* 3179 */
128'h00000000000000000000000000000000, /* 3180 */
128'h00000000000000000000000000000000, /* 3181 */
128'h00000000000000000000000000000000, /* 3182 */
128'h00000000000000000000000000000000, /* 3183 */
128'h00000000000000000000000000000000, /* 3184 */
128'h00000000000000000000000000000000, /* 3185 */
128'h00000000000000000000000000000000, /* 3186 */
128'h00000000000000000000000000000000, /* 3187 */
128'h00000000000000000000000000000000, /* 3188 */
128'h00000000000000000000000000000000, /* 3189 */
128'h00000000000000000000000000000000, /* 3190 */
128'h00000000000000000000000000000000, /* 3191 */
128'h00000000000000000000000000000000, /* 3192 */
128'h00000000000000000000000000000000, /* 3193 */
128'h00000000000000000000000000000000, /* 3194 */
128'h00000000000000000000000000000000, /* 3195 */
128'h00000000000000000000000000000000, /* 3196 */
128'h00000000000000000000000000000000, /* 3197 */
128'h00000000000000000000000000000000, /* 3198 */
128'h00000000000000000000000000000000, /* 3199 */
128'h00000000000000000000000000000000, /* 3200 */
128'h00000000000000000000000000000000, /* 3201 */
128'h00000000000000000000000000000000, /* 3202 */
128'h00000000000000000000000000000000, /* 3203 */
128'h00000000000000000000000000000000, /* 3204 */
128'h00000000000000000000000000000000, /* 3205 */
128'h00000000000000000000000000000000, /* 3206 */
128'h00000000000000000000000000000000, /* 3207 */
128'h00000000000000000000000000000000, /* 3208 */
128'h00000000000000000000000000000000, /* 3209 */
128'h00000000000000000000000000000000, /* 3210 */
128'h00000000000000000000000000000000, /* 3211 */
128'h00000000000000000000000000000000, /* 3212 */
128'h00000000000000000000000000000000, /* 3213 */
128'h00000000000000000000000000000000, /* 3214 */
128'h00000000000000000000000000000000, /* 3215 */
128'h00000000000000000000000000000000, /* 3216 */
128'h00000000000000000000000000000000, /* 3217 */
128'h00000000000000000000000000000000, /* 3218 */
128'h00000000000000000000000000000000, /* 3219 */
128'h00000000000000000000000000000000, /* 3220 */
128'h00000000000000000000000000000000, /* 3221 */
128'h00000000000000000000000000000000, /* 3222 */
128'h00000000000000000000000000000000, /* 3223 */
128'h00000000000000000000000000000000, /* 3224 */
128'h00000000000000000000000000000000, /* 3225 */
128'h00000000000000000000000000000000, /* 3226 */
128'h00000000000000000000000000000000, /* 3227 */
128'h00000000000000000000000000000000, /* 3228 */
128'h00000000000000000000000000000000, /* 3229 */
128'h00000000000000000000000000000000, /* 3230 */
128'h00000000000000000000000000000000, /* 3231 */
128'h00000000000000000000000000000000, /* 3232 */
128'h00000000000000000000000000000000, /* 3233 */
128'h00000000000000000000000000000000, /* 3234 */
128'h00000000000000000000000000000000, /* 3235 */
128'h00000000000000000000000000000000, /* 3236 */
128'h00000000000000000000000000000000, /* 3237 */
128'h00000000000000000000000000000000, /* 3238 */
128'h00000000000000000000000000000000, /* 3239 */
128'h00000000000000000000000000000000, /* 3240 */
128'h00000000000000000000000000000000, /* 3241 */
128'h00000000000000000000000000000000, /* 3242 */
128'h00000000000000000000000000000000, /* 3243 */
128'h00000000000000000000000000000000, /* 3244 */
128'h00000000000000000000000000000000, /* 3245 */
128'h00000000000000000000000000000000, /* 3246 */
128'h00000000000000000000000000000000, /* 3247 */
128'h00000000000000000000000000000000, /* 3248 */
128'h00000000000000000000000000000000, /* 3249 */
128'h00000000000000000000000000000000, /* 3250 */
128'h00000000000000000000000000000000, /* 3251 */
128'h00000000000000000000000000000000, /* 3252 */
128'h00000000000000000000000000000000, /* 3253 */
128'h00000000000000000000000000000000, /* 3254 */
128'h00000000000000000000000000000000, /* 3255 */
128'h00000000000000000000000000000000, /* 3256 */
128'h00000000000000000000000000000000, /* 3257 */
128'h00000000000000000000000000000000, /* 3258 */
128'h00000000000000000000000000000000, /* 3259 */
128'h00000000000000000000000000000000, /* 3260 */
128'h00000000000000000000000000000000, /* 3261 */
128'h00000000000000000000000000000000, /* 3262 */
128'h00000000000000000000000000000000, /* 3263 */
128'h00000000000000000000000000000000, /* 3264 */
128'h00000000000000000000000000000000, /* 3265 */
128'h00000000000000000000000000000000, /* 3266 */
128'h00000000000000000000000000000000, /* 3267 */
128'h00000000000000000000000000000000, /* 3268 */
128'h00000000000000000000000000000000, /* 3269 */
128'h00000000000000000000000000000000, /* 3270 */
128'h00000000000000000000000000000000, /* 3271 */
128'h00000000000000000000000000000000, /* 3272 */
128'h00000000000000000000000000000000, /* 3273 */
128'h00000000000000000000000000000000, /* 3274 */
128'h00000000000000000000000000000000, /* 3275 */
128'h00000000000000000000000000000000, /* 3276 */
128'h00000000000000000000000000000000, /* 3277 */
128'h00000000000000000000000000000000, /* 3278 */
128'h00000000000000000000000000000000, /* 3279 */
128'h00000000000000000000000000000000, /* 3280 */
128'h00000000000000000000000000000000, /* 3281 */
128'h00000000000000000000000000000000, /* 3282 */
128'h00000000000000000000000000000000, /* 3283 */
128'h00000000000000000000000000000000, /* 3284 */
128'h00000000000000000000000000000000, /* 3285 */
128'h00000000000000000000000000000000, /* 3286 */
128'h00000000000000000000000000000000, /* 3287 */
128'h00000000000000000000000000000000, /* 3288 */
128'h00000000000000000000000000000000, /* 3289 */
128'h00000000000000000000000000000000, /* 3290 */
128'h00000000000000000000000000000000, /* 3291 */
128'h00000000000000000000000000000000, /* 3292 */
128'h00000000000000000000000000000000, /* 3293 */
128'h00000000000000000000000000000000, /* 3294 */
128'h00000000000000000000000000000000, /* 3295 */
128'h00000000000000000000000000000000, /* 3296 */
128'h00000000000000000000000000000000, /* 3297 */
128'h00000000000000000000000000000000, /* 3298 */
128'h00000000000000000000000000000000, /* 3299 */
128'h00000000000000000000000000000000, /* 3300 */
128'h00000000000000000000000000000000, /* 3301 */
128'h00000000000000000000000000000000, /* 3302 */
128'h00000000000000000000000000000000, /* 3303 */
128'h00000000000000000000000000000000, /* 3304 */
128'h00000000000000000000000000000000, /* 3305 */
128'h00000000000000000000000000000000, /* 3306 */
128'h00000000000000000000000000000000, /* 3307 */
128'h00000000000000000000000000000000, /* 3308 */
128'h00000000000000000000000000000000, /* 3309 */
128'h00000000000000000000000000000000, /* 3310 */
128'h00000000000000000000000000000000, /* 3311 */
128'h00000000000000000000000000000000, /* 3312 */
128'h00000000000000000000000000000000, /* 3313 */
128'h00000000000000000000000000000000, /* 3314 */
128'h00000000000000000000000000000000, /* 3315 */
128'h00000000000000000000000000000000, /* 3316 */
128'h00000000000000000000000000000000, /* 3317 */
128'h00000000000000000000000000000000, /* 3318 */
128'h00000000000000000000000000000000, /* 3319 */
128'h00000000000000000000000000000000, /* 3320 */
128'h00000000000000000000000000000000, /* 3321 */
128'h00000000000000000000000000000000, /* 3322 */
128'h00000000000000000000000000000000, /* 3323 */
128'h00000000000000000000000000000000, /* 3324 */
128'h00000000000000000000000000000000, /* 3325 */
128'h00000000000000000000000000000000, /* 3326 */
128'h00000000000000000000000000000000, /* 3327 */
128'h00000000000000000000000000000000, /* 3328 */
128'h00000000000000000000000000000000, /* 3329 */
128'h00000000000000000000000000000000, /* 3330 */
128'h00000000000000000000000000000000, /* 3331 */
128'h00000000000000000000000000000000, /* 3332 */
128'h00000000000000000000000000000000, /* 3333 */
128'h00000000000000000000000000000000, /* 3334 */
128'h00000000000000000000000000000000, /* 3335 */
128'h00000000000000000000000000000000, /* 3336 */
128'h00000000000000000000000000000000, /* 3337 */
128'h00000000000000000000000000000000, /* 3338 */
128'h00000000000000000000000000000000, /* 3339 */
128'h00000000000000000000000000000000, /* 3340 */
128'h00000000000000000000000000000000, /* 3341 */
128'h00000000000000000000000000000000, /* 3342 */
128'h00000000000000000000000000000000, /* 3343 */
128'h00000000000000000000000000000000, /* 3344 */
128'h00000000000000000000000000000000, /* 3345 */
128'h00000000000000000000000000000000, /* 3346 */
128'h00000000000000000000000000000000, /* 3347 */
128'h00000000000000000000000000000000, /* 3348 */
128'h00000000000000000000000000000000, /* 3349 */
128'h00000000000000000000000000000000, /* 3350 */
128'h00000000000000000000000000000000, /* 3351 */
128'h00000000000000000000000000000000, /* 3352 */
128'h00000000000000000000000000000000, /* 3353 */
128'h00000000000000000000000000000000, /* 3354 */
128'h00000000000000000000000000000000, /* 3355 */
128'h00000000000000000000000000000000, /* 3356 */
128'h00000000000000000000000000000000, /* 3357 */
128'h00000000000000000000000000000000, /* 3358 */
128'h00000000000000000000000000000000, /* 3359 */
128'h00000000000000000000000000000000, /* 3360 */
128'h00000000000000000000000000000000, /* 3361 */
128'h00000000000000000000000000000000, /* 3362 */
128'h00000000000000000000000000000000, /* 3363 */
128'h00000000000000000000000000000000, /* 3364 */
128'h00000000000000000000000000000000, /* 3365 */
128'h00000000000000000000000000000000, /* 3366 */
128'h00000000000000000000000000000000, /* 3367 */
128'h00000000000000000000000000000000, /* 3368 */
128'h00000000000000000000000000000000, /* 3369 */
128'h00000000000000000000000000000000, /* 3370 */
128'h00000000000000000000000000000000, /* 3371 */
128'h00000000000000000000000000000000, /* 3372 */
128'h00000000000000000000000000000000, /* 3373 */
128'h00000000000000000000000000000000, /* 3374 */
128'h00000000000000000000000000000000, /* 3375 */
128'h00000000000000000000000000000000, /* 3376 */
128'h00000000000000000000000000000000, /* 3377 */
128'h00000000000000000000000000000000, /* 3378 */
128'h00000000000000000000000000000000, /* 3379 */
128'h00000000000000000000000000000000, /* 3380 */
128'h00000000000000000000000000000000, /* 3381 */
128'h00000000000000000000000000000000, /* 3382 */
128'h00000000000000000000000000000000, /* 3383 */
128'h00000000000000000000000000000000, /* 3384 */
128'h00000000000000000000000000000000, /* 3385 */
128'h00000000000000000000000000000000, /* 3386 */
128'h00000000000000000000000000000000, /* 3387 */
128'h00000000000000000000000000000000, /* 3388 */
128'h00000000000000000000000000000000, /* 3389 */
128'h00000000000000000000000000000000, /* 3390 */
128'h00000000000000000000000000000000, /* 3391 */
128'h00000000000000000000000000000000, /* 3392 */
128'h00000000000000000000000000000000, /* 3393 */
128'h00000000000000000000000000000000, /* 3394 */
128'h00000000000000000000000000000000, /* 3395 */
128'h00000000000000000000000000000000, /* 3396 */
128'h00000000000000000000000000000000, /* 3397 */
128'h00000000000000000000000000000000, /* 3398 */
128'h00000000000000000000000000000000, /* 3399 */
128'h00000000000000000000000000000000, /* 3400 */
128'h00000000000000000000000000000000, /* 3401 */
128'h00000000000000000000000000000000, /* 3402 */
128'h00000000000000000000000000000000, /* 3403 */
128'h00000000000000000000000000000000, /* 3404 */
128'h00000000000000000000000000000000, /* 3405 */
128'h00000000000000000000000000000000, /* 3406 */
128'h00000000000000000000000000000000, /* 3407 */
128'h00000000000000000000000000000000, /* 3408 */
128'h00000000000000000000000000000000, /* 3409 */
128'h00000000000000000000000000000000, /* 3410 */
128'h00000000000000000000000000000000, /* 3411 */
128'h00000000000000000000000000000000, /* 3412 */
128'h00000000000000000000000000000000, /* 3413 */
128'h00000000000000000000000000000000, /* 3414 */
128'h00000000000000000000000000000000, /* 3415 */
128'h00000000000000000000000000000000, /* 3416 */
128'h00000000000000000000000000000000, /* 3417 */
128'h00000000000000000000000000000000, /* 3418 */
128'h00000000000000000000000000000000, /* 3419 */
128'h00000000000000000000000000000000, /* 3420 */
128'h00000000000000000000000000000000, /* 3421 */
128'h00000000000000000000000000000000, /* 3422 */
128'h00000000000000000000000000000000, /* 3423 */
128'h00000000000000000000000000000000, /* 3424 */
128'h00000000000000000000000000000000, /* 3425 */
128'h00000000000000000000000000000000, /* 3426 */
128'h00000000000000000000000000000000, /* 3427 */
128'h00000000000000000000000000000000, /* 3428 */
128'h00000000000000000000000000000000, /* 3429 */
128'h00000000000000000000000000000000, /* 3430 */
128'h00000000000000000000000000000000, /* 3431 */
128'h00000000000000000000000000000000, /* 3432 */
128'h00000000000000000000000000000000, /* 3433 */
128'h00000000000000000000000000000000, /* 3434 */
128'h00000000000000000000000000000000, /* 3435 */
128'h00000000000000000000000000000000, /* 3436 */
128'h00000000000000000000000000000000, /* 3437 */
128'h00000000000000000000000000000000, /* 3438 */
128'h00000000000000000000000000000000, /* 3439 */
128'h00000000000000000000000000000000, /* 3440 */
128'h00000000000000000000000000000000, /* 3441 */
128'h00000000000000000000000000000000, /* 3442 */
128'h00000000000000000000000000000000, /* 3443 */
128'h00000000000000000000000000000000, /* 3444 */
128'h00000000000000000000000000000000, /* 3445 */
128'h00000000000000000000000000000000, /* 3446 */
128'h00000000000000000000000000000000, /* 3447 */
128'h00000000000000000000000000000000, /* 3448 */
128'h00000000000000000000000000000000, /* 3449 */
128'h00000000000000000000000000000000, /* 3450 */
128'h00000000000000000000000000000000, /* 3451 */
128'h00000000000000000000000000000000, /* 3452 */
128'h00000000000000000000000000000000, /* 3453 */
128'h00000000000000000000000000000000, /* 3454 */
128'h00000000000000000000000000000000, /* 3455 */
128'h00000000000000000000000000000000, /* 3456 */
128'h00000000000000000000000000000000, /* 3457 */
128'h00000000000000000000000000000000, /* 3458 */
128'h00000000000000000000000000000000, /* 3459 */
128'h00000000000000000000000000000000, /* 3460 */
128'h00000000000000000000000000000000, /* 3461 */
128'h00000000000000000000000000000000, /* 3462 */
128'h00000000000000000000000000000000, /* 3463 */
128'h00000000000000000000000000000000, /* 3464 */
128'h00000000000000000000000000000000, /* 3465 */
128'h00000000000000000000000000000000, /* 3466 */
128'h00000000000000000000000000000000, /* 3467 */
128'h00000000000000000000000000000000, /* 3468 */
128'h00000000000000000000000000000000, /* 3469 */
128'h00000000000000000000000000000000, /* 3470 */
128'h00000000000000000000000000000000, /* 3471 */
128'h00000000000000000000000000000000, /* 3472 */
128'h00000000000000000000000000000000, /* 3473 */
128'h00000000000000000000000000000000, /* 3474 */
128'h00000000000000000000000000000000, /* 3475 */
128'h00000000000000000000000000000000, /* 3476 */
128'h00000000000000000000000000000000, /* 3477 */
128'h00000000000000000000000000000000, /* 3478 */
128'h00000000000000000000000000000000, /* 3479 */
128'h00000000000000000000000000000000, /* 3480 */
128'h00000000000000000000000000000000, /* 3481 */
128'h00000000000000000000000000000000, /* 3482 */
128'h00000000000000000000000000000000, /* 3483 */
128'h00000000000000000000000000000000, /* 3484 */
128'h00000000000000000000000000000000, /* 3485 */
128'h00000000000000000000000000000000, /* 3486 */
128'h00000000000000000000000000000000, /* 3487 */
128'h00000000000000000000000000000000, /* 3488 */
128'h00000000000000000000000000000000, /* 3489 */
128'h00000000000000000000000000000000, /* 3490 */
128'h00000000000000000000000000000000, /* 3491 */
128'h00000000000000000000000000000000, /* 3492 */
128'h00000000000000000000000000000000, /* 3493 */
128'h00000000000000000000000000000000, /* 3494 */
128'h00000000000000000000000000000000, /* 3495 */
128'h00000000000000000000000000000000, /* 3496 */
128'h00000000000000000000000000000000, /* 3497 */
128'h00000000000000000000000000000000, /* 3498 */
128'h00000000000000000000000000000000, /* 3499 */
128'h00000000000000000000000000000000, /* 3500 */
128'h00000000000000000000000000000000, /* 3501 */
128'h00000000000000000000000000000000, /* 3502 */
128'h00000000000000000000000000000000, /* 3503 */
128'h00000000000000000000000000000000, /* 3504 */
128'h00000000000000000000000000000000, /* 3505 */
128'h00000000000000000000000000000000, /* 3506 */
128'h00000000000000000000000000000000, /* 3507 */
128'h00000000000000000000000000000000, /* 3508 */
128'h00000000000000000000000000000000, /* 3509 */
128'h00000000000000000000000000000000, /* 3510 */
128'h00000000000000000000000000000000, /* 3511 */
128'h00000000000000000000000000000000, /* 3512 */
128'h00000000000000000000000000000000, /* 3513 */
128'h00000000000000000000000000000000, /* 3514 */
128'h00000000000000000000000000000000, /* 3515 */
128'h00000000000000000000000000000000, /* 3516 */
128'h00000000000000000000000000000000, /* 3517 */
128'h00000000000000000000000000000000, /* 3518 */
128'h00000000000000000000000000000000, /* 3519 */
128'h00000000000000000000000000000000, /* 3520 */
128'h00000000000000000000000000000000, /* 3521 */
128'h00000000000000000000000000000000, /* 3522 */
128'h00000000000000000000000000000000, /* 3523 */
128'h00000000000000000000000000000000, /* 3524 */
128'h00000000000000000000000000000000, /* 3525 */
128'h00000000000000000000000000000000, /* 3526 */
128'h00000000000000000000000000000000, /* 3527 */
128'h00000000000000000000000000000000, /* 3528 */
128'h00000000000000000000000000000000, /* 3529 */
128'h00000000000000000000000000000000, /* 3530 */
128'h00000000000000000000000000000000, /* 3531 */
128'h00000000000000000000000000000000, /* 3532 */
128'h00000000000000000000000000000000, /* 3533 */
128'h00000000000000000000000000000000, /* 3534 */
128'h00000000000000000000000000000000, /* 3535 */
128'h00000000000000000000000000000000, /* 3536 */
128'h00000000000000000000000000000000, /* 3537 */
128'h00000000000000000000000000000000, /* 3538 */
128'h00000000000000000000000000000000, /* 3539 */
128'h00000000000000000000000000000000, /* 3540 */
128'h00000000000000000000000000000000, /* 3541 */
128'h00000000000000000000000000000000, /* 3542 */
128'h00000000000000000000000000000000, /* 3543 */
128'h00000000000000000000000000000000, /* 3544 */
128'h00000000000000000000000000000000, /* 3545 */
128'h00000000000000000000000000000000, /* 3546 */
128'h00000000000000000000000000000000, /* 3547 */
128'h00000000000000000000000000000000, /* 3548 */
128'h00000000000000000000000000000000, /* 3549 */
128'h00000000000000000000000000000000, /* 3550 */
128'h00000000000000000000000000000000, /* 3551 */
128'h00000000000000000000000000000000, /* 3552 */
128'h00000000000000000000000000000000, /* 3553 */
128'h00000000000000000000000000000000, /* 3554 */
128'h00000000000000000000000000000000, /* 3555 */
128'h00000000000000000000000000000000, /* 3556 */
128'h00000000000000000000000000000000, /* 3557 */
128'h00000000000000000000000000000000, /* 3558 */
128'h00000000000000000000000000000000, /* 3559 */
128'h00000000000000000000000000000000, /* 3560 */
128'h00000000000000000000000000000000, /* 3561 */
128'h00000000000000000000000000000000, /* 3562 */
128'h00000000000000000000000000000000, /* 3563 */
128'h00000000000000000000000000000000, /* 3564 */
128'h00000000000000000000000000000000, /* 3565 */
128'h00000000000000000000000000000000, /* 3566 */
128'h00000000000000000000000000000000, /* 3567 */
128'h00000000000000000000000000000000, /* 3568 */
128'h00000000000000000000000000000000, /* 3569 */
128'h00000000000000000000000000000000, /* 3570 */
128'h00000000000000000000000000000000, /* 3571 */
128'h00000000000000000000000000000000, /* 3572 */
128'h00000000000000000000000000000000, /* 3573 */
128'h00000000000000000000000000000000, /* 3574 */
128'h00000000000000000000000000000000, /* 3575 */
128'h00000000000000000000000000000000, /* 3576 */
128'h00000000000000000000000000000000, /* 3577 */
128'h00000000000000000000000000000000, /* 3578 */
128'h00000000000000000000000000000000, /* 3579 */
128'h00000000000000000000000000000000, /* 3580 */
128'h00000000000000000000000000000000, /* 3581 */
128'h00000000000000000000000000000000, /* 3582 */
128'h00000000000000000000000000000000, /* 3583 */
128'h00000000000000000000000000000000, /* 3584 */
128'h00000000000000000000000000000000, /* 3585 */
128'h00000000000000000000000000000000, /* 3586 */
128'h00000000000000000000000000000000, /* 3587 */
128'h00000000000000000000000000000000, /* 3588 */
128'h00000000000000000000000000000000, /* 3589 */
128'h00000000000000000000000000000000, /* 3590 */
128'h00000000000000000000000000000000, /* 3591 */
128'h00000000000000000000000000000000, /* 3592 */
128'h00000000000000000000000000000000, /* 3593 */
128'h00000000000000000000000000000000, /* 3594 */
128'h00000000000000000000000000000000, /* 3595 */
128'h00000000000000000000000000000000, /* 3596 */
128'h00000000000000000000000000000000, /* 3597 */
128'h00000000000000000000000000000000, /* 3598 */
128'h00000000000000000000000000000000, /* 3599 */
128'h00000000000000000000000000000000, /* 3600 */
128'h00000000000000000000000000000000, /* 3601 */
128'h00000000000000000000000000000000, /* 3602 */
128'h00000000000000000000000000000000, /* 3603 */
128'h00000000000000000000000000000000, /* 3604 */
128'h00000000000000000000000000000000, /* 3605 */
128'h00000000000000000000000000000000, /* 3606 */
128'h00000000000000000000000000000000, /* 3607 */
128'h00000000000000000000000000000000, /* 3608 */
128'h00000000000000000000000000000000, /* 3609 */
128'h00000000000000000000000000000000, /* 3610 */
128'h00000000000000000000000000000000, /* 3611 */
128'h00000000000000000000000000000000, /* 3612 */
128'h00000000000000000000000000000000, /* 3613 */
128'h00000000000000000000000000000000, /* 3614 */
128'h00000000000000000000000000000000, /* 3615 */
128'h00000000000000000000000000000000, /* 3616 */
128'h00000000000000000000000000000000, /* 3617 */
128'h00000000000000000000000000000000, /* 3618 */
128'h00000000000000000000000000000000, /* 3619 */
128'h00000000000000000000000000000000, /* 3620 */
128'h00000000000000000000000000000000, /* 3621 */
128'h00000000000000000000000000000000, /* 3622 */
128'h00000000000000000000000000000000, /* 3623 */
128'h00000000000000000000000000000000, /* 3624 */
128'h00000000000000000000000000000000, /* 3625 */
128'h00000000000000000000000000000000, /* 3626 */
128'h00000000000000000000000000000000, /* 3627 */
128'h00000000000000000000000000000000, /* 3628 */
128'h00000000000000000000000000000000, /* 3629 */
128'h00000000000000000000000000000000, /* 3630 */
128'h00000000000000000000000000000000, /* 3631 */
128'h00000000000000000000000000000000, /* 3632 */
128'h00000000000000000000000000000000, /* 3633 */
128'h00000000000000000000000000000000, /* 3634 */
128'h00000000000000000000000000000000, /* 3635 */
128'h00000000000000000000000000000000, /* 3636 */
128'h00000000000000000000000000000000, /* 3637 */
128'h00000000000000000000000000000000, /* 3638 */
128'h00000000000000000000000000000000, /* 3639 */
128'h00000000000000000000000000000000, /* 3640 */
128'h00000000000000000000000000000000, /* 3641 */
128'h00000000000000000000000000000000, /* 3642 */
128'h00000000000000000000000000000000, /* 3643 */
128'h00000000000000000000000000000000, /* 3644 */
128'h00000000000000000000000000000000, /* 3645 */
128'h00000000000000000000000000000000, /* 3646 */
128'h00000000000000000000000000000000, /* 3647 */
128'h00000000000000000000000000000000, /* 3648 */
128'h00000000000000000000000000000000, /* 3649 */
128'h00000000000000000000000000000000, /* 3650 */
128'h00000000000000000000000000000000, /* 3651 */
128'h00000000000000000000000000000000, /* 3652 */
128'h00000000000000000000000000000000, /* 3653 */
128'h00000000000000000000000000000000, /* 3654 */
128'h00000000000000000000000000000000, /* 3655 */
128'h00000000000000000000000000000000, /* 3656 */
128'h00000000000000000000000000000000, /* 3657 */
128'h00000000000000000000000000000000, /* 3658 */
128'h00000000000000000000000000000000, /* 3659 */
128'h00000000000000000000000000000000, /* 3660 */
128'h00000000000000000000000000000000, /* 3661 */
128'h00000000000000000000000000000000, /* 3662 */
128'h00000000000000000000000000000000, /* 3663 */
128'h00000000000000000000000000000000, /* 3664 */
128'h00000000000000000000000000000000, /* 3665 */
128'h00000000000000000000000000000000, /* 3666 */
128'h00000000000000000000000000000000, /* 3667 */
128'h00000000000000000000000000000000, /* 3668 */
128'h00000000000000000000000000000000, /* 3669 */
128'h00000000000000000000000000000000, /* 3670 */
128'h00000000000000000000000000000000, /* 3671 */
128'h00000000000000000000000000000000, /* 3672 */
128'h00000000000000000000000000000000, /* 3673 */
128'h00000000000000000000000000000000, /* 3674 */
128'h00000000000000000000000000000000, /* 3675 */
128'h00000000000000000000000000000000, /* 3676 */
128'h00000000000000000000000000000000, /* 3677 */
128'h00000000000000000000000000000000, /* 3678 */
128'h00000000000000000000000000000000, /* 3679 */
128'h00000000000000000000000000000000, /* 3680 */
128'h00000000000000000000000000000000, /* 3681 */
128'h00000000000000000000000000000000, /* 3682 */
128'h00000000000000000000000000000000, /* 3683 */
128'h00000000000000000000000000000000, /* 3684 */
128'h00000000000000000000000000000000, /* 3685 */
128'h00000000000000000000000000000000, /* 3686 */
128'h00000000000000000000000000000000, /* 3687 */
128'h00000000000000000000000000000000, /* 3688 */
128'h00000000000000000000000000000000, /* 3689 */
128'h00000000000000000000000000000000, /* 3690 */
128'h00000000000000000000000000000000, /* 3691 */
128'h00000000000000000000000000000000, /* 3692 */
128'h00000000000000000000000000000000, /* 3693 */
128'h00000000000000000000000000000000, /* 3694 */
128'h00000000000000000000000000000000, /* 3695 */
128'h00000000000000000000000000000000, /* 3696 */
128'h00000000000000000000000000000000, /* 3697 */
128'h00000000000000000000000000000000, /* 3698 */
128'h00000000000000000000000000000000, /* 3699 */
128'h00000000000000000000000000000000, /* 3700 */
128'h00000000000000000000000000000000, /* 3701 */
128'h00000000000000000000000000000000, /* 3702 */
128'h00000000000000000000000000000000, /* 3703 */
128'h00000000000000000000000000000000, /* 3704 */
128'h00000000000000000000000000000000, /* 3705 */
128'h00000000000000000000000000000000, /* 3706 */
128'h00000000000000000000000000000000, /* 3707 */
128'h00000000000000000000000000000000, /* 3708 */
128'h00000000000000000000000000000000, /* 3709 */
128'h00000000000000000000000000000000, /* 3710 */
128'h00000000000000000000000000000000, /* 3711 */
128'h00000000000000000000000000000000, /* 3712 */
128'h00000000000000000000000000000000, /* 3713 */
128'h00000000000000000000000000000000, /* 3714 */
128'h00000000000000000000000000000000, /* 3715 */
128'h00000000000000000000000000000000, /* 3716 */
128'h00000000000000000000000000000000, /* 3717 */
128'h00000000000000000000000000000000, /* 3718 */
128'h00000000000000000000000000000000, /* 3719 */
128'h00000000000000000000000000000000, /* 3720 */
128'h00000000000000000000000000000000, /* 3721 */
128'h00000000000000000000000000000000, /* 3722 */
128'h00000000000000000000000000000000, /* 3723 */
128'h00000000000000000000000000000000, /* 3724 */
128'h00000000000000000000000000000000, /* 3725 */
128'h00000000000000000000000000000000, /* 3726 */
128'h00000000000000000000000000000000, /* 3727 */
128'h00000000000000000000000000000000, /* 3728 */
128'h00000000000000000000000000000000, /* 3729 */
128'h00000000000000000000000000000000, /* 3730 */
128'h00000000000000000000000000000000, /* 3731 */
128'h00000000000000000000000000000000, /* 3732 */
128'h00000000000000000000000000000000, /* 3733 */
128'h00000000000000000000000000000000, /* 3734 */
128'h00000000000000000000000000000000, /* 3735 */
128'h00000000000000000000000000000000, /* 3736 */
128'h00000000000000000000000000000000, /* 3737 */
128'h00000000000000000000000000000000, /* 3738 */
128'h00000000000000000000000000000000, /* 3739 */
128'h00000000000000000000000000000000, /* 3740 */
128'h00000000000000000000000000000000, /* 3741 */
128'h00000000000000000000000000000000, /* 3742 */
128'h00000000000000000000000000000000, /* 3743 */
128'h00000000000000000000000000000000, /* 3744 */
128'h00000000000000000000000000000000, /* 3745 */
128'h00000000000000000000000000000000, /* 3746 */
128'h00000000000000000000000000000000, /* 3747 */
128'h00000000000000000000000000000000, /* 3748 */
128'h00000000000000000000000000000000, /* 3749 */
128'h00000000000000000000000000000000, /* 3750 */
128'h00000000000000000000000000000000, /* 3751 */
128'h00000000000000000000000000000000, /* 3752 */
128'h00000000000000000000000000000000, /* 3753 */
128'h00000000000000000000000000000000, /* 3754 */
128'h00000000000000000000000000000000, /* 3755 */
128'h00000000000000000000000000000000, /* 3756 */
128'h00000000000000000000000000000000, /* 3757 */
128'h00000000000000000000000000000000, /* 3758 */
128'h00000000000000000000000000000000, /* 3759 */
128'h00000000000000000000000000000000, /* 3760 */
128'h00000000000000000000000000000000, /* 3761 */
128'h00000000000000000000000000000000, /* 3762 */
128'h00000000000000000000000000000000, /* 3763 */
128'h00000000000000000000000000000000, /* 3764 */
128'h00000000000000000000000000000000, /* 3765 */
128'h00000000000000000000000000000000, /* 3766 */
128'h00000000000000000000000000000000, /* 3767 */
128'h00000000000000000000000000000000, /* 3768 */
128'h00000000000000000000000000000000, /* 3769 */
128'h00000000000000000000000000000000, /* 3770 */
128'h00000000000000000000000000000000, /* 3771 */
128'h00000000000000000000000000000000, /* 3772 */
128'h00000000000000000000000000000000, /* 3773 */
128'h00000000000000000000000000000000, /* 3774 */
128'h00000000000000000000000000000000, /* 3775 */
128'h00000000000000000000000000000000, /* 3776 */
128'h00000000000000000000000000000000, /* 3777 */
128'h00000000000000000000000000000000, /* 3778 */
128'h00000000000000000000000000000000, /* 3779 */
128'h00000000000000000000000000000000, /* 3780 */
128'h00000000000000000000000000000000, /* 3781 */
128'h00000000000000000000000000000000, /* 3782 */
128'h00000000000000000000000000000000, /* 3783 */
128'h00000000000000000000000000000000, /* 3784 */
128'h00000000000000000000000000000000, /* 3785 */
128'h00000000000000000000000000000000, /* 3786 */
128'h00000000000000000000000000000000, /* 3787 */
128'h00000000000000000000000000000000, /* 3788 */
128'h00000000000000000000000000000000, /* 3789 */
128'h00000000000000000000000000000000, /* 3790 */
128'h00000000000000000000000000000000, /* 3791 */
128'h00000000000000000000000000000000, /* 3792 */
128'h00000000000000000000000000000000, /* 3793 */
128'h00000000000000000000000000000000, /* 3794 */
128'h00000000000000000000000000000000, /* 3795 */
128'h00000000000000000000000000000000, /* 3796 */
128'h00000000000000000000000000000000, /* 3797 */
128'h00000000000000000000000000000000, /* 3798 */
128'h00000000000000000000000000000000, /* 3799 */
128'h00000000000000000000000000000000, /* 3800 */
128'h00000000000000000000000000000000, /* 3801 */
128'h00000000000000000000000000000000, /* 3802 */
128'h00000000000000000000000000000000, /* 3803 */
128'h00000000000000000000000000000000, /* 3804 */
128'h00000000000000000000000000000000, /* 3805 */
128'h00000000000000000000000000000000, /* 3806 */
128'h00000000000000000000000000000000, /* 3807 */
128'h00000000000000000000000000000000, /* 3808 */
128'h00000000000000000000000000000000, /* 3809 */
128'h00000000000000000000000000000000, /* 3810 */
128'h00000000000000000000000000000000, /* 3811 */
128'h00000000000000000000000000000000, /* 3812 */
128'h00000000000000000000000000000000, /* 3813 */
128'h00000000000000000000000000000000, /* 3814 */
128'h00000000000000000000000000000000, /* 3815 */
128'h00000000000000000000000000000000, /* 3816 */
128'h00000000000000000000000000000000, /* 3817 */
128'h00000000000000000000000000000000, /* 3818 */
128'h00000000000000000000000000000000, /* 3819 */
128'h00000000000000000000000000000000, /* 3820 */
128'h00000000000000000000000000000000, /* 3821 */
128'h00000000000000000000000000000000, /* 3822 */
128'h00000000000000000000000000000000, /* 3823 */
128'h00000000000000000000000000000000, /* 3824 */
128'h00000000000000000000000000000000, /* 3825 */
128'h00000000000000000000000000000000, /* 3826 */
128'h00000000000000000000000000000000, /* 3827 */
128'h00000000000000000000000000000000, /* 3828 */
128'h00000000000000000000000000000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00000000000000000000000000000000, /* 3840 */
128'h00000000000000000000000000000000, /* 3841 */
128'h00000000000000000000000000000000, /* 3842 */
128'h00000000000000000000000000000000, /* 3843 */
128'h00000000000000000000000000000000, /* 3844 */
128'h00000000000000000000000000000000, /* 3845 */
128'h00000000000000000000000000000000, /* 3846 */
128'h00000000000000000000000000000000, /* 3847 */
128'h00000000000000000000000000000000, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule

