/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module etherboot (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 5991;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_bffe70de,
        64'h00000000_bffe711c,
        64'h00000000_00000000,
        64'hffffffff_00000006,
        64'h00000000_bffeb428,
        64'h00000000_2f7c5c2d,
        64'h00000000_ffffffff,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_cc33aa55,
        64'h00000000_bffeb270,
        64'h00006772_615f6473,
        64'h0000646d_635f6473,
        64'h00000000_0c000000,
        64'h00000000_ffffffff,
        64'h00000000_00000000,
        64'h00000000_30000000,
        64'h00000000_004b4d47,
        64'h00004b4d_47545045,
        64'h00000003_0f060301,
        64'haaaaaaaa_aaaaaaaa,
        64'h55555555_55555555,
        64'h5851f42d_4c957f2d,
        64'h10000000_20000000,
        64'h10325476_98badcfe,
        64'hefcdab89_67452301,
        64'hcccccccc_cccccccd,
        64'h00000a0d_70617274,
        64'h00000000_000a7473,
        64'h65742065_68636143,
        64'h00000000_00000a74,
        64'h6f6f6220_50544654,
        64'h00000000_00000a74,
        64'h73657420_4d415244,
        64'h00000000_00000a74,
        64'h6f6f6220_49505351,
        64'h00000000_00000000,
        64'h0a746f6f_62204453,
        64'h00000000_0000000a,
        64'h5825203d_20646565,
        64'h73206d6f_646e6152,
        64'h000a5825_2c582520,
        64'h3d20676e_69747465,
        64'h73206863_74697753,
        64'h0000000a_5825203d,
        64'h205d6425_5b707773,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h0a646c25_2e646c25,
        64'h203d2049_5043202c,
        64'h73656c63_79632064,
        64'h6c25202c_736e6f69,
        64'h74637572_74736e69,
        64'h20646c25_202c424b,
        64'h6425203d_20746573,
        64'h5f676e69_6b726f77,
        64'h00000000_00000000,
        64'h0a2e2979_6c6e6f28,
        64'h2032206e_6f697372,
        64'h65762065_736e6563,
        64'h694c2063_696c6275,
        64'h50206c61_72656e65,
        64'h4720554e_47206568,
        64'h74207265_646e7520,
        64'h6465736e_6563694c,
        64'h00000000_0000000a,
        64'h2e6e6f62_617a6143,
        64'h2073656c_72616843,
        64'h20323130_322d3130,
        64'h30322029_43282074,
        64'h68676972_79706f43,
        64'h00000000_0000000a,
        64'h29746962_2d642528,
        64'h20302e33_2e34206e,
        64'h6f697372_65762072,
        64'h65747365_746d656d,
        64'h00000a74_73657420,
        64'h4d415244_206c6174,
        64'h656d2065_7261420a,
        64'h00000a2e_656e6f44,
        64'h00000000_000a6b6f,
        64'h0000203a_73252020,
        64'h00000073_73657264,
        64'h6441206b_63757453,
        64'h00000000_00000a3a,
        64'h00000000_0075252f,
        64'h00752520_706f6f4c,
        64'h00000000_000a7025,
        64'h7830206f_74207025,
        64'h78302073_69206567,
        64'h6e617220_74736574,
        64'h00000000_00082008,
        64'h00000000_00000008,
        64'h08080808_08080808,
        64'h08082020_20202020,
        64'h20202020_20080808,
        64'h08080808_08080808,
        64'h00000000_0000000a,
        64'h2e2e2e74_73657420,
        64'h7478656e_206f7420,
        64'h676e6970_70696b53,
        64'h00000000_000a2e78,
        64'h25783020_74657366,
        64'h666f2074_6120656e,
        64'h696c2073_73657264,
        64'h64612064_61622065,
        64'h6c626973_736f7020,
        64'h3a455255_4c494146,
        64'h00000000_00007525,
        64'h20676e69_74736574,
        64'h00000000_00007525,
        64'h20676e69_74746573,
        64'h00000000_00080808,
        64'h08080808_08080808,
        64'h00000000_00202020,
        64'h20202020_20202020,
        64'h00000000_0000000a,
        64'h7025203d_20327020,
        64'h2c702520_3d203170,
        64'h00000a2e_78257830,
        64'h20746573_66666f20,
        64'h74612078_25783020,
        64'h3d212078_25783020,
        64'h3a455255_4c494146,
        64'h00000000_000a7325,
        64'h206e6f69_74636e75,
        64'h66202c64_2520656e,
        64'h696c202c_73252065,
        64'h6c696620_2c64656c,
        64'h69616620_7325206e,
        64'h6f697472_65737361,
        64'h00000a72_6564616f,
        64'h6c20746f_6f622065,
        64'h67617473_20747372,
        64'h69662064_65736162,
        64'h20746f6f_622d750a,
        64'h00000000_5c2d2f7c,
        64'h00000000_64252065,
        64'h646f6320_68746977,
        64'h2064656c_69616620,
        64'h64616572_20666c65,
        64'h000a7972_6f6d656d,
        64'h20524444_206f7420,
        64'h666c6520_64616f6c,
        64'h00000000_00000000,
        64'h0a2e7365_74796220,
        64'h64252066_6f206e69,
        64'h622e746f_6f62206d,
        64'h6f726620_78252073,
        64'h73657264_64612079,
        64'h726f6d65_6d206f74,
        64'h20736574_79622064,
        64'h25206465_64616f4c,
        64'h00000000_216b7369,
        64'h6420746e_756f6d75,
        64'h206f7420_6c696166,
        64'h00000000_0021656c,
        64'h69662065_736f6c63,
        64'h206f7420_6c696166,
        64'h0000000a_21746f6f,
        64'h62206e65_706f206f,
        64'h74206465_6c696146,
        64'h00000000_00000000,
        64'h6e69622e_746f6f62,
        64'h00000000_00000a79,
        64'h726f6d65_6d206f74,
        64'h6e69206e_69622e74,
        64'h6f6f6220_64616f4c,
        64'h00000000_0000000a,
        64'h21726576_69726420,
        64'h44532074_6e756f6d,
        64'h206f7420_6c696146,
        64'h00000000_00000000,
        64'h0a2e6e6f_69746172,
        64'h65706f20_50544654,
        64'h206c6167_656c6c49,
        64'h00000000_000a2e64,
        64'h656c6c61_63207172,
        64'h775f656c_646e6168,
        64'h00000000_00000a2e,
        64'h646e6520_656c6966,
        64'h20657669_65636552,
        64'h00000000_00000000,
        64'h0a64253d_657a6973,
        64'h6b636f6c_62202c22,
        64'h73252220_3a717277,
        64'h00000000_0000002f,
        64'h00000000_000a646c,
        64'h25202e67_6e6f6c20,
        64'h6f6f7420_68746170,
        64'h20747365_75716552,
        64'h00000000_00000000,
        64'h0a732520_3d202964,
        64'h252c7025_2835646d,
        64'h00000000_0000000a,
        64'h6425203d_20687467,
        64'h6e656c20_656c6946,
        64'h00000000_00636d6d,
        64'h00000029_73252820,
        64'h00006425_203a7325,
        64'h00000000_434d4d65,
        64'h00000000_00004453,
        64'h00000000_00000000,
        64'h0a646e75_6f662074,
        64'h6f6e2064_25206563,
        64'h69766544_20434d4d,
        64'h0000297a_484d3030,
        64'h32282030_30325348,
        64'h00000000_00297a48,
        64'h4d383032_28203430,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282030,
        64'h35524444_20534855,
        64'h00000000_0000297a,
        64'h484d3030_31282030,
        64'h35524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282035,
        64'h32524453_20534855,
        64'h00000000_00000029,
        64'h7a484d35_32282032,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d32_35282032,
        64'h35524444_20434d4d,
        64'h0000297a_484d3235,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000029_7a484d30,
        64'h35282064_65657053,
        64'h20686769_48204453,
        64'h0000297a_484d3632,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000000_00000079,
        64'h63616765_4c204453,
        64'h00000000_00007963,
        64'h6167656c_20434d4d,
        64'h00000064_252e6425,
        64'h00000000_63256325,
        64'h63256325_63256325,
        64'h00000078_34302578,
        64'h34302520_726e5320,
        64'h78363025_206e614d,
        64'h00000000_00000a21,
        64'h646e756f_66206473,
        64'h635f7478_65206f4e,
        64'h00000000_00000000,
        64'h0a65646f_6d206120,
        64'h7463656c_6573206f,
        64'h7420656c_62616e75,
        64'h00000000_00000000,
        64'h0a217463_656c6573,
        64'h20656761_746c6f76,
        64'h206f7420_646e6f70,
        64'h73657220_746f6e20,
        64'h64696420_64726143,
        64'h0000000a_746e6573,
        64'h65727020_64726163,
        64'h206f6e20_3a434d4d,
        64'h00000000_0000000a,
        64'h64656e6f_69746974,
        64'h72617020_79646165,
        64'h726c6120_64726143,
        64'h00000000_000a7367,
        64'h6e697474_65732079,
        64'h74696c69_6261696c,
        64'h65722065_74697277,
        64'h206e6f69_74697472,
        64'h61702064_656c6c6f,
        64'h72746e6f_63207473,
        64'h6f682074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000a29_7525203e,
        64'h20752528_206d756d,
        64'h6978616d_20736465,
        64'h65637865_20657a69,
        64'h73206465_636e6168,
        64'h6e65206c_61746f54,
        64'h00000000_0000000a,
        64'h65747562_69727474,
        64'h61206465_636e6168,
        64'h6e652074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0a64656e,
        64'h67696c61_20657a69,
        64'h73207075_6f726720,
        64'h50572043_4820746f,
        64'h6e206e6f_69746974,
        64'h72617020_69255047,
        64'h0000000a_64656e67,
        64'h696c6120_657a6973,
        64'h2070756f_72672050,
        64'h57204348_20746f6e,
        64'h20616572_61206465,
        64'h636e6168_6e652061,
        64'h74616420_72657355,
        64'h00000a65_7a697320,
        64'h70756f72_67205057,
        64'h20434820_656e6966,
        64'h65642074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_000a676e,
        64'h696e6f69_74697472,
        64'h61702074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0000000a,
        64'h61657261_20617461,
        64'h64207265_73752064,
        64'h65636e61_686e6520,
        64'h726f6620_64657269,
        64'h75716572_20342e34,
        64'h203d3e20_434d4d65,
        64'h00000000_000a2978,
        64'h6c257830_2878616d,
        64'h20736465_65637865,
        64'h20786c25_78302072,
        64'h65626d75_6e206b63,
        64'h6f6c6220_3a434d4d,
        64'h00000000_00000a64,
        64'h6d632070_6f747320,
        64'h646e6573_206f7420,
        64'h6c696166_20636d6d,
        64'h00000000_000a7964,
        64'h61657220_64726163,
        64'h20676e69_74696177,
        64'h2074756f_656d6954,
        64'h0000000a_58383025,
        64'h7830203a_726f7272,
        64'h45207375_74617453,
        64'h00000000_65646f6d,
        64'h206e776f_6e6b6e55,
        64'h00000000_00006473,
        64'h5f637369_72776f6c,
        64'h00000078_25782520,
        64'h00000020_3a78250a,
        64'h00000000_0a732574,
        64'h69622d64_25203a68,
        64'h74646957_20737542,
        64'h00000000_0000203a,
        64'h79746963_61706143,
        64'h00000000_00000a73,
        64'h25203a79_74696361,
        64'h70614320_68676948,
        64'h00000a64_25203a64,
        64'h65657053_20737542,
        64'h00000000_00000a20,
        64'h63256325_63256325,
        64'h6325203a_656d614e,
        64'h00000000_00000000,
        64'h0a782520_3a4d454f,
        64'h00000000_0a782520,
        64'h3a444920_72657275,
        64'h74636166_756e614d,
        64'h00000000_000a7325,
        64'h203a6563_69766544,
        64'h00202020_3a434d4d,
        64'h00000000_52444420,
        64'h00000000_00006f4e,
        64'h00000000_00736559,
        64'h0000000a_7825203d,
        64'h2074736f_68202c78,
        64'h25207461_20646574,
        64'h61657263_20636d6d,
        64'h00000000_00000a64,
        64'h25206f74_20646567,
        64'h6e616863_206b7361,
        64'h6d202c64_65747265,
        64'h736e6920_64726143,
        64'h00000000_0000000a,
        64'h6425206f_74206465,
        64'h676e6168_63206b73,
        64'h616d202c_6465766f,
        64'h6d657220_64726143,
        64'h000a7475_6f656d69,
        64'h74207325_203a6473,
        64'h5f637369_72776f6c,
        64'h00726464_615f6573,
        64'h61625f64_73203d3d,
        64'h20657361_625f6473,
        64'h00000000_00000063,
        64'h2e636d6d_5f637369,
        64'h72776f6c_2f637273,
        64'h00000000_00000000,
        64'h66656463_62613938,
        64'h37363534_33323130,
        64'h007f7c5d_5b3f3e3d,
        64'h3c3b3a2e_2c2b2a22,
        64'h00007f7c_5d5b3f3e,
        64'h3d3c3b3a_2c2b2a22,
        64'h00000000_0a2e2e2e,
        64'h20726574_6f6f6220,
        64'h2c657962_646f6f47,
        64'h00000000_000a2e2e,
        64'h2e6d6172_676f7270,
        64'h20646564_616f6c20,
        64'h65687420_746f6f42,
        64'h00000000_00000000,
        64'h0a646c25_203d2073,
        64'h75746174_73207470,
        64'h75727265_746e6920,
        64'h74656e72_65687445,
        64'h0000000a_2e783230,
        64'h253a7832_30253a78,
        64'h3230253a_78323025,
        64'h3a783230_253a7832,
        64'h3025203d_20737365,
        64'h72646461_2043414d,
        64'h00000a78_6c253a78,
        64'h6c25203d_2043414d,
        64'h00000000_00000a78,
        64'h25203d20_5d64255b,
        64'h4d454f20_49505351,
        64'h000a7264_64612043,
        64'h414d2070_75746553,
        64'h0000000a_21747075,
        64'h72726574_6e692064,
        64'h656c646e_61686e75,
        64'h00000000_00000a78,
        64'h25783020_3d206570,
        64'h79745f6f_746f7270,
        64'h00000000_0a297825,
        64'h28206465_74726f70,
        64'h7075736e_75203d20,
        64'h6f746f72_70205049,
        64'h000a5741_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a534c50_4d203d20,
        64'h6f746f72_50205049,
        64'h00000000_000a4554,
        64'h494c5044_55203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505443_53203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a504d4f_43203d20,
        64'h6f746f72_50205049,
        64'h00000000_0000004d,
        64'h00000000_0000000a,
        64'h5041434e_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000a48,
        64'h50544545_42203d20,
        64'h6f746f72_50205049,
        64'h000a5054_4d203d20,
        64'h6f746f72_50205049,
        64'h00000a48_41203d20,
        64'h6f746f72_50205049,
        64'h000a5053_45203d20,
        64'h6f746f72_50205049,
        64'h000a4552_47203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505653_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000036,
        64'h00000000_00000000,
        64'h0a504343_44203d20,
        64'h6f746f72_50205049,
        64'h00000a50_54203d20,
        64'h6f746f72_50205049,
        64'h000a5044_49203d20,
        64'h6f746f72_50205049,
        64'h000a3a73_746e6574,
        64'h6e6f6320_74736574,
        64'h0000000a_3a726564,
        64'h61656820_74736574,
        64'h000a5055_50203d20,
        64'h6f746f72_50205049,
        64'h000a5047_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000054,
        64'h00000000_00000000,
        64'h0a504950_49203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000047,
        64'h00006425_2b544553,
        64'h46464f5f_524c5052,
        64'h00000000_3f3f3f3f,
        64'h00000000_00544553,
        64'h46464f5f_524c5052,
        64'h00000000_00544553,
        64'h46464f5f_44414252,
        64'h00000000_00005445,
        64'h5346464f_5f525352,
        64'h00000000_00544553,
        64'h46464f5f_53434652,
        64'h00544553_46464f5f,
        64'h4c525443_4f49444d,
        64'h00000000_00544553,
        64'h46464f5f_53434654,
        64'h00000000_00544553,
        64'h46464f5f_524c5054,
        64'h00000000_54455346,
        64'h464f5f49_4843414d,
        64'h00000000_54455346,
        64'h464f5f4f_4c43414d,
        64'h00000000_000a3b29,
        64'h78257830_2c302c78,
        64'h25287465_736d656d,
        64'h00000a3b_29782578,
        64'h302c7825_78302c78,
        64'h25287970_636d656d,
        64'h000a7825_203d206c,
        64'h61757463_61202c58,
        64'h25203d20_64657269,
        64'h75716572_206e656c,
        64'h00000020_3a5d6425,
        64'h5b6e6f69_74636553,
        64'h000a7325_20202020,
        64'h00786c6c_2a302520,
        64'h00003a78_6c383025,
        64'h00732542_69632520,
        64'h00000000_00732573,
        64'h65747942_20756c25,
        64'h0073257a_48632520,
        64'h00000000_646c252e,
        64'h00000000_00756c25,
        64'h00000000_00000000,
        64'h73257a48_20756c25,
        64'h00000000_00007325,
        64'h00000000_00732520,
        64'h3a646c69_7542202c,
        64'h00000000_73257325,
        64'h00000000_00000a0a,
        64'h00000058_32302520,
        64'h00000000_0000002e,
        64'h00000000_00006325,
        64'h00000000_00000020,
        64'h20202020_20202020,
        64'h000a5245_46464f5f,
        64'h50434844_20726f66,
        64'h20676e69_74696157,
        64'h00000a73_25203a73,
        64'h25206563_69766564,
        64'h206e6f20_59524556,
        64'h4f435349_44205043,
        64'h48442064_6e657320,
        64'h74276e64_6c756f43,
        64'h000a5832_30253a58,
        64'h3230253a_58323025,
        64'h3a583230_253a5832,
        64'h30253a58_32302520,
        64'h3a204341_4d207325,
        64'h00000000_30687465,
        64'h00000000_000a2973,
        64'h2528726f_72726570,
        64'h000a5952_45564f43,
        64'h5349445f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_0000000a,
        64'h64252065_646f6370,
        64'h6f205043_48442064,
        64'h656c646e_61686e55,
        64'h00000000_0a642520,
        64'h6e6f6974_706f2064,
        64'h656c646e_61686e75,
        64'h00000000_0000000a,
        64'h73252072_6f727245,
        64'h00000000_00000a64,
        64'h65737566_65722073,
        64'h73657264_64612064,
        64'h65747365_75716552,
        64'h00000000_0000000a,
        64'h4b414e20_50434844,
        64'h00000000_0a444550,
        64'h50494b53_204b4341,
        64'h000a2273_2522203d,
        64'h20656d61_6e74736f,
        64'h4820746e_65696c43,
        64'h00000a22_73252220,
        64'h3d206e69_616d6f44,
        64'h00000000_0000000a,
        64'h7364253a_6d64253a,
        64'h68642520_3d20656d,
        64'h69742065_7361654c,
        64'h000a6425_2e64252e,
        64'h64252e64_2520203a,
        64'h73736572_64646120,
        64'h6b73616d_2074654e,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h61207265_74756f52,
        64'h00000000_00000000,
        64'h0a64252e_64252e64,
        64'h252e6425_20203a73,
        64'h73657264_64412050,
        64'h49207265_76726553,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h41205049_20746e65,
        64'h696c4320_50434844,
        64'h00000000_0000000a,
        64'h4b434120_50434844,
        64'h0000000a_54534555,
        64'h5145525f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_00000000,
        64'h0a702520_2c726f72,
        64'h7265206c_616e7265,
        64'h746e6920_70636864,
        64'h00000a29_73252c73,
        64'h25287075_6b6f6f6c,
        64'h000a6563_69766564,
        64'h206e776f_6e6b6e75,
        64'h00000000_203a6425,
        64'h20656369_7665440a,
        64'h00203a64_25206563,
        64'h69766564_2073250a,
        64'h00000000_00203a64,
        64'h25206563_69766544,
        64'h00000000_00000000,
        64'h73736572_6464612d,
        64'h63616d2d_6c61636f,
        64'h6c006874_6469772d,
        64'h6f692d67_65720074,
        64'h66696873_2d676572,
        64'h00737470_75727265,
        64'h746e6900_746e6572,
        64'h61702d74_70757272,
        64'h65746e69_00646565,
        64'h70732d74_6e657272,
        64'h75630076_65646e2c,
        64'h76637369_72007974,
        64'h69726f69_72702d78,
        64'h616d2c76_63736972,
        64'h0073656d_616e2d67,
        64'h65720064_65646e65,
        64'h7478652d_73747075,
        64'h72726574_6e690073,
        64'h65676e61_7200656c,
        64'h646e6168_702c7875,
        64'h6e696c00_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h00100000_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_00000064,
        64'h6e727768_2d637369,
        64'h72776f6c_1b000000,
        64'h0e000000_03000000,
        64'h00003030_30303030,
        64'h30344064_6e727768,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h00800000_00000000,
        64'h00000030_00000000,
        64'h67000000_10000000,
        64'h03000000_00007fe3,
        64'h023e1800_47010000,
        64'h06000000_03000000,
        64'h03000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_00636d6d,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_02000000,
        64'h25010000_04000000,
        64'h03000000_02000000,
        64'h14010000_04000000,
        64'h03000000_00000100,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40636d6d,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h04000000_3a010000,
        64'h04000000_03000000,
        64'h02000000_30010000,
        64'h04000000_03000000,
        64'h01000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h00c20100_06010000,
        64'h04000000_03000000,
        64'h80f0fa02_4b000000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000010_00000000,
        64'h67000000_10000000,
        64'h03000000_00303537,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000000,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'hffff0000_01000000,
        64'hca000000_08000000,
        64'h03000000_00333130,
        64'h2d677562_65642c76,
        64'h63736972_1b000000,
        64'h10000000_03000000,
        64'h00003040_72656c6c,
        64'h6f72746e_6f632d67,
        64'h75626564_01000000,
        64'h02000000_02000000,
        64'hbb000000_04000000,
        64'h03000000_02000000,
        64'hb5000000_04000000,
        64'h03000000_03000000,
        64'hfb000000_04000000,
        64'h03000000_07000000,
        64'he8000000_04000000,
        64'h03000000_00000004,
        64'h00000000_0000000c,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h09000000_01000000,
        64'h0b000000_01000000,
        64'hca000000_10000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00000c00,
        64'h00000000_00000002,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_01000000,
        64'h03000000_01000000,
        64'hca000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6e696c63,
        64'h01000000_c3000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h01000000_bb000000,
        64'h04000000_03000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00007663_73697200,
        64'h656e6169_7261202c,
        64'h7a687465_1b000000,
        64'h13000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha8060000_59010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'he0060000_38000000,
        64'h39080000_edfe0dd0,
        64'h00000000_fffff9ba,
        64'hfffff980_fffff9a8,
        64'hfffff980_fffff996,
        64'hfffff982_fffff96e,
        64'h00000000_64726143,
        64'h2d445320_726f6620,
        64'h746f6f62_2d752064,
        64'h6573696d_696e696d,
        64'h20435349_52776f4c,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00020000_00010000,
        64'h0000c000_00008000,
        64'h00006000_00004000,
        64'h00002000_00001000,
        64'h00000800_00000400,
        64'h00000200_00000100,
        64'h00000080_00000040,
        64'h00000020_00000000,
        64'h0bebc200_0c65d400,
        64'h02faf080_05f5e100,
        64'h02faf080_017d7840,
        64'h03197500_03197500,
        64'h02faf080_018cba80,
        64'h017d7840_017d7840,
        64'h00989680_000f4240,
        64'h000186a0_00002710,
        64'h50463c37_322d2823,
        64'h1e19140f_0d0c0a00,
        64'h00000000_00000000,
        64'h00000000_10000000,
        64'h00000001_00000000,
        64'h20000000_00000002,
        64'h00000000_40000000,
        64'h00000005_00000001,
        64'h20000000_00000006,
        64'h00000001_40000000,
        64'h70000000_00000000,
        64'h70000000_00000002,
        64'h70000000_00000004,
        64'h60000000_00000005,
        64'h30000000_00000001,
        64'h30000000_00000003,
        64'h00000000_40050100,
        64'h40050000_40040500,
        64'h40040401_40040400,
        64'h40040300_40040200,
        64'h40040100_40040000,
        64'h00000000_bffeb3d8,
        64'h00000000_bffeb3c0,
        64'h00000000_bffeb3a8,
        64'h00000000_bffeb390,
        64'h00000000_bffeb378,
        64'h00000000_bffeb360,
        64'h00000000_bffeb348,
        64'h00000000_bffeb330,
        64'h00000000_bffeb318,
        64'h00000000_bffeb300,
        64'h00000000_bffeb2f0,
        64'h00000000_bffeb2e0,
        64'hffffcc04_ffffcbfe,
        64'hffffcbf8_ffffca54,
        64'hffffbbe2_ffffbbe2,
        64'hffffbbe2_ffffbbe2,
        64'hffffbbde_ffffbbda,
        64'hffffbbda_ffffbbb6,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_bffe4d62,
        64'h00000000_bffe4b04,
        64'h00000000_bffe4ef4,
        64'h00646374_65675f63,
        64'h6d6d5f64_72616f62,
        64'h00000002_0000ffff,
        64'h004c4b40_004c4b40,
        64'h00300000_20000000,
        64'h00000000_bffe9c88,
        64'h00000000_bffeafc8,
        64'h00717269_5f646e65,
        64'h5f617461_645f6473,
        64'h5f637369_72776f6c,
        64'h00000000_00007172,
        64'h695f646d_635f6473,
        64'h5f637369_72776f6c,
        64'h00007172_695f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0067616c,
        64'h665f7470_75727265,
        64'h746e695f_74696177,
        64'h5f637369_72776f6c,
        64'h00000000_646d635f,
        64'h74726174_735f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0000006e,
        64'h655f7172_695f6473,
        64'h00000000_00007475,
        64'h6f656d69_745f6473,
        64'h00000000_0000657a,
        64'h69736b6c_625f6473,
        64'h00000000_00000074,
        64'h6e636b6c_625f6473,
        64'h00000000_00000000,
        64'h74657365_725f6473,
        64'h00000000_74726174,
        64'h735f646d_635f6473,
        64'h00000000_0000676e,
        64'h69747465_735f6473,
        64'h00000000_00007669,
        64'h645f6b6c_635f6473,
        64'h00000000_00000000,
        64'h6e67696c_615f6473,
        64'h00000000_00006465,
        64'h6c5f7465_735f6473,
        64'h5f637369_72776f6c,
        64'h09020b04_0d060f08,
        64'h010a030c_050e0700,
        64'h020f0c09_0603000d,
        64'h0a070401_0e0b0805,
        64'h0c07020d_08030e09,
        64'h040f0a05_000b0601,
        64'heb86d391_2ad7d2bb,
        64'hbd3af235_f7537e82,
        64'h4e0811a1_a3014314,
        64'hfe2ce6e0_6fa87e4f,
        64'h85845dd1_ffeff47d,
        64'h8f0ccc92_655b59c3,
        64'hfc93a039_ab9423a7,
        64'h432aff97_f4292244,
        64'hc4ac5665_1fa27cf8,
        64'he6db99e5_d9d4d039,
        64'h04881d05_d4ef3085,
        64'heaa127fa_289b7ec6,
        64'hbebfbc70_f6bb4b60,
        64'h4bdecfa9_a4beea44,
        64'hfde5380c_6d9d6122,
        64'h8771f681_fffa3942,
        64'h8d2a4c8a_676f02d9,
        64'hfcefa3f8_a9e3e905,
        64'h455a14ed_f4d50d87,
        64'hc33707d6_21e1cde6,
        64'he7d3fbc8_d8a1e681,
        64'h02441453_d62f105d,
        64'he9b6c7aa_265e5a51,
        64'hc040b340_f61e2562,
        64'h49b40821_a679438e,
        64'hfd987193_6b901122,
        64'h895cd7be_ffff5bb1,
        64'h8b44f7af_698098d8,
        64'hfd469501_a8304613,
        64'h4787c62a_f57c0faf,
        64'hc1bdceee_242070db,
        64'he8c7b756_d76aa478,
        64'h02020202_02020202,
        64'h10020202_02020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02010101_01010101,
        64'h10010101_01010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h08101010_10020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02424242_42424210,
        64'h10101010_10010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h01414141_41414110,
        64'h10101010_10100404,
        64'h04040404_04040404,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h08080808_08080808,
        64'h08080808_08080808,
        64'h08082828_28282808,
        64'h08080808_08080808,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_bf5dd15f,
        64'hf0eff9bf_b0ef12e5,
        64'h05130000_2517b7e1,
        64'he2af80ef_fadfb0ef,
        64'h13050513_00002517,
        64'hbfe9c3df_f0effbff,
        64'hb0ef1325_05130000,
        64'h2517b7f5_e21ff0ef,
        64'h8522fd3f_b0ef1365,
        64'h05130000_2517a001,
        64'ha6dfe0ef_8522fe7f,
        64'hb0ef13a5_05130000,
        64'h25178782_97ba439c,
        64'h97ba078a_6a470713,
        64'h00000717_02f76463,
        64'h47190054_579b0ff4,
        64'h7413fd39_1be3816f,
        64'hc0ef2581_8552688c,
        64'h0004b823_824fc0ef,
        64'h86222401_25816080,
        64'h608ce09c_09058556,
        64'h0007c783_016907b3,
        64'h499117aa_0a130000,
        64'h2a1716aa_8a930000,
        64'h2a974000_04b7286b,
        64'h0b130000_2b174901,
        64'hdfcf80ef_fe9416e3,
        64'h868fc0ef_0405854a,
        64'h0004059b_639097ce,
        64'h00341793_449518e9,
        64'h09130000_29174000,
        64'h09b74401_9d9fe0ef,
        64'h19050513_00002517,
        64'h9b3fe0ef_e05ae456,
        64'he852ec4e_f04af426,
        64'hf822fc06_71399fbf,
        64'he06f2525_05130000,
        64'h25178082_61256be2,
        64'h7b027aa2_7a4279e2,
        64'h690664a6_644660e6,
        64'hb43fe0ef_fd4415e3,
        64'h8d8fc0ef_9456855a,
        64'hff7494e3_8e4fc0ef,
        64'h854ef0df_f0ef0485,
        64'h45890007_c50397ca,
        64'h009407b3_44818fef,
        64'hc0ef854e_f27ff0ef,
        64'h0004051b_45a10100,
        64'h0a370010_0ab7e2eb,
        64'h0b130000_2b174bc1,
        64'h097e2ca9_89930000,
        64'h19974401_4905fa94,
        64'h18e30421_ff579ae3,
        64'h070537e1_00d70023,
        64'h00f556b3_03800793,
        64'h8722f21f_f0ef454d,
        64'h45894601_0034f2df,
        64'hf0efc63e_c43a454d,
        64'h45894601_00340587,
        64'he7930127_67330147,
        64'h87bb0187_571b0087,
        64'h979b00f9_873b0004,
        64'h079b04e2_5ae1b000,
        64'h0a373009_091380b0,
        64'h09b7047e_ec5ef05a,
        64'hec86f456_f852fc4e,
        64'h08100493_69054405,
        64'he0cae4a6_e8a2711d,
        64'hab7fe06f_014160a2,
        64'h64020004_4503943e,
        64'h2a878793_00002797,
        64'h883dfedf_f0ef0045,
        64'h551b35fd_00b7d763,
        64'h842a4785_e406e022,
        64'h1141bfc1_f6180785,
        64'h00076703_97360027,
        64'h97138082_73884000,
        64'h07b7ffe5_37fdc319,
        64'h8b097a98_400006b7,
        64'h3e800793_00b76f63,
        64'h0007871b_40000637,
        64'h47812581_f7884000,
        64'h07b78d51_0106161b,
        64'h8d5d0085_979b8082,
        64'h25017b88_400007b7,
        64'h80822501_6b880007,
        64'hb8234000_07b78082,
        64'h25016388_400007b7,
        64'h8082e388_400007b7,
        64'h91011502_bff1f5df,
        64'hf0ef4541_f63ff0ef,
        64'h4521f69f_f0ef4511,
        64'hf6fff0ef_4509f75f,
        64'hf0ef4505_f7bff0ef,
        64'h4501e406_1141bf51,
        64'hc00028f3_c02026f3,
        64'hfac710e3_a94fc06f,
        64'h33850513_00002517,
        64'h02a74733_02a767b3,
        64'h02b345bb_02c74733,
        64'h40000593_02a68733,
        64'h411686b3_3e800513,
        64'hc00026f3_8e15c020,
        64'h267302b7_1d632705,
        64'hfe0813e3_97aa387d,
        64'h00078023_97aa0007,
        64'h802397aa_00078023,
        64'h97aa0007_80234000,
        64'h081387f2_45a901f6,
        64'h1e134681_48814701,
        64'h00c5131b_46058082,
        64'h80826145_69a26942,
        64'h64e27402_70a2ff24,
        64'h17e3e73f_f0ef2405,
        64'h01358533_46054685,
        64'h008495b3_497901f4,
        64'h99934441_b34fc0ef,
        64'h44850525_05130000,
        64'h2517b42f_c0ef39e5,
        64'h05130000_2517b4ef,
        64'hc0ef37a5_05130000,
        64'h2517b5af_c0ef35e5,
        64'h05130000_25170400,
        64'h0593cb7f_e0efe44e,
        64'he84aec26_f022f406,
        64'h36050513_00002517,
        64'h7179bf89_0485b86f,
        64'hc0ef0a25_05130000,
        64'h2517b7d1_4a89b96f,
        64'hc0ef3725_05130000,
        64'h25179782_852295a2,
        64'h00495613_00195593,
        64'h008a3783_bb4fc0ef,
        64'h38850513_00002517,
        64'hc985000a_358302f7,
        64'h4c636722_010a2783,
        64'hbd0fc0ef_856ee129,
        64'h952ff0ef_85226582,
        64'hbe0fc0ef_856a85e6,
        64'hbe8fc0ef_8562beef,
        64'hc0ef855e_85ce0009,
        64'h8663bfaf_c0ef855a,
        64'h85a68082_61096de2,
        64'h7d027ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_85567446,
        64'h70e6c22f_c0ef4065,
        64'h05130000_25170299,
        64'hf863d7aa_0a130000,
        64'h3a17412d_8d930000,
        64'h2d97412d_0d130000,
        64'h2d1740ac_8c930000,
        64'h2c9740ac_0c130000,
        64'h2c1740ab_8b930000,
        64'h2b9740ab_0b130000,
        64'h2b174485_4a81e03e,
        64'h00395793_c74fc0ef,
        64'he436fc86_ec6ef06a,
        64'hf466f862_fc5ee0da,
        64'he4d6e8d2_f4a64165,
        64'h05130000_251785aa,
        64'h842a892e_962af0ca,
        64'hf8a2fff5_861389b2,
        64'hecce7119_80826505,
        64'hbfb1547d_bf050d85,
        64'hf0bfe0ef_0007c503,
        64'h97ea8b8d_00078b1b,
        64'h001b079b_f1ffe0ef,
        64'h4521ef91_0ba1033d,
        64'hf7b3ff97_95e300d6,
        64'h102392c1_16c20789,
        64'h00fb8633_0006d683,
        64'h018786b3_4781e288,
        64'he6a7b023_00003797,
        64'h8d4166e2_91011402,
        64'h15028c51_0106161b,
        64'h8d5d0105_151b6642,
        64'h67a2886f_e0efe42a,
        64'h88cfe0ef_e82a892f,
        64'he0ef842a_898fe0ef,
        64'hec36b775_4a058082,
        64'h61497da2_7d427ce2,
        64'h6c066ba6_6b466ae6,
        64'h7a0679a6_794674e6,
        64'h640a60aa_8522d56f,
        64'hc0ef4da5_05130000,
        64'h251702fa_18638aa6,
        64'h8bca4785_ed4d842a,
        64'ha94ff0ef_854a85a6,
        64'h866e04fd_966396d6,
        64'h003d9693_67824d81,
        64'h898d0d13_00003d17,
        64'h9c498993_4ca1efec,
        64'h0c130000_3c174b01,
        64'h4a098ba6_ff7fe0ef,
        64'h8acae032_f46ee122,
        64'he506f86a_fc66e0e2,
        64'he4dee8da_ecd6f0d2,
        64'h69850200_051384ae,
        64'h892af4ce_f8cafca6,
        64'h7175bfb1_547dbf05,
        64'h0d8582cf_f0ef0007,
        64'hc50397ea_8b8d0007,
        64'h8b1b001b_079b840f,
        64'hf0ef4521_ef910ba1,
        64'h033df7b3_ff9795e3,
        64'h00d60023_0ff6f693,
        64'h078500fb_86330006,
        64'hc6830187_86b34781,
        64'he288f6a7_bd230000,
        64'h37978d41_66e29101,
        64'h14021502_8c510106,
        64'h161b8d5d_0105151b,
        64'h664267a2_9a8fe0ef,
        64'he42a9aef_e0efe82a,
        64'h9b4fe0ef_842a9baf,
        64'he0efec36_b7754a05,
        64'h80826149_7da27d42,
        64'h7ce26c06_6ba66b46,
        64'h6ae67a06_79a67946,
        64'h74e6640a_60aa8522,
        64'he78fc0ef_5fc50513,
        64'h00002517_02fa1863,
        64'h8aa68bca_4785ed4d,
        64'h842abb6f_f0ef854a,
        64'h85a6866e_04fd9663,
        64'h96d6003d_96936782,
        64'h4d819bad_0d130000,
        64'h3d179c49_89934ca1,
        64'h018c0c13_00003c17,
        64'h4b014a09_8ba6918f,
        64'hf0ef8aca_e032f46e,
        64'he122e506_f86afc66,
        64'he0e2e4de_e8daecd6,
        64'hf0d26985_02000513,
        64'h84ae892a_f4cef8ca,
        64'hfca67175_b7e95b7d,
        64'hb7490605_00b83023,
        64'he30c85d6_e11185e2,
        64'h00167513_80826109,
        64'h6de27d02_7ca27c42,
        64'h7be26b06_6aa66a46,
        64'h69e67906_74a6855a,
        64'h744670e6_f2cfc0ef,
        64'h68850513_00002517,
        64'hfafb90e3_04000793,
        64'h2b85fbb4_1be38c56,
        64'h2405e931_8b2ac72f,
        64'hf0ef854a_85ce6622,
        64'hf58fc0ef_856a85da,
        64'hf60fc0ef_e4328552,
        64'h06f61063_974e00e9,
        64'h08330036_17136782,
        64'h4601fffc_4a93f7ef,
        64'hc0ef8566_85da0084,
        64'h8b3bf8af_c0ef8552,
        64'h4401003b_949b0177,
        64'h9c334785_4da168ed,
        64'h0d130000_2d17686c,
        64'h8c930000_2c9767ea,
        64'h0a130000_2a17fb6f,
        64'hc0ef4b81_e03289ae,
        64'hf862e0da_e4d6f4a6,
        64'hf8a2fc86_ec6ef06a,
        64'hf466fc5e_e8d2ecce,
        64'h69850513_00002517,
        64'h892af0ca_7119bf75,
        64'h5dfdbfc5_859afe08,
        64'h0be385ba_b7610605,
        64'he10ce28c_85c60008,
        64'h036385be_008bea63,
        64'h00167813_80826109,
        64'h6de27d02_7ca27c42,
        64'h7be26b06_6aa66a46,
        64'h69e67906_74a6856e,
        64'h744670e6_82dfc0ef,
        64'h78850513_00002517,
        64'hf8f41be3_08000793,
        64'h2405ed29_8daad6af,
        64'hf0ef8526_85ca6622,
        64'h851fc0ef_856685a2,
        64'h859fc0ef_e432854e,
        64'h05461c63_96ca00d4,
        64'h85330036_16934601,
        64'hfff7c893_fff74313,
        64'h8fd5008d_16b300fd,
        64'h17b30024_079b8f5d,
        64'h00ed1733_00fd17b3,
        64'h408b07bb_408a873b,
        64'h899fc0ef_856285a2,
        64'h8a1fc0ef_854e796c,
        64'h8c930000_2c9703f0,
        64'h0b930810_0b134d05,
        64'h07f00a93_79cc0c13,
        64'h00002c17_79498993,
        64'h00002997_8cdfc0ef,
        64'h44018a32_892eec6e,
        64'hfc86f06a_f466f862,
        64'hfc5ee0da_e4d6e8d2,
        64'heccef0ca_f8a27ae5,
        64'h05130000_251784aa,
        64'hf4a67119_b7f15dfd,
        64'hbfe5e19c_e31cbf61,
        64'h0605e194_e314008c,
        64'h66638082_61096de2,
        64'h7d027ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_856e7446,
        64'h70e6933f_c0ef88e5,
        64'h05130000_3517fb54,
        64'h17e32405_e1398daa,
        64'he6cff0ef_852685ca,
        64'h6622953f_c0ef856a,
        64'h85a295bf_c0efe432,
        64'h85520566_1a63974a,
        64'h00e485b3_00361713,
        64'h4601fff6_c693fff7,
        64'hc7930089_96b300f9,
        64'h97b3408b_87bb987f,
        64'hc0ef8566_85a298ff,
        64'hc0ef8552_08000a93,
        64'h888d0d13_00003d17,
        64'h03f00c13_498507f0,
        64'h0b9388ac_8c930000,
        64'h3c97882a_0a130000,
        64'h3a179bbf_c0ef4401,
        64'h8b32892e_ec6efc86,
        64'hf06af466_f862fc5e,
        64'he0dae4d6_e8d2ecce,
        64'hf0caf8a2_89c50513,
        64'h00003517_84aaf4a6,
        64'h7119b7f1_5dfdbfe5,
        64'he298e398_bf610605,
        64'he28ce38c_008c6663,
        64'h80826109_6de27d02,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e67906,
        64'h74a6856e_744670e6,
        64'ha21fc0ef_97c50513,
        64'h00003517_fb541be3,
        64'h2405e139_8daaf5af,
        64'hf0ef8526_85ca6622,
        64'ha41fc0ef_856a85a2,
        64'ha49fc0ef_e4328552,
        64'h05661a63_97ca00f4,
        64'h86b30036_17934601,
        64'h008995b3_00e99733,
        64'h408b873b_a6dfc0ef,
        64'h856685a2_a75fc0ef,
        64'h85520800_0a9396ed,
        64'h0d130000_3d1703f0,
        64'h0c134985_07f00b93,
        64'h970c8c93_00003c97,
        64'h968a0a13_00003a17,
        64'haa1fc0ef_44018b32,
        64'h892eec6e_fc86f06a,
        64'hf466f862_fc5ee0da,
        64'he4d6e8d2_eccef0ca,
        64'hf8a29825_05130000,
        64'h351784aa_f4a67119,
        64'hbff159fd_b74d0605,
        64'he29ce31c_80826125,
        64'h6c426be2_7b027aa2,
        64'h7a4279e2_690664a6,
        64'h854e6446_60e6af7f,
        64'hc0efa525_05130000,
        64'h3517f94c_19e30c05,
        64'he91d89aa_831ff0ef,
        64'h852285a6_6622b17f,
        64'hc0ef855e_85ceb1ff,
        64'hc0efe432_854a0556,
        64'h17639726_00e406b3,
        64'h00361713_46018fd9,
        64'h038c1713_8fd9030c,
        64'h17138fd9_028c1713,
        64'h8fd9020c_17138fd9,
        64'h018c1713_0187e7b3,
        64'h8fd9008c_1793010c,
        64'h1713b63f_c0ef855a,
        64'h85ce000c_099bb6ff,
        64'hc0ef854a_10000a13,
        64'ha68b8b93_00003b97,
        64'ha60b0b13_00003b17,
        64'ha5890913_00003917,
        64'hb91fc0ef_4c018ab2,
        64'h84aefc4e_ec86e862,
        64'hec5ef05a_f456f852,
        64'he0cae4a6_a6c50513,
        64'h00003517_842ae8a2,
        64'h711db7e1_5d7db779,
        64'h0605e198_e398872a,
        64'hc291876a_00167693,
        64'hbf49000b_3d038082,
        64'h61656d42_6ce27c02,
        64'h7ba27b42_7ae26a06,
        64'h69a66946_64e6856a,
        64'h740670a6_bf5fc0ef,
        64'hb5050513_00003517,
        64'hfb441ae3_2405e529,
        64'h8d2a92ff_f0ef8526,
        64'h85ca6622_c15fc0ef,
        64'h856685a2_c1dfc0ef,
        64'he432854e_05561c63,
        64'h97ca00f4_85b30036,
        64'h1793fffd_45134601,
        64'hc39fc0ef_856285a2,
        64'h000bbd03_cba50014,
        64'h7793c4bf_c0ef854e,
        64'h04000a13_b44c8c93,
        64'h00003c97_b3cc0c13,
        64'h00003c17_e3cb8b93,
        64'h00003b97_e3cb0b13,
        64'h00003b17_b4498993,
        64'h00003997_c7dfc0ef,
        64'h44018ab2_892ee86a,
        64'hf486ec66_f062f45e,
        64'hf85afc56_e0d2e4ce,
        64'he8caf0a2_b5c50513,
        64'h00003517_84aaeca6,
        64'h7159bfc1_54fdbf59,
        64'h0605e198_e3988726,
        64'hc2918766_00167693,
        64'h80826165_6ce27c02,
        64'h7ba27b42_7ae26a06,
        64'h69a664e6_69468526,
        64'h740670a6_cddfc0ef,
        64'hc3850513_00003517,
        64'hfb541be3_2405e129,
        64'h84aaa17f_f0ef854a,
        64'h85ce6622_cfdfc0ef,
        64'h856285a2_d05fc0ef,
        64'he4328552_05661863,
        64'h97ce00f9_05b30036,
        64'h179314fd_46014090,
        64'h0cb3d23f_c0ef8885,
        64'h855e85a2_fff44493,
        64'hd31fc0ef_85520400,
        64'h0a93c2ac_0c130000,
        64'h3c17c22b_8b930000,
        64'h3b97c1aa_0a130000,
        64'h3a17d53f_c0ef4401,
        64'h8b3289ae_ec66eca6,
        64'hf486f062_f45ef85a,
        64'hfc56e0d2_e4cef0a2,
        64'hc3050513_00003517,
        64'h892ae8ca_7159bfc9,
        64'h070500a8_3023e288,
        64'h00f70533_ab1ff06f,
        64'h6121863a_69e2854e,
        64'h790274a2_70e27442,
        64'h00c71c63_96ae00d9,
        64'h88330037_16934701,
        64'h8fc59081_178265a2,
        64'h66021482_8fc18cc9,
        64'h0109179b_0105151b,
        64'h935fe0ef_84aa93bf,
        64'he0ef892a_941fe0ef,
        64'h842a947f_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7f100e8_30238f69,
        64'h00083703_e3148ee9,
        64'h07856314_b29ff06f,
        64'h6121863e_69e2854e,
        64'h790274a2_70e27442,
        64'h00c79c63_974e00e5,
        64'h88330037_97134781,
        64'h8d5d9101_178265a2,
        64'h66021502_8fc18d45,
        64'h0109179b_0105151b,
        64'h9adfe0ef_84aa9b3f,
        64'he0ef892a_9b9fe0ef,
        64'h842a9bff_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7f100e8_30238f49,
        64'h00083703_e3148ec9,
        64'h07856314_ba1ff06f,
        64'h6121863e_69e2854e,
        64'h790274a2_70e27442,
        64'h00c79c63_974e00e5,
        64'h88330037_97134781,
        64'h8d5d9101_178265a2,
        64'h66021502_8fc18d45,
        64'h0109179b_0105151b,
        64'ha25fe0ef_84aaa2bf,
        64'he0ef892a_a31fe0ef,
        64'h842aa37f_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7d100e8_302302a7,
        64'h57330008_3703e314,
        64'h02a6d6b3_07856314,
        64'h4505e111_c21ff06f,
        64'h6121863e_69e2854e,
        64'h790274a2_70e27442,
        64'h00c79c63_974e00e5,
        64'h88330037_97134781,
        64'h8d5d9101_178265a2,
        64'h66021502_8fc18d45,
        64'h0109179b_0105151b,
        64'haa5fe0ef_84aaaabf,
        64'he0ef892a_ab1fe0ef,
        64'h842aab7f_e0ef89aa,
        64'hec4ef04a_f426f822,
        64'hfc06e032_e42e7139,
        64'hb7e100e8_302302a7,
        64'h07330008_3703e314,
        64'h02a686b3_07856314,
        64'hc9dff06f_6121863e,
        64'h69e2854e_790274a2,
        64'h70e27442_00c79c63,
        64'h974e00e5_88330037,
        64'h97134781_8d5d9101,
        64'h178265a2_66021502,
        64'h8fc18d45_0109179b,
        64'h0105151b_b21fe0ef,
        64'h84aab27f_e0ef892a,
        64'hb2dfe0ef_842ab33f,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7f100e8,
        64'h30238f09_00083703,
        64'he3148e89_07856314,
        64'hd15ff06f_6121863e,
        64'h69e2854e_790274a2,
        64'h70e27442_00c79c63,
        64'h974e00e5_88330037,
        64'h97134781_8d5d9101,
        64'h178265a2_66021502,
        64'h8fc18d45_0109179b,
        64'h0105151b_b99fe0ef,
        64'h84aab9ff_e0ef892a,
        64'hba5fe0ef_842ababf,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7f100e8,
        64'h30238f29_00083703,
        64'he3148ea9_07856314,
        64'hd8dff06f_6121863e,
        64'h69e2854e_790274a2,
        64'h70e27442_00c79c63,
        64'h974e00e5_88330037,
        64'h97134781_8d5d9101,
        64'h178265a2_66021502,
        64'h8fc18d45_0109179b,
        64'h0105151b_c11fe0ef,
        64'h84aac17f_e0ef892a,
        64'hc1dfe0ef_842ac23f,
        64'he0ef89aa_ec4ef04a,
        64'hf426f822_fc06e032,
        64'he42e7139_b7ad0485,
        64'hb23ff0ef_0007c503,
        64'h97e20039_f7930985,
        64'hb33ff0ef_4521ef81,
        64'h00adb023_00acb023,
        64'h8d419101_14021502,
        64'h01a46433_00a96533,
        64'h010d1d1b_0105151b,
        64'h0344f7b3_c79fe0ef,
        64'h892ac7ff_e0ef8d2a,
        64'hc85fe0ef_842ac8bf,
        64'he0efe47f_f06f6165,
        64'h7ae28556_7b4264e6,
        64'h85da8626_6da26d42,
        64'h6ce27c02_7ba26a06,
        64'h69a66946_70a67406,
        64'h948fd0ef_0cc50513,
        64'h00003517_03749b63,
        64'h00fb0cb3_00fa8db3,
        64'h00349793_474c0c13,
        64'h00003c17_9c4a0a13,
        64'h4981bc5f_f0ef4481,
        64'h8bb28b2e_e46ee86a,
        64'hec66e8ca_f0a2f486,
        64'hf062f45e_f85ae4ce,
        64'heca60200_05138aaa,
        64'h6a05fc56_e0d27159,
        64'hb75107a1_05858082,
        64'h61616ba2_6b426ae2,
        64'h7a0279a2_794274e2,
        64'h640660a6_557d9bef,
        64'hd0ef0fa5_05130000,
        64'h35179caf_d0ef0ce5,
        64'h05130000_3517058e,
        64'h02d60b63_fff7c693,
        64'hc31986be_8b056390,
        64'h00858733_bf6d07a1,
        64'h07056394_e390fff7,
        64'hc613c299_863e8a85,
        64'h008706b3_a0a94501,
        64'ha08fd0ef_16450513,
        64'h00003517_fd4417e3,
        64'h04050325_99634581,
        64'h87a6a22f_d0ef855a,
        64'h85dea2af_d0ef854e,
        64'h03271863_470187a6,
        64'ha38fd0ef_855685de,
        64'h00040b9b_a44fd0ef,
        64'h854e4a41_13cb0b13,
        64'h00003b17_134a8a93,
        64'h00003a97_12c98993,
        64'h00003997_a64fd0ef,
        64'h4401892e_e45ee486,
        64'he85aec56_f052f44e,
        64'hf84ae0a2_13c50513,
        64'h00003517_84aafc26,
        64'h715dbf5d_0785a001,
        64'ha90fd0ef_13c50513,
        64'h00003517_85a28626,
        64'haa0fd0ef_12450513,
        64'h00003517_6090600c,
        64'h02e80363_60980004,
        64'h38038082_61054501,
        64'h64a26442_60e200c7,
        64'h986300d5_043300d5,
        64'h84b30037_96934781,
        64'he426e822_ec061101,
        64'hc2dff06f_80824501,
        64'h80824501_80828082,
        64'h80828082_45098082,
        64'h45098082_4509bff9,
        64'h26052004_04136622,
        64'hea3fc0ef_e4328522,
        64'h85b28082_61454501,
        64'h64e27402_70a20096,
        64'h186300c6_84bb842e,
        64'hf406ec26_f0227179,
        64'h80824505_80824505,
        64'h80824505_80820141,
        64'h8d7d6402_60a29522,
        64'h408007b3_f57ff0ef,
        64'he406952e_842ae022,
        64'h1141a001_d2dff0ef,
        64'h4505b62f_d0efe406,
        64'h1b050513_00003517,
        64'h85aa862e_86b28736,
        64'h11418082_02f55533,
        64'h47a9b000_25738082,
        64'h45018082_45018082,
        64'h01414501_60a2f51f,
        64'hc0ef2000_0537b9ef,
        64'hd0efe406_1c450513,
        64'h00003517_11418082,
        64'h80826105_644260e2,
        64'h85229daf_f0ef4581,
        64'h6622c509_842afd1f,
        64'hf0efe432_8532ec06,
        64'he8221101_02b50633,
        64'h8082953e_055e10d0,
        64'h0513e308_95360017,
        64'h86930075_6513157d,
        64'h631cafa7_07130000,
        64'h47178082_45018082,
        64'h24050513_000f4537,
        64'ha001ddbf_f0efe406,
        64'h25011141_90020000,
        64'h0023e8df_f0efc1ef,
        64'hd0ef9fa5_05130000,
        64'h3517bddd_c2cfd0ef,
        64'h22850513_00003517,
        64'hc981c62e_0005059b,
        64'h8d6f90ef_01849513,
        64'h85a2c4af_d0ef22e5,
        64'h05130000_3517c56f,
        64'hd0ef1f25_05130000,
        64'h351785a2_01849613,
        64'h86a20bf0_0493bf1d,
        64'h1f050513_00003517,
        64'hc5112501_d79fa0ef,
        64'h4501efa5_85930000,
        64'h35974605_bf911de5,
        64'h05130000_3517bfb9,
        64'h20050513_00003517,
        64'hc9192501_c6efb0ef,
        64'h54020808_f3f99cbd,
        64'h47b225a0_10ef854e,
        64'hdbfff0ef_00044503,
        64'h9452dc9f_f0ef880d,
        64'h45210004_099b00c4,
        64'hd41be505_2501fbbf,
        64'ha0ef0808_95ca6605,
        64'h00749181_02049593,
        64'h300a0a13_00003a17,
        64'h09620bf0_0913e12d,
        64'h44812501_e53fa0ef,
        64'h08082425_85930000,
        64'h35974605_d0cfd0ef,
        64'h23050513_00003517,
        64'h80822701_01132401,
        64'h3a032481_39832501,
        64'h39032581_34832601,
        64'h34032681_3083d36f,
        64'hd0ef23a5_05130000,
        64'h3517c515_2501e43f,
        64'ha0ef2541_30232531,
        64'h34232521_38232491,
        64'h3c232681_30232611,
        64'h3423c725_05130000,
        64'h4517fe25_85930000,
        64'h35974605_d9010113,
        64'h8302037e_c4458593,
        64'h00002597_4305f140,
        64'h25730ff0_000f0000,
        64'h100f8082_610560e2,
        64'he9fff0ef_00914503,
        64'hea7ff0ef_00814503,
        64'hf13ff0ef_ec06002c,
        64'h11018082_61456942,
        64'h64e27402_70a2fe94,
        64'h10e3ec9f_f0ef0091,
        64'h4503ed1f_f0ef3461,
        64'h00814503_f3fff0ef,
        64'h0ff57513_002c0089,
        64'h553354e1_03800413,
        64'h892af406_e84aec26,
        64'hf0227179_80826145,
        64'h694264e2_740270a2,
        64'hfe9410e3_f0bff0ef,
        64'h00914503_f13ff0ef,
        64'h34610081_4503f81f,
        64'hf0ef0ff5_7513002c,
        64'h0089553b_54e14461,
        64'h892af406_e84aec26,
        64'hf0227179_80826105,
        64'h644260e2_f43ff0ef,
        64'h00914503_f4bff0ef,
        64'h00814503_fb7ff0ef,
        64'h0ff47513_002cf5df,
        64'hf0ef0091_4503f65f,
        64'hf0ef0081_4503fd1f,
        64'hf0efec06_8121842a,
        64'h002ce822_11018082,
        64'h00f58023_00e580a3,
        64'h0007c783_00074703,
        64'h97aa973e_811100f5,
        64'h7713d027_87930000,
        64'h2797b7f5_0405fa5f,
        64'hf0ef8082_01416402,
        64'h60a2e509_00044503,
        64'h842ae406_e0221141,
        64'h808200e7_88230200,
        64'h071300e7_8423fc70,
        64'h071300e7_8623470d,
        64'h00078223_00e78023,
        64'h476d00e7_8623f800,
        64'h07130007_82231000,
        64'h07b78082_00a70023,
        64'hdfe50207_f7930147,
        64'h47831000_07378082,
        64'h02057513_0147c503,
        64'h100007b7_80820005,
        64'h45038082_00b50023,
        64'h80826105_690264a2,
        64'h644260e2_f47dfa1f,
        64'hf0ef4124_0433854a,
        64'h89260084_f3638922,
        64'h68048493_842ae04a,
        64'hec06e822_009894b7,
        64'he4261101_80826105,
        64'h690264a2_644260e2,
        64'hfe856ee3_f45ff0ef,
        64'h0405944a_02855433,
        64'h24040413_000f4437,
        64'h02a48533_370000ef,
        64'h892af63f_f0ef84aa,
        64'he04ae426_e822ec06,
        64'h11018082_02a7d533,
        64'h01419101_15026402,
        64'h60a202f4_07b32407,
        64'h8793000f_47b73a20,
        64'h00ef842a_f95ff0ef,
        64'he022e406_11418082,
        64'h610564a2_8d0502a7,
        64'hd5336442_60e29101,
        64'h150202f4_07b33e80,
        64'h07933ce0_00ef842a,
        64'hfc1ff0ef_84aae426,
        64'he822ec06_11018082,
        64'h45018082_01418d5d,
        64'h91011782_150260a2,
        64'h1007e783_10a7a223,
        64'h10e1a023_27051001,
        64'ha70300e5_7763878e,
        64'h1041e703_492000ef,
        64'he4061141_8082cf3f,
        64'hf06fd0a5_85930000,
        64'h45974611_cb81f227,
        64'hd7830000_47978082,
        64'h24010113_22013903,
        64'h22813483_23013403,
        64'h23813083_f63ff0ef,
        64'h8522002c_ec2ff0ef,
        64'he802c44a_08282040,
        64'h061385a6_e84ff0ef,
        64'h22113c23_00282180,
        64'h06134581_893284ae,
        64'h842a2321_30232291,
        64'h34232281_3823dc01,
        64'h0113ebff_f06f6145,
        64'h05c170a2_41907402,
        64'hd8dff06f_614570a2,
        64'h65a27402_85228a7f,
        64'hd0efe42e_57450513,
        64'h00003517_842a8b7f,
        64'hd06f6145_59c50513,
        64'h00003517_70a27402,
        64'h02f70a63_478d00d7,
        64'h0e6301e1_570300e1,
        64'h0f230115_c70300e1,
        64'h0fa34689_0105c703,
        64'hf022f406_71798082,
        64'h61056902_64a26442,
        64'h60e2d5ff_f06f6105,
        64'h690264a2_60e26442,
        64'h909fd0ef_5bc50513,
        64'h00003517_0087cf63,
        64'h278d439c_00c78793,
        64'h00004797_00f71c23,
        64'h00004717_27850007,
        64'hd7830267_87930000,
        64'h47972400_00ef0200,
        64'h0513d33f_f0ef4515,
        64'h03c5d583_00004597,
        64'h256000ef_4535e2bf,
        64'hf0ef854a_e4458593,
        64'h00004597_e4a79723,
        64'h00004797_4611d25f,
        64'hf0ef0665_55030000,
        64'h4517e6a7_91230000,
        64'h4797d39f_f0ef4511,
        64'hdc1ff0ef_00448513,
        64'hffc4059b_06a79a63,
        64'h25010024_d783d55f,
        64'hf0ef0965_55030000,
        64'h451708a7_95632501,
        64'h0004d783_d6bff0ef,
        64'h84ae450d_892a08c7,
        64'hdf638432_478de04a,
        64'he426ec06_e8221101,
        64'hb7990c87_93230000,
        64'h4797eaff_f0ef854e,
        64'hec858593_00004597,
        64'h4611eca7_9a230000,
        64'h4797da9f_f0ef4501,
        64'heea79023_00004797,
        64'hdb7ff0ef_10f73223,
        64'h00004717_10f73223,
        64'h00004717_451101f4,
        64'h17934405_a1dfd0ef,
        64'h6b050513_00003517,
        64'h858a4390_11c78793,
        64'h00004797_e1cff0ef,
        64'h850a85a2_e24ff0ef,
        64'h850a6ca5_85930000,
        64'h359700f7_096302f0,
        64'h07930129_4703e10f,
        64'hf0ef850a_4d458593,
        64'h00003597_885ff0ef,
        64'h850a4581_10000613,
        64'hb75516f7_21230000,
        64'h47172000_07938082,
        64'h615569b2_695264f2,
        64'h741270b2_a8dfd0ef,
        64'h6f850513_00003517,
        64'h00a405b3_f4cff0ef,
        64'h51850513_00003517,
        64'h842af5af_f0ef8522,
        64'h04a7f263_0ff00793,
        64'h9526f6af_f0ef5365,
        64'h05130000_351784aa,
        64'hf78ff0ef_85221aa7,
        64'haf230000_479704e7,
        64'hee631ff0_0793fff5,
        64'h071beabf_f0ef9526,
        64'h0505f9af_f0ef8526,
        64'h00a404b3_0505fa6f,
        64'hf0ef892e_ea4aee26,
        64'hf6068522_89aae64e,
        64'h01258413_f2227169,
        64'h80824501_80820141,
        64'h640260a2_8522547d,
        64'h00850363_830fa0ef,
        64'h8432e406_e0221141,
        64'h83026105_25011fe5,
        64'h85930000_25976902,
        64'h834a64a2_60e26442,
        64'hf1402573_0ff0000f,
        64'h0000100f_b55fd0ef,
        64'h7a850513_00003517,
        64'h862286aa_608ce41f,
        64'hc0ef85a2_6088b6ff,
        64'hd0ef85a2_4124043b,
        64'hec067b25_05130000,
        64'h35170004_b9036380,
        64'he04ae822_28448493,
        64'h00004497_29478793,
        64'h00004797_e4261101,
        64'h80826105_64a26442,
        64'he00c95a6_60e2600c,
        64'ha1fff0ef_ec066008,
        64'h85aa84ae_862ee426,
        64'h2c040413_00004417,
        64'he8221101_80822cf7,
        64'h37230000_47172cf7,
        64'h37230000_471707fe,
        64'h47854e80_006f0305,
        64'h05130141_60a26402,
        64'h02a4753b_4529fe7f,
        64'hf0ef357d_02b455bb,
        64'h45a900b7_f86347a5,
        64'h00a04563_842ee406,
        64'he0221141_b7c50505,
        64'hfd07879b_9fb902f6,
        64'h07bb00b6_e763fd07,
        64'h059b2701_8082853e,
        64'he3190005_47034629,
        64'h46a54781_80820141,
        64'h91411542_11418d5d,
        64'h05220085_579bfa5f,
        64'hf06f4581_d7dff06f,
        64'h01410505_45814629,
        64'h60a26402_f77d8b11,
        64'h00074703_973e0005,
        64'h4703fea4_7ae3157d,
        64'h80820141_557d6402,
        64'h60a2e719_8b110007,
        64'h4703973e_fff58513,
        64'hd9878793_00002797,
        64'hfff5c703_00a405b3,
        64'h951ff0ef_e589842a,
        64'he406e022_1141bfd5,
        64'h0789bff1_052a052a,
        64'hb7e9e01c_078d00e6,
        64'h98630420_07130027,
        64'hc683fce6_9fe3052a,
        64'h06900713_0017c683,
        64'hfed716e3_06b00693,
        64'h02d70763_04d00693,
        64'h80820141_640260a2,
        64'h02d70e63_04700693,
        64'h00e6ea63_02d70463,
        64'h0007c703_04b00693,
        64'h601cf87f_f0ef842e,
        64'he406e022_1141b7e1,
        64'he008b7cd_fc97879b,
        64'h0ff7f793_fe07079b,
        64'hc6098a09_b7d196be,
        64'h050502d5_86b3feb7,
        64'hf4e3fd07_879b0008,
        64'h8b630046_78938082,
        64'h61058536_644260e2,
        64'hec050008_98630446,
        64'h78930006_460300f8,
        64'h06330007_079b0005,
        64'h4703e728_08130000,
        64'h28174681_00c16583,
        64'he0dff0ef_c632ec06,
        64'h006c842e_e8221101,
        64'hbfd50789_bff1052a,
        64'h052ab7e9_e01c078d,
        64'h00e69863_04200713,
        64'h0027c683_fce69fe3,
        64'h052a0690_07130017,
        64'hc683fed7_16e306b0,
        64'h069302d7_076304d0,
        64'h06938082_01416402,
        64'h60a202d7_0e630470,
        64'h069300e6_ea6302d7,
        64'h04630007_c70304b0,
        64'h0693601c_f0dff0ef,
        64'h842ee406_e0221141,
        64'h80820141_40a00533,
        64'h60a2f23f_f0efe406,
        64'h05051141_f2dff06f,
        64'h00e68463_02d00713,
        64'h00054683_b7e94501,
        64'he088fcf7_18e347a9,
        64'hfd279be3_07858f81,
        64'hcb010007_c703fe87,
        64'h82e367e2_f5dff0ef,
        64'h8522082c_892a862e,
        64'h80826121_790274a2,
        64'h744270e2_5529e901,
        64'h65a2b03f_f0ef84b2,
        64'h842ae42e_00063023,
        64'hf04afc06_f426f822,
        64'h7139b7e1_e008b7cd,
        64'hfc97879b_0ff7f793,
        64'hfe07079b_c6098a09,
        64'hb7d196be_050502d5,
        64'h86b3feb7_f4e3fd07,
        64'h879b0008_8b630046,
        64'h78938082_61058536,
        64'h644260e2_ec050008,
        64'h98630446_78930006,
        64'h460300f8_06330007,
        64'h079b0005_4703fc68,
        64'h08130000_28174681,
        64'h00c16583_f61ff0ef,
        64'hc632ec06_006c842e,
        64'he8221101_8082fae7,
        64'h8fe34741_bfed47a9,
        64'h8082c19c_47a1a809,
        64'h050900e7_9c630780,
        64'h07130ff7_f7930207,
        64'h879bc709_8b050007,
        64'h4703973e_01470713,
        64'h00002717_00154783,
        64'h02f71f63_03000793,
        64'h00054703_c19c47c1,
        64'hcf950447_f7930007,
        64'hc78397ba_00254703,
        64'h04d71763_07800693,
        64'h0ff77713_0207071b,
        64'hc6898a85_0006c683,
        64'h00e786b3_05c78793,
        64'h00002797_00154703,
        64'h06f71e63_03000793,
        64'h00054703_e7c9419c,
        64'hb7f1377d_87aabfa5,
        64'hfef51be3_0785f8b7,
        64'h12e30007_c70300d8,
        64'h0a630087_85130007,
        64'hb803bfcd_367d0785,
        64'hf8b71fe3_0007c703,
        64'hd24d8a1d_eb1187aa,
        64'h27018edd_00365713,
        64'h02079693_8fd90107,
        64'h179300b7_e7330085,
        64'h97938e19_953a9301,
        64'h1702fed8_19e30007,
        64'h869b0785_fcb69de3,
        64'h0007c683_87aa00a7,
        64'h083b9f1d_4721c39d,
        64'h00757793_b7f5367d,
        64'h0785feb7_1ce30007,
        64'hc7038082_853e4781,
        64'he60187aa_260100c7,
        64'hef630ff5_f59347c1,
        64'hb7ed853e_feb70be3,
        64'h00150793_00054703,
        64'h80824501_00c51463,
        64'h0ff5f593_962abfe1,
        64'h0405d17d_f83ff0ef,
        64'h852285ca_86268082,
        64'h614569a2_694264e2,
        64'h740270a2_85224401,
        64'h0097db63_408987bb,
        64'h008509bb_d0dff0ef,
        64'h8522c899_0005049b,
        64'hd19ff0ef_892ee44e,
        64'hf406e84a_ec26852e,
        64'h842af022_7179bfc5,
        64'h0505feb7_8de30005,
        64'h47838082_00c51363,
        64'h962a8082_853ed3f5,
        64'h9f950705_0006c683,
        64'h0007c783_00e586b3,
        64'h00e507b3_a8214781,
        64'h00e61463_4701b7e5,
        64'h00b70023_97220005,
        64'hc58300e6_85b300f8,
        64'h0733fef6_05e317fd,
        64'h4781fff6_461386ae,
        64'h88328082_01416402,
        64'h60a28522_f53ff0ef,
        64'h00a5e963_842ae406,
        64'he0221141_80826145,
        64'h64e26942_85267402,
        64'h70a20004_0023f75f,
        64'hf0ef944a_864a8522,
        64'hfff60913_00c56463,
        64'h6582892a_ce1184aa,
        64'h6622dd3f_f0efe02e,
        64'he84af406_e432ec26,
        64'h852e842a_f0227179,
        64'hb7e50106_80230785,
        64'h00f706b3_0006c803,
        64'h00f586b3_808200f6,
        64'h13634781_00f50733,
        64'h963a95be_078e02e7,
        64'h87335761_00365793,
        64'hfed765e3_40f606b3,
        64'h0106b023_07a100f5,
        64'h06b30006_b80300f5,
        64'h86b3a811_471d4781,
        64'heb9d872a_8b9d00b5,
        64'h67b304b5_0463b7f5,
        64'hfeb78fa3_0785bfe9,
        64'hfee7bc23_07a18082,
        64'h00c79763_963e963a,
        64'h97aa078e_02e78733,
        64'h57610036_57930106,
        64'hee6340f8_8833469d,
        64'h00c508b3_87aaffed,
        64'h8f5537fd_07220ff5,
        64'hf69347a1_eb0587aa,
        64'h00757713_80824501,
        64'hb7e50789_00d780a3,
        64'h00e78023_8082e311,
        64'h0017c703_ce810007,
        64'hc68387aa_cf990005,
        64'h4783c11d_80826105,
        64'h64a28526_644260e2,
        64'he0080505_00050023,
        64'hc501f73f_f0ef8526,
        64'h842ac891_e822ec06,
        64'h6104e426_1101bfd9,
        64'h70a7bc23_00004797,
        64'h05050005_0023c781,
        64'h00054783_c519f9ff,
        64'hf0ef8522_85a68082,
        64'h610564a2_644260e2,
        64'h85224401_7407b223,
        64'h00004797_ef810004,
        64'h4783942a_fa1ff0ef,
        64'h85a68522_cc116380,
        64'h76078793_00004797,
        64'he519842a_84aeec06,
        64'he426e822_1101bfd5,
        64'h87aeb7e5_0505fafd,
        64'h0007c683_0785fee6,
        64'h8fe38082_4501eb19,
        64'h00054703_b7c50785,
        64'h8082853e_fa7d0007,
        64'h46030705_00d60863,
        64'ha021872e_ca890007,
        64'h468300f5_07334781,
        64'hbfd5872e_b7d50785,
        64'hfa7d0007_46030705,
        64'hfed60ee3_8082853e,
        64'hea990007_468300f5,
        64'h07334781_b7fd0785,
        64'h808240a7_8533e701,
        64'h0007c703_00b78563,
        64'h87aa95aa_80826105,
        64'h644260e2_4501fe85,
        64'h7be3157d_00b78663,
        64'h00054783_0ff5f593,
        64'h952265a2_fe5ff0ef,
        64'hec06842a_e42ee822,
        64'h1101bfcd_07858082,
        64'h40a78533_e7010007,
        64'hc70387aa_bfcd0505,
        64'hdffd8082_00b79363,
        64'h00054783_0ff5f593,
        64'h80824501_bfcd0505,
        64'hc3998082_00b79363,
        64'h00054783_0ff5f593,
        64'h8082853e_fee10705,
        64'he3994187_d79b0187,
        64'h979b40f6_87bb0007,
        64'hc78300e5_87b30007,
        64'hc68300e5_07b3a015,
        64'h478100e6_14634701,
        64'h8082853e_f37d0505,
        64'he3994187_d79b0187,
        64'h979b40f7_07bbfff5,
        64'hc7830005_47030585,
        64'h80820007_8023fec7,
        64'h99e3d375_fee78fa3,
        64'h0785fff5_c7030585,
        64'h963efb7d_00178693,
        64'h0007c703_87b68082,
        64'he21987aa_b7d587b6,
        64'h8082fb75_fee78fa3,
        64'h0785fff5_c7030585,
        64'heb090017_86930007,
        64'hc70387aa_8082f76d,
        64'h00e68023_078500f5,
        64'h06b30007_470300f5,
        64'h873300c7_8c634781,
        64'h8082fb75_fee78fa3,
        64'h0785fff5_c7030585,
        64'h87aa8082_01416402,
        64'h60a28d41_15029001,
        64'hfd1ff0ef_14020005,
        64'h041bfdbf_f0efe022,
        64'he4061141_80820141,
        64'h25016402_60a28d41,
        64'h0105151b_fe9ff0ef,
        64'h842afeff_f0efe022,
        64'he4061141_fc3ff06f,
        64'h96050513_00005517,
        64'h80822501_8d5d00f7,
        64'h17bb40f0_07bb00f7,
        64'h553b93ed_836d8f3d,
        64'h0127d713_e1189736,
        64'h00176713_02d786b3,
        64'h65186294_611c68e6,
        64'h86930000_46971220,
        64'h106f8082_61056902,
        64'h64a26442_60e28522,
        64'he99ff0ef_10f40023,
        64'h0247c783_85220ea4,
        64'h2e23681c_18f43423,
        64'h21478793_00001797,
        64'h18f43023_22478793,
        64'h00001797_16f43c23,
        64'h8fa78793_fffff797,
        64'he65ff0ef_04052823,
        64'h03253023_e90410f5,
        64'h02a34785_0ef52c23,
        64'h4799c57c_57fdcd21,
        64'h842a1660_10ef4505,
        64'h1c000593_84aa892e,
        64'hc7ad639c_c7bd651c,
        64'hcbad511c_cbbd4d5c,
        64'hcfad4401_4d1cc141,
        64'h4401e04a_e426ec06,
        64'he8221101_b7716000,
        64'h290010ef_71c50513,
        64'h00003517_01a98863,
        64'hd80fe0ef_856685e2,
        64'h00978e63_601cd8ef,
        64'he0ef855e_85ca0009,
        64'h0663d9af_e0ef638c,
        64'h855a0fc4_2603681c,
        64'h89560007_c3638952,
        64'h4c1cc791_4901541c,
        64'hdb8fe06f_61252d65,
        64'h05130000_45176d02,
        64'h6ca26c42_6be27b02,
        64'h7aa27a42_79e26906,
        64'h64a660e6_64460294,
        64'h15634d29_794c8c93,
        64'h00003c97_00050c1b,
        64'h218b8b93_00004b97,
        64'h218b0b13_00004b17,
        64'h218a8a93_00004a97,
        64'h218a0a13_00004a17,
        64'h89aae0ca_ec86e06a,
        64'he466e862_ec5ef05a,
        64'hf456f852_fc4e6080,
        64'he8a2aea4_84930000,
        64'h5497e4a6_711d8082,
        64'he308e518_e11ce788,
        64'h6798b027_87930000,
        64'h5797e508_80829407,
        64'hab230000_5797e79c,
        64'he39cb1a7_87930000,
        64'h5797b7d5_6000a8cf,
        64'hf0ef8522_c78119a4,
        64'h47838082_610564a2,
        64'h644260e2_00941763,
        64'h84beec06_e4266380,
        64'he822b4a7_87930000,
        64'h57971101_80824388,
        64'h9a078793_00005797,
        64'h80820f85_05138082,
        64'hc3980015_071b4388,
        64'h9b878793_00005797,
        64'hbfd55535_80826105,
        64'h64a26442_60e2e080,
        64'h0f840413_e501ce0f,
        64'hf0ef842a_cd09f7df,
        64'hf0ef84ae_e822ec06,
        64'he4261101_bfcdf840,
        64'h0513bfe5_45018082,
        64'h610560e2_5535e97f,
        64'he06f6105_60e200f7,
        64'h0c630ff0_07930815,
        64'h470302b7_006365a2,
        64'h10354703_c105fbdf,
        64'hf0efe42e_ec061101,
        64'h41488082_853ebfd1,
        64'h87b600a6_04630fc7,
        64'ha6038082_0141853e,
        64'h478160a2_f3cfe0ef,
        64'he4063325_05130000,
        64'h451785aa_114102e7,
        64'h90636394_631cc167,
        64'h07130000_57178082,
        64'h45018082_01414501,
        64'h640260a2_0dc000ef,
        64'h13e000ef_02c00513,
        64'hfc5ff0ef_85220005,
        64'h5563ac0f_e0ef8522,
        64'h12a000ef_c4f72423,
        64'h00005717_842ae406,
        64'he0224785_1141ef9d,
        64'h439cc5e7_87930000,
        64'h57978082_18b50d23,
        64'h8082557d_8082557d,
        64'h80824501_c56c8702,
        64'h972a4318_972a8379,
        64'hca050513_00003517,
        64'h1702ef05_6863450d,
        64'h0007081b_377d8b3d,
        64'h01a6571b_f0e51c63,
        64'h40000737_06bba423,
        64'h06dba223_06fba023,
        64'h04cbae23_018ba503,
        64'h45e646d6_47c64636,
        64'he8051763_842a90ff,
        64'he0efc4be_855e0107,
        64'h979b008c_460107cb,
        64'hd783c2be_479d04f1,
        64'h102347a5_06fb9e23,
        64'h04e15783_0007d663,
        64'h018ba783_ec051163,
        64'h842a943f_e0efc2be,
        64'h47d5855e_c4be0107,
        64'h979b008c_460107cb,
        64'hd78304f1_1023478d,
        64'h6ce000ef_06cb8513,
        64'h00ec4641_ef2ff06f,
        64'hfa100413_bf6d1187,
        64'h25839752_83790207,
        64'h9713fcfc_65e34581,
        64'hbfa1d171_d13fe0ef,
        64'h855e4585_0b700613,
        64'h0ff6f693_bb35f53d,
        64'h9d9fe0ef_855ec9af,
        64'hf0ef855e_460118fb,
        64'hae2308bb_a2230017,
        64'hb79317ed_088ba583,
        64'hef8d1afb_a823409c,
        64'he79d0046_f7930089,
        64'h2683f14d_feffe0ef,
        64'h855e408c_913fe0ef,
        64'h855e02eb_aa230017,
        64'hb71341b7_87b301a7,
        64'h86634711_00d78963,
        64'h47214000_06b70009,
        64'h2783bfa5_fb9910e3,
        64'h0931941f_e0ef855e,
        64'h035baa23_08fba223,
        64'h180bae23_1a0ba823,
        64'h088ba783_dabfe0ef,
        64'h855e4585_0b700613,
        64'h4681c90d_dbbfe0ef,
        64'h855e0fb6_f6934585,
        64'h0b700613_00894683,
        64'hc3a12781_8ff900f9,
        64'hf7b30009_270340dc,
        64'h04f71963_0017b793,
        64'h17ed0049_4703409c,
        64'h10000db7_20000d37,
        64'hf1090913_00003917,
        64'hbd2197bf_e0ef3fe5,
        64'h05130000_4517ff64,
        64'h98e304a1_eb992781,
        64'h00f9f7b3_00fa97bb,
        64'h409cf76c_8c930000,
        64'h3c974c2d_f44b0b13,
        64'h00003b17_4a85f2e4,
        64'h84930000_3497daaf,
        64'hf0ef2981_855e00f9,
        64'hf9b34601_088ba583,
        64'h044ba783_040ba983,
        64'he6f769e3_400407b7,
        64'h04fba023_00c7e793,
        64'h040ba783_d7dd8b85,
        64'h04dba023_0106e693,
        64'h040ba683_04dba023,
        64'h0216869b_c58900c7,
        64'hf593cd91_0027f593,
        64'h1abba423_03f7f593,
        64'h0c464783_04fba023,
        64'h0016879b_700006b7,
        64'hb1294c25_05130000,
        64'h4517e611_b5f1e225,
        64'hecf769e3_400407b7,
        64'h00f77863_1a0bb603,
        64'h400407b7_04fba023,
        64'h27851000_07b7b0cd,
        64'h02fba423_47857680,
        64'h10ef8526_a39fe0ef,
        64'h8a3d8abd_0146561b,
        64'h0106569b_06248513,
        64'h55058593_00004597,
        64'h074ba603_a59fe0ef,
        64'h04d48513_55458593,
        64'h00004597_0186d69b,
        64'h0ff77713_0ff7f793,
        64'h0ff6f813_0106d71b,
        64'h0086d79b_06cbc603,
        64'h077bc883_070ba683,
        64'ha8dfe0ef_fef53623,
        64'h02450513_57458593,
        64'h00004597_84aa06fb,
        64'hc603074b_d68307ab,
        64'hd70302c7_d7b3ed10,
        64'h92010a8b_b783d11c,
        64'h9fb90712_00e03733,
        64'h8f750207_161376c1,
        64'h9fb5068e_00d036b3,
        64'h8ef9f006_8693ff01,
        64'h06b79fb5_068a00d0,
        64'h36b38ef9_0f068693,
        64'hf0f0f6b7_9fb500f0,
        64'h37b30686_00d036b3,
        64'h27818ef9_8ff9ccc6,
        64'h8693aaa7_8793cccc,
        64'hd6b7aaaa_b7b708cb,
        64'ha7030005_06230005,
        64'h15234a00_00ef855e,
        64'h08fba823_08fba623,
        64'h20000793_c79919cb,
        64'ha7831afb_aa231b0b,
        64'ha7830adb_a2230afb,
        64'ha02302d6_06bb02f7,
        64'h57bb8a8d_0106d69b,
        64'h02e6073b_3e800613,
        64'hc30503f7_77130126,
        64'hd71bc78d_27818fd1,
        64'h8ff90186_d61b17fd,
        64'h67c100cd_a68308fb,
        64'hae230087_171b1487,
        64'ha78397b6_078a0966,
        64'h86930000_369704d6,
        64'h1c638003_06b7018b,
        64'ha60300f6_f8638bbd,
        64'h00c7579b_46a5008d,
        64'ha703fda5_9ee3fefd,
        64'h2e238fd9_8ff58f51,
        64'h0087d79b_8e690087,
        64'h961b8f51_0187971b,
        64'h0187d61b_0d11000d,
        64'h2783f006_869300ff,
        64'h0537040d_059366c1,
        64'hbf911187_25839752,
        64'h83790207_9713f6f7,
        64'h62e34581_472db575,
        64'hdef98be3_10bc0991,
        64'h81dff0ef_855e8405,
        64'h85934601_180bae23,
        64'h096ba223_1afba823,
        64'h017d85b7_4785f3f5,
        64'h37fd6702_67a2c521,
        64'hd51fe0ef_e03ac93a,
        64'he556e16a_e43e855e,
        64'h110c0110_04000713,
        64'h4791d502_8dead33a,
        64'h0af11023_fe0c7d13,
        64'h47b56702_ed05d7ff,
        64'he0efd53e_e03ad33a,
        64'h855e110c_0107979b,
        64'h46014755_07cbd783,
        64'h0af11023_03700793,
        64'h895ff0ef_855e4601,
        64'h18fbae23_08bba223,
        64'h0017b793_17ed088b,
        64'ha583efd9_1afba823,
        64'h409c09b7_90638bbd,
        64'h010cc783_e541dcff,
        64'he0efc93e_e556e166,
        64'h855e110c_04000793,
        64'h0110d53e_00fde7b3,
        64'h17c12d81_810007b7,
        64'hd33e47d5_0af11023,
        64'h47994d85_0ae79d63,
        64'h470d00e7_86634705,
        64'h409cd41f_e0ef855e,
        64'h02fbaa23_001d3793,
        64'h40fd0d33_100007b7,
        64'h00ed0863_47912000,
        64'h073700ed_0d6347a1,
        64'h40000737_0e051963,
        64'h8daa8bff_f0ef855e,
        64'h0015b593_40bd05b3,
        64'h100005b7_00fd0863,
        64'h45912000_07b700fd,
        64'h0d6345a1_400007b7,
        64'h12078e63_278101a7,
        64'hf7b300f9_77b30009,
        64'had0340dc_840b0b1b,
        64'h06010993_017d8b37,
        64'hbf0104fb_a0230087,
        64'he793040b_a783f207,
        64'h50e302e7_97138fd5,
        64'h8ff90087_d79b0087,
        64'h969bf007_07136741,
        64'h44dcfbe1_8b8583a5,
        64'h4cdce605_1de3eb7f,
        64'he0efdc3e_f84af426,
        64'hc556855e_010c0400,
        64'h07931030_c33e47d5,
        64'h08f11023_47990209,
        64'h886339fd_09053ac5,
        64'h49959881_19020100,
        64'h0ab70ff1_04934905,
        64'hbfa98003_0737b785,
        64'h80020737_00074563,
        64'h03079713_b7bda007,
        64'h071b8001_1737b949,
        64'hdf400413_e15fe0ef,
        64'h89850513_00005517,
        64'hfef493e3_3a478793,
        64'h00003797_04a1ebc5,
        64'h278100f9_77b300e7,
        64'h97bb4785_40980a85,
        64'h83f97913_02079a93,
        64'h478500f9_7933fe0c,
        64'h7c933c24_84930000,
        64'h3497044b_a783f0be,
        64'h0ff10c13_040ba903,
        64'h639c02a7_87930000,
        64'h579708f7_13638001,
        64'h07b7018b_a70304fb,
        64'ha0238fd9_20000737,
        64'h040ba783_00075963,
        64'h02d79713_00ebac23,
        64'h80010737_08d70e63,
        64'h4689c701_09270d63,
        64'h8b3d0187_d71b04eb,
        64'hac238f55_8f718ecd,
        64'h0087571b_8de90087,
        64'h159b8ecd_0187169b,
        64'h0187559b_40d804fb,
        64'haa232781_8fd58ef1,
        64'hf0070613_8fd16741,
        64'h0087569b_8e698fd5,
        64'h0087161b_0187179b,
        64'h0187569b_00ff0537,
        64'h4098bd79_8a9d9381,
        64'h00f6d69b_17828fd9,
        64'h01e6d71b_8ff90027,
        64'h979b1771_6705b545,
        64'h08bba823_00b515bb,
        64'h89bd0165_d59bbd91,
        64'h40040737_bda94003,
        64'h0737bd89_40020737,
        64'hbb75842a_fe0996e3,
        64'h39fdc529_844ff0ef,
        64'hd05aec56_e826855e,
        64'h108c0810_4b210a85,
        64'h4991d482_06f11023,
        64'h98810209_1a930330,
        64'h07930bf1_04934905,
        64'hd2caed05_874ff0ef,
        64'hd4bed2ca_855e0107,
        64'h979b108c_460107cb,
        64'hd78306f1_10230370,
        64'h079304fb_a0232789,
        64'h100007b7_54075963,
        64'h018ba703_e20515e3,
        64'h842aff3f_e0ef855e,
        64'h00b54583_113000ef,
        64'h855ee405_10e3842a,
        64'hc94ff0ef_855e08fb,
        64'h80a357fd_08fbaa23,
        64'h4785e405_1ce3842a,
        64'h8d8ff0ef_c4bec2ca,
        64'h855e008c_0107979b,
        64'h46014955_07cbd783,
        64'h04f11023_479d8f6f,
        64'hf0efc282_c4be04e1,
        64'h1023855e_008c4601,
        64'h0107979b_471100e7,
        64'h8e63577d_04cba783,
        64'hc21508fb_a82300e7,
        64'hf4632000_0793090b,
        64'ha70308fb_a6230107,
        64'hd4632000_07930afb,
        64'hb8230e0b_b0230c0b,
        64'hbc230c0b_b8230c0b,
        64'hb4230c0b_b0230a0b,
        64'hbc230307_87b300d7,
        64'h97b32689_078546a1,
        64'h8fd90106_d79b8f7d,
        64'h003f0737_0107979b,
        64'h14070f63_02cba703,
        64'h090ba823_1408dd63,
        64'h090ba623_00e5183b,
        64'h8b3d0107_d71b08eb,
        64'ha22308eb_a42304cb,
        64'ha823180b_ae231a0b,
        64'ha8238a05_00c7d61b,
        64'h02c7073b_018ba883,
        64'h45050f87_47031086,
        64'h26039652_9752060a,
        64'h8b3d5aaa_0a130000,
        64'h3a178a1d_0036571b,
        64'h00ebac23_4007071b,
        64'h40010737_a0292007,
        64'h071b4001_0737bf05,
        64'h06fb9e23_478502fb,
        64'ha6238b85_41e7d79b,
        64'h048ba783_00fbac23,
        64'h400007b7_bfe91bf0,
        64'h10ef0640_051308a9,
        64'h6fe31310_10ef8526,
        64'h0007cc63_048ba783,
        64'hf155842a_b1eff0ef,
        64'h855e4585_3e800913,
        64'h90810205_14931550,
        64'h10ef4501_afeff0ef,
        64'h855e0407_c163180b,
        64'h8c23048b_a7838082,
        64'h615d6db6_6d566cf6,
        64'h7c167bb6_7b567af6,
        64'h6a1a69ba_695a64fa,
        64'h741a70ba_8522d55d,
        64'h842ad99f_f0ef855e,
        64'ha031020b_a423f4fd,
        64'h34fd1005_0de3842a,
        64'ha88ff0ef_855e008c,
        64'h46014495_cf818b85,
        64'h1b8ba783_12050ae3,
        64'h842aaa2f_f0efc482,
        64'hc2be855e_008c479d,
        64'h460104f1_10234789,
        64'he7b5180b_8ca3198b,
        64'hc783c7b1_199bc783,
        64'h1e7010ef_45018baa,
        64'he3b54401_e6eeeaea,
        64'heee6f2e2_f6defada,
        64'hfed6e352_e74eeb4a,
        64'hef26f706_f3227161,
        64'h551cb585_84aab595,
        64'hfa100493_9fcff0ef,
        64'hc5050513_00005517,
        64'hd965c04f_f0ef8522,
        64'h4585bfd1_18f40c23,
        64'h47850007_d663443c,
        64'hed09c1cf_f0ef8522,
        64'h4581becf_f0ef8522,
        64'h02f51f63_f9200793,
        64'hb55d18f4_0ca34785,
        64'h06041e23_d45c8b85,
        64'h41e7d79b_c43ccc18,
        64'h80010737_00e68563,
        64'h80020737_4c14bf45,
        64'h319010ef_3e800513,
        64'h06090863_397d0007,
        64'hca6347b2_ed1db76f,
        64'hf0ef8522_858a4601,
        64'hc43e0197_e7b30187,
        64'h1563c43e_0177f7b3,
        64'hc25a4bdc_01511023,
        64'h4c18681c_e13db9ef,
        64'hf0efc402_c2520131,
        64'h10238522_858a4601,
        64'h40000cb7_80020c37,
        64'h00ff8bb7_4b050290,
        64'h0a934a55_03700993,
        64'h3e900913_cc1c8002,
        64'h07b700f7_15630aa0,
        64'h079300c1_4703e911,
        64'hbe0ff0ef_c23ec43a,
        64'h8522858a_460147d5,
        64'h0aa00713_e3991aa0,
        64'h07138ff9_4bdc00ff,
        64'h8737681c_00f11023,
        64'h47a10005_05a346d0,
        64'h00ef8522_f14984aa,
        64'hcdaff0ef_8522f13f,
        64'hf0ef8522_45814601,
        64'hb5eff0ef_8522d85c,
        64'h478508f4_22231a04,
        64'h28231804_2e230884,
        64'h2783f945_84aa9782,
        64'h6b9c679c_8522681c,
        64'h409010ef_7d000513,
        64'hb8eff0ef_85220204,
        64'h2c2302f4_08234785,
        64'h1af42c23_478df93f,
        64'hf0eff3e5_4481541c,
        64'h80826109_7ca27c42,
        64'h7be26b06_6aa66a46,
        64'h69e674a6_79068526,
        64'h744670e6_f8500493,
        64'hb98ff0ef_dd450513,
        64'h00005517_02042423,
        64'heb8d6b9c_679c681c,
        64'hc509f07f_f0ef842a,
        64'hc17c8fd9_f466f862,
        64'hfc5ee0da_e4d6e8d2,
        64'heccef0ca_f4a6fc86,
        64'hf8a2070d_4b9c7119,
        64'h10000737_691c8082,
        64'h8082c18f_f06f02c5,
        64'h0823dd0c_0007859b,
        64'h87ba00d5_f3630007,
        64'h069b0007_859b4f18,
        64'h87ae00d5_f3630007,
        64'h869b4f5c_6918e215,
        64'hb7cdc402_fef414e3,
        64'h47858082_61217902,
        64'h74a27442_70e2d26f,
        64'hf0ef8526_858a4601,
        64'hc43e4789_00f41f63,
        64'h4791c24a_00f11023,
        64'h4799ed19_d44ff0ef,
        64'hc43ec24a_8526858a,
        64'h46010107_979b4955,
        64'h842e07c4_d78300f1,
        64'h10230370_079304f5,
        64'h92635529_478500f5,
        64'h866384aa_4791f04a,
        64'hf822fc06_f4267139,
        64'h80820141_640260a2,
        64'h45058302_014160a2,
        64'h64028522_00030763,
        64'h0187b303_679c681c,
        64'h00055e63_ffdfe0ef,
        64'h842ae406_e0221141,
        64'hb325842a_b335dd79,
        64'h842a941f_f0ef8526,
        64'h45850a70_061386ca,
        64'hb381842a_953ff0ef,
        64'h85264585_09b00613,
        64'h46850127_9b630a79,
        64'hc783d4fb_0ee34785,
        64'hed19971f_f0ef8526,
        64'h458509c0_061386de,
        64'hfdba18e3_0c110ffa,
        64'h7a132a0d_ffac90e3,
        64'h0ffafa93_2ca12a85,
        64'he139999f_f0ef8526,
        64'h0ff6f693_0196d6bb,
        64'h45858656_000c2683,
        64'h4c818ad2_09b00d93,
        64'h4d6108f0_0a13ff9a,
        64'h10e32a05_e92d9c5f,
        64'hf0ef8526_45850ff6,
        64'h76130ff6_f693f8ca,
        64'h061b00da_d6bb003a,
        64'h169b4c8d_fdbd1fe3,
        64'h2d05e945_8a2a9edf,
        64'hf0ef8526_45850ff6,
        64'h76130ff6_f693f88d,
        64'h061b00dc_d6bb003d,
        64'h169b4d91_4d0108f4,
        64'haa2300a7_979b0e09,
        64'hc7830af9_87a34785,
        64'he579a21f_f0ef8526,
        64'h45850af0_06134685,
        64'he3958b85_0af9c783,
        64'he20b05e3_b535547d,
        64'hdb8ff0ef_fd450513,
        64'h00005517_cb898b85,
        64'h09b9c783_bfd100f9,
        64'h7933fff7_c793b5a9,
        64'h2f8020ef_fa450513,
        64'h00005517_ef898b85,
        64'h0a69c783_02d90263,
        64'hfcb614e3_87b20ff9,
        64'h79130127_e933c70d,
        64'h4189591b_4187d79b,
        64'h8b050189_191b0187,
        64'h979b0027_571b00c5,
        64'h17bbc39d_8b850017,
        64'h579b4b98_97d2078e,
        64'h0017861b_45914505,
        64'h47810016_e913c399,
        64'h0fe6f913_8b89c719,
        64'h89360017_f7130a79,
        64'hc683008a_4783b5c9,
        64'he50ff0ef_fec50513,
        64'h00005517_85ca0126,
        64'h7a63963e_09d9c783,
        64'h9e3d0087_979b0106,
        64'h161b09e9_c78309f9,
        64'hc603ee05_1ae3842a,
        64'hf8aff0ef_852685ce,
        64'hee068de3_ff450513,
        64'h00005517_8a89000b,
        64'h8963fa65_96e387ae,
        64'h06110521_0128893b,
        64'h0ffbfb93_00fbebb3,
        64'h00be17bb_cb898b85,
        64'h0107c783_97d2078e,
        64'h02080063_01162023,
        64'h02e858bb_b7f14b81,
        64'h4a814c81_b7c9ed6f,
        64'hf0ef0125_05130000,
        64'h55170008_8d6302e8,
        64'h78bb0017_859b0005,
        64'h28034311_4e054781,
        64'h89568662_00ca0513,
        64'h8c0a009c_9c9be399,
        64'h4b8502ea_dabb54dc,
        64'hb7615429_f14ff0ef,
        64'h01850513_00005517,
        64'hcb8902ec_f7bb0005,
        64'hac83e791_02eaf7bb,
        64'h060a8063_fe09f993,
        64'h02f10993_0045aa83,
        64'hdb4501a5_05130000,
        64'h55170984_a7038082,
        64'h2a010113_23813d83,
        64'h24013d03_24813c83,
        64'h25013c03_25813b83,
        64'h26013b03_26813a83,
        64'h27013a03_27813983,
        64'h28013903_28813483,
        64'h29013403_29813083,
        64'h8522f840_0413f8ef,
        64'hf0ef0425_05130000,
        64'h5517e7b9_0016f793,
        64'h07e4c683_00e7eb63,
        64'h02050513_00005517,
        64'h8a2e8b32_84aabfe7,
        64'h87933ffc_07b79f3d,
        64'hbff7879b_bffc07b7,
        64'h4d180ac7_ed634789,
        64'h23b13c23_25a13023,
        64'h25913423_25813823,
        64'h25713c23_27613023,
        64'h27513423_27413823,
        64'h27313c23_29213023,
        64'h28913423_28813823,
        64'h28113c23_d6010113,
        64'h80826145_69a26942,
        64'h64e27402_70a28522,
        64'h013505a3_17a010ef,
        64'h8526842a_86dff0ef,
        64'h852685ca_00091c63,
        64'h00f51e63_842a57b5,
        64'hc519cc1f_f0ef84aa,
        64'h45850b30_06138edd,
        64'h892e9be1_0079f693,
        64'h0ff5f993_08154783,
        64'hf022f406_e44ee84a,
        64'hec267179_bfd984aa,
        64'hb7554685_fef760e3,
        64'h54a94705_ffc5879b,
        64'h80822401_01132281,
        64'h34832201_39038526,
        64'h23013403_23813083,
        64'hdf400493_e3990b94,
        64'h4783e915_9a7ff0ef,
        64'h854a85a2_980101f1,
        64'h0413ed91_258199f5,
        64'hffe4059b_e11d84aa,
        64'hd3fff0ef_892a4585,
        64'h0b900613_842eed85,
        64'h54a94681_04b7ec63,
        64'h06f58463_47892321,
        64'h30232291_34232281,
        64'h38232211_3c23dc01,
        64'h0113b765_5929b775,
        64'h5951bf45_1a04b023,
        64'h54c020ef_dd4d1a04,
        64'hb503892a_b75d08f4,
        64'haa2302f7_07bb2785,
        64'h27058bfd_8b7d0057,
        64'hd79b00a7_d71b50fc,
        64'hf3dd8b85_0af44783,
        64'h80822501_01132281,
        64'h39832301_39032381,
        64'h3483854a_24013403,
        64'h24813083_08f48023,
        64'h0a744783_08f4ac23,
        64'h00a7979b_02e787bb,
        64'h0dd44703_0e044783,
        64'hf8dc07a6_0d442783,
        64'h00098663_c79954dc,
        64'h08f4aa23_00a7979b,
        64'h0e044783_0af407a3,
        64'h4785e141_e0bff0ef,
        64'h85264585_0af00613,
        64'h4685c6b5_e3918bfd,
        64'h09c44783_c7898b85,
        64'h0a044783_f4fc07a6,
        64'hc319f4fc_54d89fb9,
        64'h08844703_9fb90087,
        64'h171b0894_47039fb9,
        64'h0107171b_0187979b,
        64'h08a44703_08b44783,
        64'hf8fc07ce_02e787b3,
        64'h0dd44783_02f70733,
        64'h0e044703_97ba08c4,
        64'h47039fb9_0087171b,
        64'h0107979b_468508d4,
        64'h470308e4_47830409,
        64'h8f63fce5_14e30621,
        64'h070de21c_07ce02b7,
        64'h87b30dd4_478302f5,
        64'h85b30e04_45830009,
        64'h8c634685_c39197ae,
        64'hffe74583_9fad0105,
        64'h959b0087_979b0007,
        64'h4583fff7_4783e0fc,
        64'h07c64681_09d40513,
        64'h0a844783_fcdc07c6,
        64'h0c848613_09140713,
        64'h0e244783_06f48fa3,
        64'h09c44783_c7898b89,
        64'h0a044783_00098a63,
        64'h08f480a3_0b344783,
        64'hc7890e24_4783e781,
        64'h0019f993_8b8506f4,
        64'h8f2309b4_49830a04,
        64'h4783f8dc_00d77363,
        64'h0147d693_07a68007,
        64'h07136705_0d442783,
        64'h00e7fd63_cc981ff7,
        64'h87934004_07b753b8,
        64'h97ba078a_fa470713,
        64'h00004717_1cf76d63,
        64'h47210c04_478313d0,
        64'h10ef85a2_20000613,
        64'h1e050563_1a04b503,
        64'h1aa4b023_6ee020ef,
        64'h20000513_e7991a04,
        64'hb7831e05_1a63892a,
        64'hc03ff0ef_84aa85a2,
        64'h980101f1_04131ce7,
        64'hf3634901_3ffc0737,
        64'h23313423_22913c23,
        64'h24813023_24113423,
        64'h9fb92321_3823bffc,
        64'h07b7db01_01134d18,
        64'hbfcdfc79_347d8082,
        64'h612174a2_744270e2,
        64'hd8bff0ef_85263e80,
        64'h0593e919_c4dff0ef,
        64'h8526858a_4601440d,
        64'hc432c23e_84aafc06,
        64'hf426f822_47f58e55,
        64'h00f11023_030006b7,
        64'h8e554799_71390106,
        64'h161b0086_969b8082,
        64'h61216aa2_6a4269e2,
        64'h74a27902_85267442,
        64'h70e2fc09_99e39aa2,
        64'h02878433_9a224089,
        64'h89b308c9_6783fc85,
        64'h1ae3f01f_f0ef854a,
        64'h85d68652_86a2844e,
        64'h0089f363_0207e403,
        64'h01093783_89a6f96d,
        64'hecdff0ef_854a08c9,
        64'h2583a089_4481bd7f,
        64'hf0ef4225_05130000,
        64'h551700b6_7a630144,
        64'h85b36810_00054d63,
        64'h869fa0ef_852200b4,
        64'h4583c11d_892a4a40,
        64'h10ef8ab6_84b28a2e,
        64'h4148842a_ce05e456,
        64'he852ec4e_f04af426,
        64'hf822fc06_7139b7c5,
        64'h4401b7d5_0004841b,
        64'hb74d02f6_063bbf61,
        64'h47c58082_61256906,
        64'h64a66446_60e68522,
        64'hc41ff0ef_46c50513,
        64'h00005517_c11dd4ff,
        64'hf0efd23e_d402854a,
        64'h100c47f5_460102f1,
        64'h102347b1_0497f063,
        64'h4785e529_842ad6ff,
        64'hf0efc83e_ca26d23a,
        64'h854a100c_47850030,
        64'hcc3ee42e_4755d432,
        64'hcf3108c9_27832601,
        64'h02f11023_02c92703,
        64'h47c906d7_f66384b6,
        64'h892a4785_e8a2ec86,
        64'he0cae4a6_711d8082,
        64'h4501bfd5_45018082,
        64'h612174a2_744270e2,
        64'hf8ed34fd_c901dc7f,
        64'hf0ef8522_858a4601,
        64'h4495cb91_8b891b84,
        64'h2783c11d_dddff0ef,
        64'hc23e842a_f426fc06,
        64'hf822858a_460147d5,
        64'hc42e00f1_102347c1,
        64'h7139e7a9_19c52783,
        64'hbf6df920_0513d07f,
        64'hf0ef5125_05130000,
        64'h5517fc80_47e34501,
        64'h8456b74d_84565d60,
        64'h20ef3e80_05130080,
        64'h5863fff4_0a9bfe04,
        64'hc5e334fd_80826125,
        64'h7b027aa2_7a4279e2,
        64'h690664a6_644660e6,
        64'hfba00513_d4dff0ef,
        64'h54050513_00005517,
        64'hc7950125_f7b30547,
        64'h95630135_f7b3c789,
        64'h1005f793_45b2ed15,
        64'he71ff0ef_855a858a,
        64'h4601e00a_0a13e009,
        64'h89930809_09134495,
        64'hc43e842e_8b2af456,
        64'hec86f05a_e4a6e8a2,
        64'h6a056989_fdf94937,
        64'h0107979b_f852fc4e,
        64'he0ca07c5_5783c23e,
        64'h47d500f1_102347b5,
        64'h711d8082_61457402,
        64'h70a2c43c_47b2e119,
        64'hec9ff0ef_8522858a,
        64'h4601c43e_8fd94000,
        64'h07378fd9_8f756000,
        64'h06b78ff5_8ff9f806,
        64'h86934bdc_008006b7,
        64'h4538691c_c195842a,
        64'hc402c23e_f406f022,
        64'h478500f1_10234785,
        64'h71798082_61457402,
        64'h70a28522_6cc020ef,
        64'h7d000513_e509842a,
        64'hf21ff0ef_c202c402,
        64'h00011023_858a4601,
        64'h85226ea0_20eff406,
        64'h3e800513_842af022,
        64'h71798082_4501bf65,
        64'h4501fd45_59b010ef,
        64'h0d448513_0d440593,
        64'h4611fcf7_15e30e04,
        64'h47830e04_c703fcf7,
        64'h1be30c04_47830c04,
        64'hc703fef7_11e30dd4,
        64'h47830dd4_c7038082,
        64'h24010113_22813483,
        64'h23013403_23813083,
        64'hfb600513_00f70d63,
        64'h0a044783_0a04c703,
        64'he909fadf_f0ef1a05,
        64'h34832211_3c232291,
        64'h342385a2_980101f1,
        64'h04132281_3823dc01,
        64'h011308e6_e0634004,
        64'h07374d14_80826161,
        64'h60a6fd3f_f0efcc3e,
        64'hd402e486_100c2000,
        64'h07930030_e83ee42e,
        64'h07851782_4785d23e,
        64'h47d502f1_102347a1,
        64'h715d8302_0007b303,
        64'h679c691c_80826e65,
        64'h05130000_55178082,
        64'h6108953e_81753fe7,
        64'h87930000_47971502,
        64'h00a7eb63_47ad8082,
        64'h557d8082_01416402,
        64'h60a24501_83020141,
        64'h60a26402_85220003,
        64'h07630207_b303679c,
        64'h681c0005_5e63ff5f,
        64'hf0ef842a_e406e022,
        64'h11418082_557d8082,
        64'h557db7f1_659c95aa,
        64'h058e05e1_35f1bfe1,
        64'h617cbff1_7d5c8082,
        64'h61054501_6442e900,
        64'h64a260e2_02945433,
        64'h0e7010ef_90811482,
        64'h7540f55c_08c52483,
        64'h795c8782_97b6e426,
        64'he822ec06_1101431c,
        64'h97360025_97134666,
        64'h86930000_469704b7,
        64'hec63479d_80824501,
        64'h83020003_03630087,
        64'hb303679c_691c8082,
        64'h61356452_60f28522,
        64'h125020ef_0808842a,
        64'he3fff0ef_e436eec6,
        64'heac2e6be_e2baea22,
        64'hee060808_10000593,
        64'h1234862a_fe36fa32,
        64'hf62e710d_80826161,
        64'h60e2e69f_f0efe436,
        64'he4c6e0c2_fc3ef83a,
        64'hec061000_05931014,
        64'h862ef436_f032715d,
        64'h80826161_60e2e8df,
        64'hf0efe436_e4c6e0c2,
        64'hfc3ef83a_ec061034,
        64'hf436715d_b7f18522,
        64'h02010393_0005059b,
        64'h501010ef_85220124,
        64'h74336000_00840b13,
        64'hb5fd845a_d89ff0ef,
        64'h00840b13_02010393,
        64'h00044503_a809dd1f,
        64'hf0ef0028_02010393,
        64'h0005059b_e31ff0ef,
        64'h400845a9_46010016,
        64'hb6930038_00840b13,
        64'hf8b50693_a81145c1,
        64'h00163613_46850038,
        64'h00840b13_fa850613,
        64'hf6e510e3_07800713,
        64'h02e50063_07500713,
        64'ha00d4601_46850038,
        64'h00840b13_f6e51ee3,
        64'h07000713_00a76c63,
        64'h06e50e63_07300713,
        64'hb74d048d_0024c503,
        64'h80826109_0007051b,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_744670e6,
        64'hf55d08f5_09630630,
        64'h079304d5_0f630580,
        64'h069302a6_eb6306d5,
        64'h0f630640_06930489,
        64'h0014c503_478100f6,
        64'hf36346a5_0ff7f793,
        64'hfd07879b_cb9d0004,
        64'hc7830355_10634781,
        64'h04890545_0f630014,
        64'hc503bfe1_e71ff0ef,
        64'h02010393_04850135,
        64'h086304d7_ff639381,
        64'h17827682_0017079b,
        64'hc52d8f1d_0004c503,
        64'h77a27742_02095913,
        64'h03000a93_06c00a13,
        64'h02500993_f82af02e,
        64'hf42afc3e_843684b2,
        64'he0dafc86_e4d6e8d2,
        64'heccef4a6_f8a2597d,
        64'h011cf0ca_7119b7e1,
        64'h01178023_00660023,
        64'h06850006_48830007,
        64'hc30300d7_063397ba,
        64'h93811782_40f807bb,
        64'hb7d1feb5_0fa30505,
        64'hbf4500c8_063b8082,
        64'h00b7ea63_0006879b,
        64'hfff5081b_46810015,
        64'h559b9d19_00050023,
        64'h050500f5_002302d0,
        64'h07930003_076302f6,
        64'he96300a6_06bb0300,
        64'h059340e0_063b8536,
        64'hfcb8ffe3_02b8d53b,
        64'hfec68fa3_06850ff6,
        64'h76130306_061b04ae,
        64'h6a630ff5_761302b8,
        64'hf53b0005_089b3859,
        64'h86ba4e25_0ff6f813,
        64'h04100693_c2190610,
        64'h06934305_40a0053b,
        64'he6810005_56634301,
        64'hbfd900d7_00230785,
        64'h0006c683_00f506b3,
        64'h00d3b823_00170693,
        64'h8082852e_00070023,
        64'h00b6e663_0103b703,
        64'h0007869b_47819d9d,
        64'hfff7059b_00c6f563,
        64'h8e9dfff7_06930003,
        64'hb7038f99_92010205,
        64'h96130103_b7830083,
        64'hb7038082_45018082,
        64'h00078023_45050103,
        64'hb78300a7_002300f3,
        64'hb8230017_079300d7,
        64'hfe639381_17822785,
        64'h40f707b3_0003b683,
        64'h0083b783_0103b703,
        64'h80826145_45016a02,
        64'h69a26942_64e27402,
        64'h70a22f20_00ef00e5,
        64'h05130000_6517fd24,
        64'h1de33020_00ef8191,
        64'h00f5f613_0405854e,
        64'h0007c583_008487b3,
        64'h318000ef_8552e781,
        64'h0004059b_01f47793,
        64'h20000913_af498993,
        64'h00006997_af4a0a13,
        64'h00006a17_4401ed9f,
        64'hf0ef8526_45813460,
        64'h00efaf25_05130000,
        64'h6517dca6_06130000,
        64'h6617e789_a6c60613,
        64'h00006617_584c19c4,
        64'h2783d65f_b0ef0865,
        64'h85930000_65977448,
        64'h098030ef_b1450513,
        64'h00006517_384000ef,
        64'hb0850513_00006517,
        64'ha9058593_00006597,
        64'hc789aa25_85930000,
        64'h6597545c_3a4000ef,
        64'hb1850513_00006517,
        64'h5c0c3b20_00ef0186,
        64'h561b0ff6_f6930ff7,
        64'h77130ff6_77930106,
        64'h569b0086_571bb265,
        64'h05130000_651706c4,
        64'h45835830_3dc000ef,
        64'h91c115c2_0085d59b,
        64'hb3050513_00006517,
        64'h546c3f20_00efb265,
        64'h05130000_651706f4,
        64'h45834020_00ef638c,
        64'hb2850513_00006517,
        64'h681c2240_10ef842a,
        64'h4bf010ef_45014790,
        64'h10ef0001_b5031460,
        64'h30efb425_05130000,
        64'h651784aa_03e030ef,
        64'he052e44e_e84aec26,
        64'hf022f406_20000513,
        64'h71797a00_006f6105,
        64'h468560e2_66226442,
        64'h85a25010_10efe42e,
        64'hec064501_842ae822,
        64'h11018082_01416402,
        64'h60a2557d_e3914505,
        64'h703c1040_30efade5,
        64'h05130000_6517ace5,
        64'h85930000_659734c0,
        64'h06139126_86930000,
        64'h569702f4_02632000,
        64'h07b7e406_6380e022,
        64'h1141711c_80822501,
        64'h638897aa_200007b7,
        64'h050ef73f_f06f2000,
        64'h05374581_46098082,
        64'hb7f9c45c_4785d8f1,
        64'h45018885_bfe94501,
        64'hc45c4789_c7890024,
        64'hf793f404_01242423,
        64'he01c2000_07b78082,
        64'h614569a2_694264e2,
        64'h740270a2_557d1520,
        64'h30ef8522_00099d63,
        64'h508000ef_bec50513,
        64'h00006517_862285aa,
        64'h89aa7b30_10ef9765,
        64'h05130000_551785a2,
        64'hc41d5551_842a1380,
        64'h30ef892e_84b2e44e,
        64'hf406e84a_ec26f022,
        64'h04800513_717908b0,
        64'h41635535_b7dd87ca,
        64'h14e109a1_3c2020ef,
        64'he43e002c_4621854e,
        64'h639c0087_8913dcd5,
        64'h01096483_00093983,
        64'h97a667a1_bf41b1bf,
        64'hf0ef8522_b77100f9,
        64'h26230009_b783dbd9,
        64'h8b85bd85_645020ef,
        64'h4505d809_8ce3c43f,
        64'hf0ef8522_484cc85c,
        64'h9bf54985_485cb4bf,
        64'hf0ef8522_ef8d8b85,
        64'h00892783_00090963,
        64'h04043023_246030ef,
        64'h855a85d6_0ca00613,
        64'ha0868693_00005697,
        64'h01848c63_04043903,
        64'h6004cc9d_49858889,
        64'hc85c9bf9_485cc85c,
        64'h0027e793_485ccbb5,
        64'h603cfeb6_90e30791,
        64'h872a2685_c3988f51,
        64'h8361ff87_37030106,
        64'h8763c390_0086161b,
        64'hff870513_63104591,
        64'h480d4681_00c90793,
        64'h01898713_08e69f63,
        64'h0037f693_470d0204,
        64'h3c230049_2783cba9,
        64'h7c1c2c40_30ef855a,
        64'h85d609c0_0613a6e6,
        64'h86930000_56970189,
        64'h8c630384_39030004,
        64'h3983cfb5_0014f793,
        64'h660000ef_d1c50513,
        64'h00006517_85cad1bf,
        64'hf0ef85ca_29010049,
        64'h6913ff39_79138522,
        64'h01442903_c39d0084,
        64'hf79368a0_00efd1e5,
        64'h05130000_651785ca,
        64'hd45ff0ef_85ca2901,
        64'h00896913_ff397913,
        64'h85220144_2903c39d,
        64'h0044f793_b29ff0ef,
        64'h85224581_b71ff0ef,
        64'h85224581_cc5cf920,
        64'h0793c781_7c1c00f7,
        64'h6f630c89_37830209,
        64'h37031404_80632481,
        64'h8cfd4981_485c0709,
        64'h34833740_30ef855a,
        64'h85d60f20_061386e6,
        64'h01890963_00043903,
        64'hb7117020_00efd7e5,
        64'h05130000_6517b065,
        64'h85930000_5597000b,
        64'h9d633bfd_20000c37,
        64'h8bd2bd61_00c4e493,
        64'hbd853b40_30efd8e5,
        64'h05130000_6517d7e5,
        64'h85930000_65971490,
        64'h0613b226_86930000,
        64'h5697b765_47014781,
        64'h2585e31c_97469381,
        64'h83751782_170200be,
        64'h873b8fd9_8fe90107,
        64'h67330087_d79b01c8,
        64'h78330087_981b0107,
        64'h67330187_971b0187,
        64'hd81bf2e5_00670363,
        64'h16fd0605_27810107,
        64'he7b301e8_183b0705,
        64'h00371f1b_00064803,
        64'hec0689e3_6e89f005,
        64'h051300ff_0e374311,
        64'h47014781_45816390,
        64'h0107e683_65410004,
        64'h3883603c_ee079be3,
        64'h8b85449c_df5ff0ef,
        64'h8522488c_db9ff0ef,
        64'he0248522_44cc8082,
        64'h61654501_6ce27c02,
        64'h7ba27b42_7ae26a06,
        64'h69a66946_64e67406,
        64'h70a6efe9_485ce5eb,
        64'h0b130000_6b17e4ea,
        64'h8a930000_6a97ebbf,
        64'hf0ef2581_0015e593,
        64'hc30c8c93_00005c97,
        64'h85220d89_b583cdbf,
        64'hf0ef8522_4585e9bf,
        64'hf0ef8522_24058593,
        64'h000f45b7_d31ff0ef,
        64'h85224581_46054685,
        64'h4705cfff_f0ef8522,
        64'h4581cc7f_f0ef8522,
        64'h85a6c8bf_f0ef681a,
        64'h0a138522_00095583,
        64'hc55ff0ef_00989a37,
        64'h85220089_2583be3f,
        64'hf0ef8522_4581d73f,
        64'hf0ef8522_45814605,
        64'h46814705_0144e493,
        64'h16078663_8b85008a,
        64'h2783000a_09638cdd,
        64'h03243c23_4c1c4485,
        64'he391448d_8b89c709,
        64'h0017f713_44810049,
        64'h278316f9_9a630404,
        64'h3a032000_07b70004,
        64'h3983bf7f_f0ef4585,
        64'h60080e04_9c636f60,
        64'h20ef00c9_05134581,
        64'h4611d01c_e03084b2,
        64'h892e0005_d7830204,
        64'h08a3ec66_f062f45e,
        64'hf85afc56_e0d2e4ce,
        64'hf486e8ca_eca67100,
        64'hf0a27159_80826105,
        64'h690264a2_644260e2,
        64'hc8440499_3c235a80,
        64'h30eff825_05130000,
        64'h6517f725_85930000,
        64'h65970760_0613d066,
        64'h86930000_569702f9,
        64'h026384ae_842a2000,
        64'h07b7ec06_e426e822,
        64'h00053903_e04a1101,
        64'h80826105_64a26442,
        64'h60e2e424_5ee030ef,
        64'hfc850513_00006517,
        64'hfb858593_00006597,
        64'h06f00613_d3c68693,
        64'h00005697_02f40263,
        64'h84ae2000_07b7ec06,
        64'he4266100_e8221101,
        64'h80826105_64a26442,
        64'h60e2e0a0_90511452,
        64'h632030ef_00c50513,
        64'h00006517_ffc58593,
        64'h00006597_06800613,
        64'hd7068693_00005697,
        64'h02f48263_842e2000,
        64'h07b7ec06_e8226104,
        64'he4261101_80826105,
        64'h64a26442_60e2fc80,
        64'h90411442_676030ef,
        64'h05050513_00006517,
        64'h04058593_00006597,
        64'h06100613_da468693,
        64'h00005697_02f48263,
        64'h842e2000_07b7ec06,
        64'he8226104_e4261101,
        64'hd4dff06f_01414581,
        64'h60a26402_6008f23f,
        64'hf0ef4605_46854705,
        64'h45818522_ef1ff0ef,
        64'h45818522_f39ff0ef,
        64'h842a4581_04053023,
        64'h02053c23_46054681,
        64'h4705e022_e4061141,
        64'h80820141_45016402,
        64'h60a2d97f_f0ef4581,
        64'h6008f67f_f0ef4581,
        64'h46054685_47058522,
        64'hf35ff0ef_45818522,
        64'hf7dff0ef_e4064581,
        64'h85224605_46814705,
        64'h7100e022_11418082,
        64'h612169e2_790274a2,
        64'h744270e2_0289b823,
        64'h8c4588a1_01246433,
        64'h0034949b_8c590049,
        64'h79130029_191b8b05,
        64'h88090014_141b6722,
        64'h75a030ef_e43a1365,
        64'h05130000_65171265,
        64'h85930000_659705a0,
        64'h0613e7a6_86930000,
        64'h569702f9_84638436,
        64'h893284ae_200007b7,
        64'hfc06f04a_f426f822,
        64'h00053983_ec4e7139,
        64'h80826105_64a26442,
        64'h60e2f404_7a6030ef,
        64'h18050513_00006517,
        64'h17058593_00006597,
        64'h05300613_eb468693,
        64'h00005697_02f40263,
        64'h84ae2000_07b7ec06,
        64'he4266100_e8221101,
        64'h80826105_64a26442,
        64'h60e2f004_7e6030ef,
        64'h1c050513_00006517,
        64'h1b058593_00006597,
        64'h04c00613_ee468693,
        64'h00005697_02f40263,
        64'h84ae2000_07b7ec06,
        64'he4266100_e8221101,
        64'h80826105_64a26442,
        64'h60e2ec80_90011402,
        64'h02b030ef_20450513,
        64'h00006517_1f458593,
        64'h00006597_04500613,
        64'hdd068693_00007697,
        64'h02f48263_842e2000,
        64'h07b7ec06_e8226104,
        64'he4261101_80826105,
        64'h64a26442_60e2e880,
        64'h90011402_06f030ef,
        64'h24850513_00006517,
        64'h23858593_00006597,
        64'h03e00613_e1c68693,
        64'h00007697_02f48263,
        64'h842e2000_07b7ec06,
        64'he8226104_e4261101,
        64'h80826105_64a26442,
        64'h60e2e404_0af030ef,
        64'h28850513_00006517,
        64'h27858593_00006597,
        64'h03600613_f9c68693,
        64'h00005697_02f40263,
        64'h84ae2000_07b7ec06,
        64'he4266100_e8221101,
        64'h80826105_64a26442,
        64'h60e2e004_0ef030ef,
        64'h2c850513_00006517,
        64'h2b858593_00006597,
        64'h02f00613_fcc68693,
        64'h00005697_02f40263,
        64'h84ae2000_07b7ec06,
        64'he4266100_e8221101,
        64'h80826105_64a26442,
        64'h60e2fc24_12f030ef,
        64'h30850513_00006517,
        64'h2f858593_00006597,
        64'h08800613_ff468693,
        64'h00005697_02f50263,
        64'h84ae842a_200007b7,
        64'hec06e426_e8221101,
        64'h8082556d_bfe50007,
        64'hac238082_4501cf98,
        64'h02000713_00d71763,
        64'h469100d7_0d63711c,
        64'h46a15958_80826149,
        64'h640a60aa_f83ff0ef,
        64'h0808f01f_f0ef0808,
        64'he85ff0ef_080885a2,
        64'h6622f71f_f0efe42e,
        64'he5060808_842ae122,
        64'h71758082_61051c65,
        64'h05130000_751760e2,
        64'hfca71de3_fef68fa3,
        64'hfec68f23_0007c783,
        64'h97ae0006_46038bbd,
        64'h962e0047_d6130705,
        64'h06890007_c78300e1,
        64'h07b34541_39458593,
        64'h00006597_20468693,
        64'h00007697_47013e50,
        64'h20efec06_850a4641,
        64'h05050593_11018082,
        64'he13cb807_87930000,
        64'h0797ed3c_639cf4e7,
        64'h87930000_7797e93c,
        64'h04053423_639cf567,
        64'h87930000_77978082,
        64'h614569a2_694264e2,
        64'h740270a2_fd24fde3,
        64'h45019782_8522603c,
        64'hfc1c078e_643c0124,
        64'hf5633f30_20ef9522,
        64'h45819201_16020006,
        64'h091b40a9_863b449d,
        64'h04000993_00e78023,
        64'h97a2f800_07130017,
        64'h8513e84a_f406e44e,
        64'hec26842a_03f7f793,
        64'hf0227179_653c8082,
        64'h61616ba2_6b426ae2,
        64'h7a0279a2_794274e2,
        64'h640660a6_b7c99782,
        64'h44018526_60bc0174,
        64'h176399d6_41590933,
        64'h4a7020ef_0144043b,
        64'h86560084_853385ce,
        64'h020ada93_020a1a93,
        64'h00090a1b_00f97463,
        64'h93811782_00078a1b,
        64'h408b07bb_04000b93,
        64'h04000b13_e53c8932,
        64'h89ae84aa_97b203f7,
        64'hf413ec56_f052e486,
        64'he45ee85a_f44ef84a,
        64'hfc26e0a2_715d653c,
        64'h80826105_692264c2,
        64'hcd70cd34_c97c0505,
        64'h282300c8_863b00d3,
        64'h06bb00fe_07bb010e,
        64'h883b6462_f3ff1de3,
        64'h00e587bb_0005869b,
        64'h0003861b_0f918f5d,
        64'h0157171b_00b7579b,
        64'h9f3d0077_47339fa1,
        64'h8f4dfff7_47130007,
        64'h081b00b3_85bb4080,
        64'h9fa18dd5_0115d59b,
        64'h94aa00f5_969b048a,
        64'h9db5ffc2_a4038db9,
        64'h02c10075_e5b3fff7,
        64'hc593023f_c4839ead,
        64'h00c703bb_00c3e633,
        64'h400c9ead_0166561b,
        64'h00a6139b_0082a583,
        64'h9e2d8e3d_8e59fff6,
        64'hc6139db1_00f8073b,
        64'h01076833_01a8581b,
        64'h0003a583_9e2d0068,
        64'h171b0107_083b0042,
        64'ha5839f2d_942a040a,
        64'h418c95aa_058a93aa,
        64'h038a020f_c5839f2d,
        64'h022fc403_021fc383,
        64'h0002a703_00d745b3,
        64'h8f5dfff6_47132462,
        64'h82930000_5297f45f,
        64'h17e300e4_07bb0004,
        64'h069b0005_861b0291,
        64'h8f5d0177_171b0097,
        64'h579b9f3d_8f219fa5,
        64'h8f2d0007_081b00d5,
        64'h843b8ec1_00092483,
        64'h0106d69b_9fa50106,
        64'h941b992a_9ea1090a,
        64'h8ead00e7_c6b3ffc3,
        64'ha4839c35_00c705bb,
        64'h03c18e4d_0156561b,
        64'h0132c903_00b6159b,
        64'h40809e2d_9ea194aa,
        64'h8db9048a_00f8073b,
        64'h0083a403_9e210107,
        64'h683301c8_581b0048,
        64'h171b0122_c4830107,
        64'h083b4080_9e2194aa,
        64'h048a0043_a4039f21,
        64'h0112c483_9f254000,
        64'h00c5c4b3_942a040a,
        64'h00d7c5b3_0003a703,
        64'h0102c403_2c438393,
        64'h00005397_82fe34ef,
        64'h8f930000_5f97f25f,
        64'h1ee300e4_07bb0004,
        64'h069b0003_861b0005,
        64'h881b8f5d_0147171b,
        64'h00c7579b_9f3d0077,
        64'h47338f6d_0083c733,
        64'h9fb900d3_843b8ec1,
        64'h40980126_d69b9fb9,
        64'h00e6941b_94aa048a,
        64'hffcfa703_9eb90fc1,
        64'h8eadffff_44838efd,
        64'h0075c6b3_0f119f35,
        64'h00c583bb_00c3e633,
        64'h40189eb9_0176561b,
        64'h0096139b_008fa703,
        64'h9e398e3d_8e7500b7,
        64'hc6339f31_00f805bb,
        64'h0105e833_0003a703,
        64'h01b8581b_9e390058,
        64'h159b0105_883b004f,
        64'ha7039db9_942a040a,
        64'h4318972a_070a93aa,
        64'h038a000f_47039db9,
        64'h002f4403_001f4383,
        64'h000fa583_00b6c733,
        64'h8df100d7_c5b342e2,
        64'h82930000_5297366f,
        64'h8f930000_5f9742ef,
        64'h0f130000_5f17f45f,
        64'h17e300e3_87bb0003,
        64'h869b0005_881b0f41,
        64'h8f5d0167_171b00a7,
        64'h579b9f3d_8f2d9fa1,
        64'h00777733_8f2d0007,
        64'h061b00d7_03bbffcf,
        64'ha4039fa1_00d3e6b3,
        64'h0116969b_00f6d39b,
        64'h007686bb_8ebd00cf,
        64'h24038ef9_00b7c6b3,
        64'h00d383bb_00c5873b,
        64'h008383bb_8e590146,
        64'h561b00c6_171b9e39,
        64'h008f2383_8e358e6d,
        64'h00f6c633_9f3100f8,
        64'h05bb0077_073b0105,
        64'he8330198_581b0078,
        64'h159b0105_883b004f,
        64'h2703ff4f_a3839db9,
        64'h007585bb_0fc1008f,
        64'ha403000f_2583000f,
        64'ha38300b6_47338dfd,
        64'h00c6c5b3_3ecf8f93,
        64'h00005f97_887687f2,
        64'h869a8646_04050293,
        64'h8f2ae44a_e826ec22,
        64'h110105c5_28830585,
        64'h23030545_2e030505,
        64'h2e83bf81_842abdd1,
        64'h00e785a3_47216786,
        64'ha8dfd0ef_082c462d,
        64'h6506ab7f_d0ef4581,
        64'h02000613_6506f835,
        64'h0005041b_a19fe0ef,
        64'h1028d3c1_01814783,
        64'h02f51b63_4791b771,
        64'h0005041b_8b2fe0ef,
        64'h00f50223_47857522,
        64'h00f50023_5795b7c5,
        64'h078500c6_802396be,
        64'h0834b77d_f0f713e3,
        64'h0e500793_01814703,
        64'h00d77963_0007869b,
        64'h02000613_47299381,
        64'h02061793_f8f6e9e3,
        64'h0007069b_00d58023,
        64'h070595ba_082cfe67,
        64'h02e3b7dd_ffc81be3,
        64'h00080563_0005c803,
        64'h05858082_61256446,
        64'h60e68522_4419feb0,
        64'h45e34185_d59b0185,
        64'h959ba831_00068e1b,
        64'h8f858593_00007597,
        64'h92c116c2_36810108,
        64'hec630308_58131842,
        64'hf9f6881b_92c10305,
        64'h96930017_061b0006,
        64'hc58300e5_06b3432d,
        64'h48e54701_fec686e3,
        64'h0006c683_96aa9281,
        64'h02071693_fff7871b,
        64'hb77d87ba_b7452785,
        64'ha0e900e7_8ca30007,
        64'h8ba30007_8b230460,
        64'h071300e7_8c230210,
        64'h07136786_bb1fd0ef,
        64'h082c462d_c7e56506,
        64'h01814783_10051563,
        64'h2501ac3f_e0ef1028,
        64'h4585e045_0005041b,
        64'hbccfe0ef_da021028,
        64'h4581ebb1_02000613,
        64'heb290007_4703972a,
        64'h93010207_97134781,
        64'h00010c23_6522e471,
        64'h0005041b_eddfd0ef,
        64'hec86e8a2_1028002c,
        64'h4605e42a_711db7d5,
        64'h842abf55_00048023,
        64'h00f51563_47918082,
        64'h61256906_64a66446,
        64'h60e68522_00a92023,
        64'hc15fd0ef_953e0347,
        64'h87930270_079300e6,
        64'h84630005_46830430,
        64'h0793470d_6562e015,
        64'h0005041b_e63fd0ef,
        64'h510c6562_02090a63,
        64'hfec783e3_177d0007,
        64'hc78397a6_93811782,
        64'h0007869b_fff6879b,
        64'hce890007_00230200,
        64'h061346ad_00b48713,
        64'hc8dfd0ef_8526462d,
        64'h75c2e93d_2501b97f,
        64'he0ef0828_4585e559,
        64'h2501c9ef_e0efd202,
        64'h08284581_c4b9e051,
        64'h0005041b_f95fd0ef,
        64'hec86e8a2_08284601,
        64'h002c8932_84aee42a,
        64'he0cae4a6_711d8082,
        64'h61256446_60e62501,
        64'hacefe0ef_00f50223,
        64'h478500e7_8ca30087,
        64'h571b00e7_8c230044,
        64'h570300e7_8ba30087,
        64'h571b00e7_8b237522,
        64'h00645703_cb856786,
        64'heb950207_f79300b7,
        64'hc7834519_67a6e129,
        64'h250199df_e0efe4be,
        64'h1028083c_65a2e929,
        64'h250180af_e0efec86,
        64'h1028002c_4605842e,
        64'he42ae8a2_711dbfcd,
        64'h47a18082_614d853e,
        64'h64ea740a_70aa0005,
        64'h079bb48f_e0ef6506,
        64'he7910005_079be18f,
        64'he0ef0088_00f70223,
        64'h06d707a3_478506f7,
        64'h04a30086_d69b0106,
        64'hd69b0087_d79b0107,
        64'hd79b0107_979b06f7,
        64'h04230107_d79b06f7,
        64'h07230107_969b57d6,
        64'h02f69c63_05574683,
        64'h02e00793_6706efa9,
        64'h0005079b_fbbfd0ef,
        64'h8522c1bd_47890005,
        64'h059bca4f_e0ef8522,
        64'h0005059b_f25fd0ef,
        64'h85a60004_450306f7,
        64'h076357d6_4736cbb5,
        64'h8bc100b4_c78300f4,
        64'h02234785_00f485a3,
        64'h0207e793_64060281,
        64'h4783df7f_d0ef00d4,
        64'h851302a1_0593464d,
        64'h648aebdd_0005079b,
        64'hdcbfe0ef_10a80ce7,
        64'h92634711_cbf10005,
        64'h079ba9df_e0ef10a8,
        64'h65820c05_4c6347ad,
        64'hefdfd0ef_850ae33f,
        64'hd0ef10a8_008c0280,
        64'h0613e3ff_d0ef1028,
        64'h05ad4655_0e058d63,
        64'h479165e6_10071163,
        64'h02077713_479900b7,
        64'hc7037786_10079963,
        64'h0005079b_ae7fe0ef,
        64'hf0be083c_f4be0088,
        64'h65a26786_12079563,
        64'h0005079b_95cfe0ef,
        64'hed26f122_f5060088,
        64'h002c4605_e02ee42a,
        64'h71718082_616564e6,
        64'h740670a6_2501c94f,
        64'he0ef00f5_02234785,
        64'h008705a3_8c3d0274,
        64'h74138c65_8cbd7522,
        64'h00b74783_c30d6706,
        64'he39d0207_f79300b7,
        64'hc7834519_67a6e915,
        64'h2501b55f_e0efe4be,
        64'h1028083c_65a2e131,
        64'h25019c2f_e0eff486,
        64'h10284605_002c8432,
        64'h84aee42a_eca6f0a2,
        64'h7159b7c5_44218082,
        64'h614d6d46_6ce67c06,
        64'h7ba67b46_7ae66a0a,
        64'h69aa694a_64ea740a,
        64'h70aa8522_f2bfe0ef,
        64'h85a67522_441db749,
        64'h8c6a0ffb_fb93f53f,
        64'hd0ef3bfd_855a4581,
        64'h20000613_ec090005,
        64'h041b8d4f_e0ef0195,
        64'h02230385_2823001c,
        64'h0d1b7522_a82d0005,
        64'h041bd50f_e0ef00f5,
        64'h02234785_01278aa3,
        64'h01578a23_01378da3,
        64'h01478d23_00e78ca3,
        64'h00078ba3_00078b23,
        64'h04600713_00e78c23,
        64'h02100713_00e785a3,
        64'h75224741_6786e835,
        64'h0005041b_f5ffe0ef,
        64'h1028040b_99634c85,
        64'h00274b83_06f404a3,
        64'h06d407a3_0087d79b,
        64'h0086d69b_0107d79b,
        64'h0106d69b_0107979b,
        64'h06f40423_0107d79b,
        64'h0107969b_06f40723,
        64'h478100f6_93635714,
        64'h00d61663_57d20007,
        64'h4603468d_05740aa3,
        64'h7722ff7f_d0ef0544,
        64'h051385da_052404a3,
        64'h05540423_053407a3,
        64'h05440723_040405a3,
        64'h04040523_03740a23,
        64'h02000613_04f406a3,
        64'h0089591b_0089d99b,
        64'h04600793_0ff4fa13,
        64'h04f40623_02e00b93,
        64'h0109591b_02100793,
        64'h0109d99b_02f40fa3,
        64'h0109191b_0104999b,
        64'h0ff97a93_47c187af,
        64'he0ef855a_02000593,
        64'h462d886f_e0ef855a,
        64'h00050c1b_45812000,
        64'h06130344_0b13f60f,
        64'he0ef8522_0104d91b,
        64'h85a67422_16041263,
        64'h0005041b_a8cfe0ef,
        64'h16f48863_440557fd,
        64'h16f48c63_44097522,
        64'h47851804_80630005,
        64'h049bb33f_e0ef4581,
        64'h75221807_9d630207,
        64'hf79300b7_c7834419,
        64'h67a61af4_15634791,
        64'h1c040763_0005041b,
        64'hd53fe0ef_e4be1028,
        64'h083c65a2_1c041263,
        64'h0005041b_bc4fe0ef,
        64'he8eaece6_f0e2f4de,
        64'hf8dafcd6_e152e54e,
        64'he94aed26_f506f122,
        64'h1028002c_4605e42a,
        64'h7171b7ed_f5512501,
        64'h91eff0ef_85a27502,
        64'hbf612501_f12fe0ef,
        64'h7502e411_f1552501,
        64'h9e3fe0ef_1008faf5,
        64'h18e34791_d94d2501,
        64'h838ff0ef_00a84581,
        64'hf1612501_941fe0ef,
        64'hcaa200a8_4589952f,
        64'he0ef00a8_100c0280,
        64'h0613fc87_8de30149,
        64'h2783c89d_88c1cc0d,
        64'h0005041b_accfe0ef,
        64'h00094503_79028082,
        64'h61497946_74e6640a,
        64'h60aa451d_cb810014,
        64'hf79300b5_c483c599,
        64'h75e2eb89_0207f793,
        64'h00b7c783_45196786,
        64'he1052501_e27fe0ef,
        64'he0be1008_081c65a2,
        64'he9052501_c94fe0ef,
        64'hf8cafca6_e122e506,
        64'h1008002c_4605e42a,
        64'h7175b7b1_00f40523,
        64'hfbf7f793_00a44783,
        64'hf55d2501_67a040ef,
        64'h03040593_0017c503,
        64'h46854c50_601cdba5,
        64'h0407f793_00a44783,
        64'hfcf96ae3_4d1c6008,
        64'hfcf900e3_45094785,
        64'hb769449d_b7e12501,
        64'ha1eff0ef_85ca6008,
        64'hf9792501_b25fe0ef,
        64'h167d1000_06374c0c,
        64'hb7dd4505_02f91463,
        64'h57fd0005_091b941f,
        64'he0ef4c0c_bf7d84aa,
        64'h00a405a3_c5390004,
        64'h2a232501_a5aff0ef,
        64'h484cef01_600800f4,
        64'h0523c818_0207e793,
        64'hfed772e3_48144458,
        64'hcf390027_f71300a4,
        64'h47838082_610564a2,
        64'h69028526_644260e2,
        64'h0007849b_cb9100b4,
        64'h4783e491_0005049b,
        64'hbb8fe0ef_842ae04a,
        64'hec06e426_e8221101,
        64'hbfad8a2a_bfbd4a09,
        64'hb7494a05_b7c539f1,
        64'h09112485_e1116582,
        64'h01557533_2501aa2f,
        64'he0efe02e_854ab745,
        64'hfc0c94e3_3cfd39f9,
        64'h09092485_e3918fd9,
        64'h0087979b_00094703,
        64'h00194783_038b9163,
        64'h20000993_03440913,
        64'h85cee921_2501d04f,
        64'he0ef0015_899b8522,
        64'h00099e63_1afd4c09,
        64'h44814981_49011000,
        64'h0ab7504c_b74d009b,
        64'h202300f4_02a30017,
        64'he793c804_00544783,
        64'hfef963e3_29054c1c,
        64'h2485e111_09550863,
        64'h09350863_2501a49f,
        64'he0ef8522_85ca4a85,
        64'h59fd4481_490902fb,
        64'h9f634785_00044b83,
        64'h80826165_6ce27c02,
        64'h7ba27b42_7ae26a06,
        64'h69a66946_64e68552,
        64'h740670a6_00fb2023,
        64'h02f76263_ffec871b,
        64'h481c0184_2c836000,
        64'h000a1c63_00050a1b,
        64'he70fe0ef_ec66f062,
        64'hf45efc56_e4cee8ca,
        64'heca6f486_e0d28522,
        64'h002c4601_8b2ee42a,
        64'hf85a8432_f0a27159,
        64'hbfcd4419_80826165,
        64'h64e67406_70a68522,
        64'hc00fe0ef_102885a6,
        64'hc489cf81_6786e801,
        64'h0005041b_85eff0ef,
        64'he4be1028_083c65a2,
        64'he00d0005_041becef,
        64'he0eff486_f0a21028,
        64'h002c4601_84aee42a,
        64'heca67159_bf6584aa,
        64'hd16dbf7d_00042a23,
        64'h00f51663_47912501,
        64'hf77fe0ef_85224581,
        64'hc58fe0ef_852285ca,
        64'h00042a23_02f51363,
        64'h47912501_b34ff0ef,
        64'h85224581_02243023,
        64'h80826145_64e26942,
        64'h85267402_70a20005,
        64'h049bc4ff_e0ef8522,
        64'h45810009_1f63e889,
        64'h0005049b_d8cfe0ef,
        64'h892e842a_f406e84a,
        64'hec26f022_71798082,
        64'h01416402_60a20004,
        64'h3023e119_2501daef,
        64'he0ef842a_e406e022,
        64'h1141b7c1_fcf501e3,
        64'h4791bfdd_45258082,
        64'h61217442_70e2f971,
        64'hfcf50be3_47912501,
        64'hcadfe0ef_00f41423,
        64'h0067d783_85224581,
        64'h67e2c448_e24fe0ef,
        64'h0007c503_67e2a02d,
        64'h00043023_4515e789,
        64'h8bc100b5_c783cd99,
        64'h6c0ce529_2501968f,
        64'hf0eff01c_101ce01c,
        64'h852265a2_67e2e115,
        64'h2501fdaf_e0ef0828,
        64'h002c4601_842ac52d,
        64'he42ef822_fc067139,
        64'hb7bdc45c_013787bb,
        64'h413484bb_cc0c445c,
        64'hfaf5fae3_4f9c601c,
        64'hfabafee3_fd4588e3,
        64'h0005059b_c3ffe0ef,
        64'hbf6984ce_e5990005,
        64'h059bfcbf_e0efcb81,
        64'h8b896008_00a44783,
        64'hb765cc0c_c84cb5ed,
        64'h490500f4_05a34785,
        64'h00f59763_57fdbded,
        64'h490900f4_05a34789,
        64'h00f59763_47850005,
        64'h059b802f_f0efe595,
        64'h484cbfb1_9ca90094,
        64'hd49bcd11_2501c79f,
        64'he0ef6008_d7b51ff4,
        64'hf793c45c_9fa5445c,
        64'h0499ea63_4a855a7d,
        64'hd1c19c9d_c45c2781,
        64'h4c0c8ff9_413007bb,
        64'h02c6ed63_0337563b,
        64'h0336d6bb_fff4869b,
        64'h377dc729_0097999b,
        64'h00254783_6008bf59,
        64'hcc44ed35_250124b0,
        64'h40ef85ce_0017c503,
        64'h86264685_601c00f4,
        64'h0523fbf7_f79300a4,
        64'h4783ed51_250129d0,
        64'h40ef0017_c50385ce,
        64'h4685601c_c3850407,
        64'hf7930304_099300a4,
        64'h4783fc96_0ee34c50,
        64'hd3e51ff7_f793445c,
        64'h4481bf7d_00f40523,
        64'h0207e793_00a44783,
        64'hc81cfcf7_78e34818,
        64'h445ce4bd_00042623,
        64'h445884ba_e3918b89,
        64'h00a44783_00977763,
        64'h48188082_61216aa2,
        64'h6a4269e2_790274a2,
        64'h854a7442_70e20007,
        64'h891bcf89_00b44783,
        64'h00091763_0005091b,
        64'hfa8fe0ef_84ae842a,
        64'he456e852_ec4efc06,
        64'hf04af426_f8227139,
        64'hb721fe94_65e3fee7,
        64'h8fa32405_07850007,
        64'h47039736_92810204,
        64'h16936722_0789bdf5,
        64'h4545b7e9_00e60023,
        64'hfc974703_972a1088,
        64'h93011702_0007059b,
        64'hfff5871b_b7e12785,
        64'hbf199c3d_01260023,
        64'hfff7c793_e989963a,
        64'h93010206_97136622,
        64'h36fd86a2_85be04e4,
        64'h60630037_871be705,
        64'hfc974703_97361094,
        64'h93010207_97134781,
        64'hf48fe0ef_1828100c,
        64'hb7614509_f6e512e3,
        64'h67a24711_dd612501,
        64'ha86ff0ef_18284581,
        64'h01350e63_2501897f,
        64'he0ef0007_c50365c6,
        64'h77e2e105_2501e46f,
        64'hf0ef1828_4581f951,
        64'h2501f4ff_e0ef1828,
        64'h4581c2aa_8bdfe0ef,
        64'h0007c503_65c677e2,
        64'hf55d2501_e6cff0ef,
        64'h18284581_fd4d2501,
        64'hf75fe0ef_18284585,
        64'h80826149_79a67946,
        64'h74e6640a_60aa0007,
        64'h8023078d_00e78123,
        64'h02f00713_0e941563,
        64'h00e780a3_03a00713,
        64'h00e78023_0307071b,
        64'h3d874703_00008717,
        64'he50567a2_45010409,
        64'h91634996_c2be4bdc,
        64'h02f00913_842677e2,
        64'hecbe081c_e5212501,
        64'hab9fe0ef_1828002c,
        64'h460184ae_00050023,
        64'hf4cef8ca_e122e506,
        64'he42afca6_7175bfd9,
        64'h4415fcf4_1ee34791,
        64'hb7c5c8c8_965fe0ef,
        64'h0004c503_74a2cb99,
        64'h8bc100b5_c7838082,
        64'h616564e6_740670a6,
        64'h8522cbd8_575277a2,
        64'he9916586_e41d0005,
        64'h041bcb4f_f0efe4be,
        64'h1028083c_65a2ec19,
        64'h0005041b_b25fe0ef,
        64'heca6f486_f0a21028,
        64'h002c4601_e42a7159,
        64'hbfe5452d_80826105,
        64'h60e24501_48a78623,
        64'h00008797_00054a63,
        64'h945fe0ef_ec060028,
        64'he42a1101_80820141,
        64'h640260a2_00043023,
        64'he1192501_9b5fe0ef,
        64'h8522e901_2501f01f,
        64'hf0ef842a_e406e022,
        64'h11418082_01416402,
        64'h60a24505_ea3fe06f,
        64'h014160a2_640200f5,
        64'h02234785_00f40523,
        64'hfdf7f793_600800a4,
        64'h47830007_89a30007,
        64'h892300e7_8ca300d7,
        64'h8da30460_07130086,
        64'hd69b00e7_8c230210,
        64'h07130106_d69b00e7,
        64'h8aa30087_571b0107,
        64'h571b0107_171b00e7,
        64'h8a230107_571b0107,
        64'h169b00e7_8d230007,
        64'h8ba30007_8b234858,
        64'h00e78fa3_00d78f23,
        64'h0187571b_0107569b,
        64'h00d78ea3_00e78e23,
        64'h0086d69b_0106d69b,
        64'h0107169b_481800e7,
        64'h85a30207_671300b7,
        64'hc703741c_e1552501,
        64'hb5ffe0ef_6008500c,
        64'h00f40523_fbf7f793,
        64'h00a44783_ed4d2501,
        64'h607040ef_03040593,
        64'h0017c503_46854c50,
        64'h601cc395_0407f793,
        64'hcf610207_f71300a4,
        64'h4783e16d_2501ab7f,
        64'he0ef842a_e406e022,
        64'h1141bd15_499db5f1,
        64'hc81cbf41_00f40523,
        64'h0407e793_00a44783,
        64'h9b5fe0ef_952285d2,
        64'h86260305_05130007,
        64'h049b0127_746340ab,
        64'h873b1ff5_75130009,
        64'h049b4448_01b42e23,
        64'hfd012501_649040ef,
        64'h85da4685_0017c503,
        64'h00d77a63_44584814,
        64'h00c70e63_4c58bdc9,
        64'h00faa023_9fa5000a,
        64'ha783c45c_9fa54099,
        64'h093b445c_9a3e9381,
        64'h02049793_0094949b,
        64'h00f40523_fbf7f793,
        64'h00a44783_a29fe0ef,
        64'h855a95d2_20000613,
        64'h91811582_0097959b,
        64'h0297f263_41b587bb,
        64'h4c4cf149_25016e50,
        64'h40ef85d2_86a60017,
        64'hc50341a6_84bb00e6,
        64'hf4630104_873b0099,
        64'h549b0027_c683072c,
        64'h7a6367a2_8db200a8,
        64'h063b000d_081bd159,
        64'h2501964f_f0efe43e,
        64'h853e4c0c_601c00f4,
        64'h0523fbf7_f79300a4,
        64'h4783f969_25017350,
        64'h40ef85da_0017c503,
        64'h46854c50_601cc38d,
        64'h0407f793_00a44783,
        64'hc85ce311_cc1c4858,
        64'hbf894985_00f405a3,
        64'h47850197_9763b785,
        64'h00f40523_0207e793,
        64'h00a44783_12f76b63,
        64'h4818445c_f3fd0005,
        64'h079bd6af_f0ef4c0c,
        64'hb7494989_00f405a3,
        64'h478902e7_98634705,
        64'hcb914581_485cef01,
        64'h040d1a63_0ffd7d13,
        64'h01a7fd33_37fd0025,
        64'h47830097_5d1b6008,
        64'h14079463_1ff77793,
        64'h04090463_44585cfd,
        64'h03040b13_1ff00c13,
        64'h20000b93_04f76e63,
        64'h0127873b_445c1a07,
        64'h82638b89_00a44783,
        64'h80826109_6de27d02,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e67906,
        64'h74a6854e_744670e6,
        64'h0007899b_c39d00b4,
        64'h47830009_97630005,
        64'h099bca3f_e0ef8ab6,
        64'h89328a2e_842a0006,
        64'ha023ec6e_f06af466,
        64'hf862fc5e_e0daf4a6,
        64'hfc86e4d6_e8d2ecce,
        64'hf0caf8a2_7119b585,
        64'h499dbf9d_bb1fe0ef,
        64'h855295a2_86260305,
        64'h85930007_049b0127,
        64'h746340bb_873b1ff5,
        64'hf5930009_049b444c,
        64'h01b42e23_f10d2501,
        64'h044050ef_85da0017,
        64'hc5038642_4685601c,
        64'h00f40523_fbf7f793,
        64'h682200a4_4783f131,
        64'h25010980_50efe442,
        64'h85da4685_0017c503,
        64'hc30d0407_771300a4,
        64'h47030506_01634c50,
        64'hbf3900fa_a0239fa5,
        64'h000aa783_c45c9fa5,
        64'h4099093b_445c9a3e,
        64'h93810204_97930094,
        64'h949bc3ff_e0ef9552,
        64'h85da2000_06139101,
        64'h15020097_951b0097,
        64'hfc6341b5_07bb4c48,
        64'hc3850407_f79300a4,
        64'h4783f945_25010d20,
        64'h50ef85d2_864286a6,
        64'h0017c503_41a684bb,
        64'h00e6f463_00c4873b,
        64'h0099549b_0027c683,
        64'h072c7a63_67a28dc2,
        64'h00a6083b_000d061b,
        64'hd5792501_b86ff0ef,
        64'he43e853e_4c0c601c,
        64'hcc08b795_498500f4,
        64'h05a34785_01951763,
        64'hb7e52501_bc6ff0ef,
        64'h4c0cbfb5_498900f4,
        64'h05a34789_00a7ec63,
        64'h47854848_eb11020d,
        64'h19630ffd_7d1301a7,
        64'hfd3337fd_00254783,
        64'h00975d1b_60081207,
        64'h91631ff7_77934458,
        64'hfa090ae3_5cfd0304,
        64'h0b131ff0_0c132000,
        64'h0b930006_091b00f6,
        64'h7463893e_40f907bb,
        64'h445c0104_29031607,
        64'h8c638b85_00a44783,
        64'h80826109_6de27d02,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e67906,
        64'h74a6854e_744670e6,
        64'h0007899b_c39d6622,
        64'h00b44783_00099863,
        64'h0005099b_e85fe0ef,
        64'h8ab6e432_8a2e842a,
        64'h0006a023_ec6ef06a,
        64'hf466f862_fc5ee0da,
        64'hf0caf4a6_fc86e4d6,
        64'he8d2ecce_f8a27119,
        64'hbdd14525_bf51ec07,
        64'h9ee3451d_8b85fa09,
        64'h00e30029_7913ee07,
        64'h16e30107_f7134511,
        64'h00b44783_ee051de3,
        64'hbdf54501_00f49423,
        64'h0124b023_0004ae23,
        64'h0004a623_c8880069,
        64'h5783daff_e0ef01c4,
        64'h0513c8c8_f35fe0ef,
        64'h00094503_000485a3,
        64'hd09c0134_8523f480,
        64'h03092783_85a27922,
        64'h0209e993_c3990089,
        64'hf793f139_250180cf,
        64'hf0ef0125_262385d6,
        64'h397d7522_fd212501,
        64'he1fff0ef_030a2a83,
        64'h855285ca_02090363,
        64'h00fa0223_0005091b,
        64'h00040aa3_00040a23,
        64'h00040da3_00040d23,
        64'h4785f9bf_e0ef85a2,
        64'h000a4503_00040fa3,
        64'h00040f23_00040ea3,
        64'h00040e23_000405a3,
        64'h00e40c23_00040ba3,
        64'h00040b23_00e40823,
        64'h000407a3_00040723,
        64'h00f40ca3_00f408a3,
        64'h02100713_04600793,
        64'h7a220089_e9936406,
        64'ha0210809_0a630089,
        64'h7913fff9_45210049,
        64'h7793f3fd_8bc5451d,
        64'h00b44783_80826149,
        64'h6ae67a06_79a67946,
        64'h74e6640a_60aac905,
        64'h2501e7df_f0ef1028,
        64'h00f51763_4791c115,
        64'h10078e63_01f97993,
        64'h01c97793_4519e011,
        64'he1196406_2501b61f,
        64'hf0efe4be_1028083c,
        64'h65a2e91d_25019cef,
        64'hf0ef1028_002c8a79,
        64'h84aa8932_00053023,
        64'h16050c63_e42eecd6,
        64'hf0d2f4ce_f8cafca6,
        64'he122e506_7175bfe5,
        64'h452d8082_612170e2,
        64'h2501a02f_f0ef0828,
        64'h080c4601_00f61863,
        64'h4785cb11_4501e398,
        64'h97aa0007_0023c319,
        64'h67620007_0023c319,
        64'h66226318_00a78733,
        64'h050eb6a7_87930000,
        64'h97970405_4263832f,
        64'hf0eff42e_e432e82e,
        64'hfc061028_ec2a7139,
        64'h80824509_bf4d4505,
        64'hbf5d4509_bf65faf4,
        64'he7e30004_891b4c1c,
        64'h00f402a3_0017e793,
        64'h00544783_c81c2785,
        64'h01378a63_481cfd71,
        64'h25018abf_f0ef8522,
        64'h85ca4601_03348c63,
        64'h03448c63_80826145,
        64'h6a0269a2_694264e2,
        64'h740270a2_4501e891,
        64'h0005049b_ed6ff0ef,
        64'h852285ca_59fd4a05,
        64'h06f5f063_892e842a,
        64'he052e44e_ec26f406,
        64'he84af022_71794d1c,
        64'h08b7f063_47858082,
        64'h610564a2_85266442,
        64'h60e200e7_82234705,
        64'h601c80ef_f0ef462d,
        64'h6c08700c_838ff0ef,
        64'h45810200_06136c08,
        64'he0850005_049ba34f,
        64'hf0ef6008_484ce49d,
        64'h0005049b_fa9ff0ef,
        64'h842aec06_e426e822,
        64'h11018082_610564a2,
        64'h644260e2_451d00f5,
        64'h13634791_dd792501,
        64'hbb7ff0ef_85224585,
        64'hcb990097_8d630007,
        64'hc7836c1c_ed092501,
        64'ha7eff0ef_6008484c,
        64'h0e500493_e50d2501,
        64'h87dff0ef_842ae426,
        64'hec06e822_45811101,
        64'hbfe54511_b7cd0004,
        64'h2a23d945_2501bfdf,
        64'hf0ef8522_45818082,
        64'h614569a2_694264e2,
        64'h740270a2_45010097,
        64'h9a630017_b79317e1,
        64'h8bfd0337_80630327,
        64'h026303f7_f79300b7,
        64'hc783c321_0007c703,
        64'h6c1ce129_2501aecf,
        64'hf0ef6008_a0b1c90d,
        64'he199484c_49bd0e50,
        64'h09134511_84aef406,
        64'h842ae44e_e84aec26,
        64'hf0227179_bdc10ff7,
        64'h77130017_e7933701,
        64'heca8efe3_0ff57513,
        64'hf9f7051b_eea8f3e3,
        64'h0ff57513_fbf7051b,
        64'hb5754519_ef0719e3,
        64'h00080663_00054803,
        64'hee050513_00008517,
        64'h00054c63_4185551b,
        64'h0187151b_02b6f263,
        64'hfd370ae3_f35709e3,
        64'hf3470be3_f2e37de3,
        64'h00074703_97229301,
        64'h17020017_061b8732,
        64'h45ad46a1_0ff7f793,
        64'h0027979b_05659a63,
        64'hb5a1c4c8_ae4ff0ef,
        64'h0007c503_609cdbe5,
        64'h8bc100b5_c7836c8c,
        64'hfbe58b91_b7054515,
        64'hf315bfd9_4511b72d,
        64'h4501e607_0ae30004,
        64'hbc230004_a623cb99,
        64'h0207f793_0047f713,
        64'hf4e513e3_4711c515,
        64'h00b7c783_709cf127,
        64'h9de3b7c5_01066613,
        64'hfed714e3_46850037,
        64'hf713bded_00c905a3,
        64'h00866613_00e79463,
        64'h47118bb1_0ff7f793,
        64'h0027979b_01659f63,
        64'h00e90023_471500e6,
        64'h95630e50_07130009,
        64'h4683c6e5_460100e5,
        64'h73634611_94320200,
        64'h05139201_1602a865,
        64'h268500e5_0023954a,
        64'h91010206_95130027,
        64'he793a211_0505a8c9,
        64'h48e50200_03134781,
        64'h45a14701_4681b78d,
        64'h02400793_943a12f6,
        64'he7630200_0693f757,
        64'h87e3b7b5_4709b73d,
        64'h04058082_61216b02,
        64'h6aa26a42_69e27902,
        64'h74a27442_70e20004,
        64'hbc232501_a81ff0ef,
        64'h85264581_bf35c55c,
        64'h4bdc611c_a0e1dd5d,
        64'h2501df9f_f0ef8526,
        64'h45810cd6_0a63fff6,
        64'h46030006_c68300f5,
        64'h86330785_00f706b3,
        64'h708cef89_8ba100b7,
        64'h47831207_80630007,
        64'h47836c98_10051163,
        64'h2501ce0f_f0ef6088,
        64'h48cc492d_10051963,
        64'h2501adff_f0ef8526,
        64'h458100f9_05a30200,
        64'h0793943a_09479b63,
        64'h470d1d37_89630024,
        64'h478300f9_00a302e0,
        64'h07930b37_94630014,
        64'h47830139_00230d37,
        64'h96630004_4783b42f,
        64'hf0ef854a_02000593,
        64'h462d0204_b9030d57,
        64'h84630d47_86630004,
        64'h47834b21_02e00993,
        64'h05c00a93_02f00a13,
        64'h0ce7f063_47fd0004,
        64'h47030004_a6230405,
        64'h0ce79463_05c00713,
        64'h00e78663_842e84aa,
        64'h02f00713_0005c783,
        64'he05ae456_e852ec4e,
        64'hf04afc06_f426f822,
        64'h7139b7e9_db1c2785,
        64'h5b1c2a85_6018f141,
        64'h2501d24f_f0ef0145,
        64'h0223b7b9_c848a89f,
        64'hf0ef85a6_c8046008,
        64'hd91c4157_87bb591c,
        64'h00faed63_00254783,
        64'h60084a05_02aa2823,
        64'haabff0ef_855285a6,
        64'h00043a03_bf0ff0ef,
        64'h03450513_45812000,
        64'h06136008_f5792501,
        64'hde0ff0ef_6008fcf4,
        64'h8de357fd_fcf48be3,
        64'h4785d4bd_451d0005,
        64'h049be83f_f0ef480c,
        64'hf60a0ee3_06f4e063,
        64'h4d1c6008_b7614505,
        64'h00f49463_57fdbf49,
        64'h45090097_e4634785,
        64'h0005049b_b2fff0ef,
        64'hfc0a9fe3_0157fab3,
        64'h37fd0049_5a9b0025,
        64'h4783bf5d_4501ec1c,
        64'h97ce0347_87930124,
        64'h15230996_601cfcf7,
        64'h75e30009_071b0085,
        64'h5783e18d_c85c6108,
        64'h2785480c_00099d63,
        64'h842a8a2e_00f97993,
        64'hd7ed495c_80826121,
        64'h6aa26a42_69e27902,
        64'h74a27442_70e24511,
        64'heb9993c1_e456e852,
        64'hec4ef426_03091793,
        64'h2905f822_fc0600a5,
        64'h5903f04a_7139b795,
        64'h547df6f5_14e34785,
        64'hdd612501_dbdff0ef,
        64'h852685ce_8622bfb5,
        64'h00f482a3_0017e793,
        64'h0054c783_c89c37fd,
        64'hf8e788e3_577dc4c0,
        64'h489c0209_9063e905,
        64'h2501debf_f0ef8526,
        64'h85a2167d_10000637,
        64'hb7cdfd24_1de3fb45,
        64'h0ae30555_0a63c901,
        64'h2501c0df_f0ef8526,
        64'h85a24409_b7e94401,
        64'h012a6463_00f46763,
        64'h24054c9c_5afd4a05,
        64'h844afef4_61e3894e,
        64'h4c9c08f4_026357fd,
        64'h80826121_6aa26a42,
        64'h69e27902_74a27442,
        64'h70e28522_44050087,
        64'hed634785_0005041b,
        64'hc5bff0ef_a8154905,
        64'h02f96d63_4d1c0009,
        64'h056300c5_2903e991,
        64'h89ae84aa_e456e852,
        64'hf04af822_fc06ec4e,
        64'hf4267139_bf79012a,
        64'h81a300fa_81230189,
        64'h591b0109_579b00fa,
        64'h80a30087_d79b0324,
        64'h0a230107_d79b9426,
        64'h0109179b_29010125,
        64'h69338d71_f0000637,
        64'h2501d96f_f0ef8556,
        64'h9aa60344_0a931fc4,
        64'h74130024_141bf80a,
        64'h16e30005_0a1bfdcf,
        64'hf0ef9dbd_0075d59b,
        64'h515cbf79_01348223,
        64'h03240aa3_0089591b,
        64'h0109591b_0109191b,
        64'h03240a23_94261fe4,
        64'h74130014_141bfc0a,
        64'h12e30005_0a1b815f,
        64'hf0ef9dbd_0085d59b,
        64'h515cb7e9_0127e933,
        64'h9bc100f9_79130089,
        64'h591b0347_c7830154,
        64'h87b38082_61216aa2,
        64'h6a4269e2_790274a2,
        64'h85527442_70e200f4,
        64'h82234785_032a8a23,
        64'h9aa60ff9_79130049,
        64'h591bc40d_1ffafa93,
        64'h000a1f63_00050a1b,
        64'h86fff0ef_9dbd8526,
        64'h009ad59b_50dc00f4,
        64'h82234785_02f98a23,
        64'h99a60ff7_f7938fd9,
        64'h8ff50049_179b00f7,
        64'hf71316c1_66850347,
        64'hc7830134_87b3cc19,
        64'h1ff9f993_0ff97793,
        64'h00198a9b_8805060a,
        64'h16630005_0a1b8bdf,
        64'hf0ef9dbd_0099d59b,
        64'h00b989bb_515c0015,
        64'hd99b0937_94630ee7,
        64'h8863470d_0ae78f63,
        64'h842e8932_47090005,
        64'h47830af5_f0634a09,
        64'h84aa4d1c_0ab9f563,
        64'h4a094985_e456f04a,
        64'hf426f822_fc06e852,
        64'hec4e7139_80826105,
        64'h64a28526_644260e2,
        64'h00e78223_4705601c,
        64'h00e78023_57156c1c,
        64'hf3cff0ef_45810200,
        64'h06136c08_ec990005,
        64'h049b939f_f0ef6008,
        64'h484ce495_0005049b,
        64'hf35ff0ef_842aec06,
        64'he426e822_110100a5,
        64'h5583b795_4505bfc1,
        64'h4134043b_f6f4f7e3,
        64'h4f9c0009_3783f69a,
        64'hfce30144_8c630005,
        64'h049be75f_f0efbf7d,
        64'h2501e5df_f0ef0134,
        64'h766385a6_00093503,
        64'h09924a85_5a7d0027,
        64'hc98384ba_b75d4501,
        64'h00893c23_943e0347,
        64'h87930416_883d0009,
        64'h378300f9_2a239fa9,
        64'h0044579b_d1710099,
        64'h28235788_fce477e3,
        64'h0087d703_eb0d5798,
        64'h00e69463_470d0007,
        64'hc683e0a9_842efee4,
        64'hf4e34f98_611c8082,
        64'h61216aa2_6a4269e2,
        64'h790274a2_744270e2,
        64'h450900f4_9c63892a,
        64'h478500b5_1523e456,
        64'he852ec4e_f822fc06,
        64'hf04a4544_f4267139,
        64'h8082853e_4785bfb9,
        64'h02455793_1512ffaf,
        64'hf0ef954a_03450513,
        64'h1fc57513_0024151b,
        64'hf93d2501_a3bff0ef,
        64'h9dbd0075_d59b515c,
        64'hb7618fc9_0087979b,
        64'h03494503_03594783,
        64'h99221fe4_74130014,
        64'h141bf145_2501a65f,
        64'hf0ef9dbd_0085d59b,
        64'h515cbf4d_93d117d2,
        64'hbf658391_c0198fc5,
        64'h0087979b_88050349,
        64'h4783994e_1ff9f993,
        64'hf5792501_a93ff0ef,
        64'h0344c483_854a9dbd,
        64'h94ca1ff4_f4930099,
        64'hd59b0014_899b0249,
        64'h27838082_6145853e,
        64'h69a26942_64e27402,
        64'h70a257fd_c9112501,
        64'hac7ff0ef_9dbd0094,
        64'hd59b9cad_515c0015,
        64'hd49b00f7_1e6308d7,
        64'h0d63468d_06d70b63,
        64'h842e4689_00054703,
        64'h02e5f963_892ae44e,
        64'hec26f022_f406e84a,
        64'h71794d18_0eb7f563,
        64'h47858082_45018082,
        64'h9d3d02b7_87bb5548,
        64'h00254783_00e7f963,
        64'h377985be_ffe5879b,
        64'h4d188082_610564a2,
        64'h644260e2_00a03533,
        64'h25015cd0_50ef4581,
        64'h46010014_45030004,
        64'h02a35d90_50ef85a6,
        64'h4685d810_22f401a3,
        64'h22e40123_20d40ca3,
        64'h20d40c23_0187d79b,
        64'h0107d71b_260522e4,
        64'h00a322f4_00230720,
        64'h06930014_45030087,
        64'h571b0107_571b0107,
        64'h971b5010_20e40f23,
        64'h445c20f4_0fa30187,
        64'hd79b0107_d71b20e4,
        64'h0ea320f4_0e230087,
        64'h571b0107_571b0107,
        64'h971b20e4_0d2302e4,
        64'h0ba30410_0713481c,
        64'h20f40da3_02f40b23,
        64'h06100793_02f40aa3,
        64'h02f40a23_05200793,
        64'h22f409a3_faa00793,
        64'h22f40923_05500793,
        64'h9fdff0ef_85264581,
        64'h20000613_03440493,
        64'h0af71b63_47850054,
        64'h47030cf7_1063478d,
        64'h00044703_ed692501,
        64'hc01ff0ef_842ae426,
        64'hec06e822_1101bdcd,
        64'h9cbd0017_d79b8885,
        64'h029787bb_478db709,
        64'h0014949b_00f91563,
        64'h4789d41c_9fb5e00a,
        64'h84e3b545_a19ff0ef,
        64'h05440513_b5b10005,
        64'h099ba27f_f0ef0584,
        64'h0513b351_47810004,
        64'h2a230124_002300f4,
        64'h132368f7_12230000,
        64'h971793c1_17c22785,
        64'h6927d783_00009797,
        64'hc448a57f_f0ef2204,
        64'h0513c808_a61ff0ef,
        64'h21c40513_00f51c63,
        64'h27278793_25016141,
        64'h77b7a77f_f0ef2184,
        64'h051302f5_17632527,
        64'h87932501_416157b7,
        64'ha8dff0ef_03440513,
        64'h04e79263_a5570713,
        64'h4107d79b_776d0107,
        64'h979b8fd9_0087979b,
        64'h000402a3_23244703,
        64'h23344783_e13d2501,
        64'hce7ff0ef_8522001a,
        64'h059b06e7_9b634705,
        64'h4107d79b_0107979b,
        64'h8fd90087_979b0644,
        64'h47030654_478308f9,
        64'h1963478d_00f402a3,
        64'hf8000793_c45cc81c,
        64'h57fdee99_e6e30094,
        64'hd49b1ff4_849b0024,
        64'h949bd408_b09ff0ef,
        64'h06040513_f00a93e3,
        64'h10e91163_470dd05c,
        64'h03442023_cc04d458,
        64'h014787bb_24890147,
        64'h073b0909_00b93933,
        64'h19556941_00b67763,
        64'h49051655_6605f326,
        64'h6ce384ae_032655bb,
        64'h40c5063b_f4c563e3,
        64'h873200d7_063b9f3d,
        64'h004ad71b_27810334,
        64'h86bbdfa9_8fd90087,
        64'h979b2501_04244703,
        64'h04344783_14050e63,
        64'h8d5d0085_151b0474,
        64'h47830484_4503ffbd,
        64'h00faf793_01541423,
        64'h00faeab3_008a9a9b,
        64'h04544783_04644a83,
        64'hffc100f9_77b3fff9,
        64'h079b2901_fa0903e3,
        64'h01240123_04144903,
        64'hfaf769e3_0ff7f793,
        64'h009401a3_fff4879b,
        64'h47050134_2e230444,
        64'h44832981_1a098763,
        64'h00f9e9b3_0089999b,
        64'h04a44783_04b44983,
        64'hfee791e3_20000713,
        64'h4107d79b_0107979b,
        64'h8fd90087_979b03f4,
        64'h47030404_4783b785,
        64'h47b5c119_4a01f6e5,
        64'h05e34785_470dbf85,
        64'h00e51963_4785470d,
        64'hfe9915e3_0491c10d,
        64'hea1ff0ef_852285d2,
        64'h000a0763_45090004,
        64'haa030104_8913ff2a,
        64'h14e30991_094100a9,
        64'ha0232501_c51ff0ef,
        64'h854ac789_4501ffc9,
        64'h478389a6_23a40a13,
        64'h1fa40913_848a04f5,
        64'h1a634785_ee5ff0ef,
        64'h85224581_f5718911,
        64'h00090463_fb79478d,
        64'h00157713_092060ef,
        64'h00a400a3_00040023,
        64'h0ff4f513_80826161,
        64'h853e6ae2_7a0279a2,
        64'h794274e2_640660a6,
        64'h47a9c111_89110009,
        64'h0563e385_00157793,
        64'h17e060ef_00144503,
        64'hc79d0004_47830089,
        64'hb023c015_47b184aa,
        64'h638097ba_90c78793,
        64'h0000a797_00351713,
        64'h02054e63_47adddbf,
        64'hf0ef8932_852e89aa,
        64'h00053023_ec56f052,
        64'hfc26e0a2_e486f44e,
        64'hf84a715d_bfcd450d,
        64'h80826105_690264a2,
        64'h644260e2_00a03533,
        64'h8d050125_75332501,
        64'hd25ff0ef_08640513,
        64'h00978c63_45010127,
        64'hf7b31465_04930054,
        64'h4537fff5_09130100,
        64'h05370005_079bd4bf,
        64'hf0ef06a4_051302e7,
        64'h9f63a557_07134107,
        64'hd79b776d_0107979b,
        64'h8fd90087_979b4509,
        64'h23244703_23344783,
        64'he52d2501_fa3ff0ef,
        64'h842ad91c_00050223,
        64'h57fde04a_e426ec06,
        64'he8221101_80826105,
        64'h690264a2_644260e2,
        64'h85220324_a823597d,
        64'h4405c119_25012320,
        64'h60ef0344_8593864a,
        64'h46850014_c503ec19,
        64'h0005041b_fddff0ef,
        64'h892e84aa_02b78763,
        64'h4401e04a_e426ec06,
        64'he8221101_591c8082,
        64'h4501f8df_f06fc399,
        64'h00454783_b7f94505,
        64'hb7e5397d_2aa060ef,
        64'h85ce8626_9cbd4685,
        64'h00144503_4c5cff2a,
        64'h74e34a05_00344903,
        64'h80826145_6a0269a2,
        64'h694264e2_740270a2,
        64'h450100e7_eb6340f4,
        64'h87bb0004_02234c58,
        64'h505ce131_25012ec0,
        64'h60ef85ce_86264685,
        64'h00154503_842a0345,
        64'h0993e052_e84af406,
        64'h5904e44e_ec26f022,
        64'h71798082_853e2781,
        64'h8fd50107_979b8fd1,
        64'h0087179b_0145c603,
        64'h0155c703_00e51d63,
        64'h0006879b_8edd0087,
        64'h979b470d_01a5c683,
        64'h01b5c783_80824525,
        64'h80820141_60a24525,
        64'hc3914501_00157793,
        64'h35e060ef_0017c503,
        64'he4061141_02e69063,
        64'h00855703_0067d683,
        64'hc70d0007_c703cb85,
        64'h611cc915_bfd5b067,
        64'h47030000_a7178082,
        64'h853ae11c_0006871b,
        64'h078900b6_66630ff6,
        64'hf593fd06_869b577d,
        64'h46050007_c683b7dd,
        64'h0705a00d_577d00d7,
        64'h06630017_869300c6,
        64'h986302d5_fc630007,
        64'h468303a0_06130200,
        64'h0593cf99_873e611c,
        64'h80826105_690264a2,
        64'h644260e2_00040023,
        64'h00f49323_8fd90087,
        64'h979b0169_47030179,
        64'h478300f4_92238fd9,
        64'h0087979b_01894703,
        64'h01994783_c088f4bf,
        64'hf0ef00f5_842384ae,
        64'h01c90513_00b94783,
        64'hfcd79be3_07850405,
        64'h00e40023_04050114,
        64'h00230103_15630007,
        64'h831b0e50_071300a7,
        64'h146302c7_00630007,
        64'h470300f9_073346ad,
        64'h02e00893_48214515,
        64'h02000613_47810185,
        64'h3903cfb5_00958413,
        64'he04ae426_ec06e822,
        64'h1101495c_bfc5feb5,
        64'h0fa30505_808200f6,
        64'h13630005_079b9e29,
        64'hb7d500d7_00230785,
        64'h00f50733_00074683,
        64'h00f58733_808200e6,
        64'h13630007_871b4781,
        64'h80822501_8d5d0562,
        64'h8fd907c2_00354503,
        64'h00254783_8f5d07a2,
        64'h00054703_00154783,
        64'h80820141_60a23020,
        64'h00730ff0_000f0000,
        64'h100f7ca0_30efdc65,
        64'h05130000_95173417,
        64'h907307fe_47853007,
        64'h90738fd9_88070713,
        64'h67093000_27f37ee0,
        64'h30efdca5_05130000,
        64'h95177fa0_30efdae5,
        64'h05130000_95178307,
        64'hb58382e7_b823f007,
        64'h07136705_80e7b423,
        64'h8f75e406_16fd1141,
        64'hff8006b7_8087b703,
        64'h300017b7_b7d914fd,
        64'hb7e9bf9f_f0efbfc1,
        64'h710a8493_00a060ef,
        64'h4501dff1_54fd000a,
        64'h2783bfc5_c13ff0ef,
        64'hfc075de3_03379713,
        64'h83093783_02074563,
        64'h03379713_83093783,
        64'h5a0b0493_efbfe0ef,
        64'h8522e78d_0009a783,
        64'he4a9cc07_a1230000,
        64'ha797cc07_a7230000,
        64'ha797cc07_ad230000,
        64'ha797cc07_a9230000,
        64'ha797cc07_9f230000,
        64'ha797d0f7_03a30000,
        64'ha7170054_4783d0f7,
        64'h09230000_a7170044,
        64'h4783d0f7_0ea30000,
        64'ha7170034_4783d2f7,
        64'h04230000_a7173000,
        64'h19370026_2b370024,
        64'h4783d2f7_0da30000,
        64'ha7176a89_d2ca0a13,
        64'h0000aa17_00144783,
        64'hd4f70823_0000a717,
        64'hd3898993_0000a997,
        64'h44810004_4783d5e4,
        64'h04130000_a41710f0,
        64'h30efe925_05130000,
        64'h9517d725_c5830000,
        64'ha597d7b6_46030000,
        64'ha617d846_c6830000,
        64'ha697d8f8_48030000,
        64'ha817d967_c7830000,
        64'ha797d9d7_47030000,
        64'ha71714b0_30efebe5,
        64'h05130000_951780e7,
        64'hb423e05a_e456e852,
        64'hec4ef04a_f426f822,
        64'hfc068f4d_91c115c2,
        64'h00800737_71398087,
        64'hb5838007_b6033000,
        64'h17b78082_61616ae2,
        64'h7a0279a2_794274e2,
        64'h82f6b423_47a16406,
        64'h60a68086_b7838006,
        64'hb78380f6_b42393c1,
        64'h80a6b023_17c29101,
        64'h300016b7_8fd91502,
        64'h0ff77713_8ff18321,
        64'h0087179b_f0060613,
        64'h01000637_4722f43f,
        64'hf0ef4512_043050ef,
        64'h0028e325_85930000,
        64'ha5974609_053050ef,
        64'h0048e445_85930000,
        64'ha5974611_fc941ee3,
        64'h1f9030ef_00c78023,
        64'h0ff67613_00ca5633,
        64'h0286061b_0405854a,
        64'h0004059b_013407b3,
        64'h028a863b_4499f769,
        64'h09130000_9917e7e9,
        64'h89930000_a9975ae1,
        64'h44012330_30eff7e5,
        64'h05130000_95178a2a,
        64'h017070ef_c63eec56,
        64'hf052f44e_f84afc26,
        64'he0a2e486_04b00513,
        64'h45854601_00740207,
        64'h879b0700_07b7715d,
        64'h80822501_8d5d8d79,
        64'h00ff0737_0085151b,
        64'h8fd98f75_0085571b,
        64'hf0068693_8fd966c1,
        64'h0185579b_0185171b,
        64'h80829141_15428d5d,
        64'h05220085_579b8082,
        64'h614564e2_740270a2,
        64'h85228b8f_f0eff065,
        64'h05130000_a5170450,
        64'h0693efe7_57030000,
        64'ha717efa8_88930000,
        64'ha89785a6_862247b2,
        64'h0007a803_f1478793,
        64'h0000a797_14b050ef,
        64'hf4060068_f5c58593,
        64'h0000a597_461184ae,
        64'h8432ec26_f0227179,
        64'hbfc14785_ec3ff0ef,
        64'h80826105_64a26442,
        64'h60e2c3c0_0c2007b7,
        64'h311030ef_04450513,
        64'h00009517_e7990206,
        64'hc1630337_16938304,
        64'hb7033000_14b74781,
        64'h2401ec06_e42643c0,
        64'he8220c20_07b71101,
        64'h80826101_01135f81,
        64'h34838526_60013403,
        64'h60813083_8287b823,
        64'h300017b7_0405a9bf,
        64'hf0ef8626_fef845e3,
        64'h0006881b_ff063c23,
        64'h06210685_00083803,
        64'h983a0036_98139742,
        64'h85b24681_4037d79b,
        64'h30000837_860a2785,
        64'h0077e793_37ed02d5,
        64'h1e638066_86936685,
        64'hc6918005_069b0001,
        64'h550300d1_00230086,
        64'hd69b0106_d69b0106,
        64'h969b00d1_00a345d4,
        64'h95ba070e_9f318006,
        64'h871b7007_76130084,
        64'h171beb3d_43180267,
        64'h07130000_a717c349,
        64'h27018f71_fff74713,
        64'h00c5163b_10100513,
        64'h8a1d0905_6c63ffc7,
        64'h849b5f20_0513fee7,
        64'h881b2781_60113423,
        64'h5e913c23_639c97ae,
        64'h300005b7_9fad8406,
        64'h879b0387_f5930034,
        64'h179b6685_8387b703,
        64'h00f67413_26016081,
        64'h30239f01_01138307,
        64'hb6033000_17b7bba5,
        64'h46014430_30ef15e5,
        64'h05130000_951785aa,
        64'hb36900f4_16236080,
        64'h079300f4_1f230024,
        64'hd78300f4_1e230004,
        64'hd78302f4_142301e4,
        64'h578302f4_132302a0,
        64'h061301c4_57832ed0,
        64'h50ef8522_85ca4619,
        64'h2f7050ef_00640513,
        64'h0f058593_0000a597,
        64'h46193090_50ef854e,
        64'h10058593_0000a597,
        64'h46193190_50ef854a,
        64'h85ce4619_00f59a23,
        64'h01658993_02058913,
        64'h20000793_eaf719e3,
        64'h1427d783_0000a797,
        64'h0285d703_ecf711e3,
        64'h15048493_0000a497,
        64'h1587d783_0000a797,
        64'h0265d703_b1e91d65,
        64'h05130000_9517b9d1,
        64'h1c850513_00009517,
        64'hb9f91a25_05130000,
        64'h9517b1e5_18c50513,
        64'h00009517_b9cd17e5,
        64'h05130000_9517b9f5,
        64'h16050513_00009517,
        64'hb31915a5_05130000,
        64'h9517bb01_14450513,
        64'h00009517_bb291365,
        64'h05130000_9517b315,
        64'h12050513_00009517,
        64'hb33d11a5_05130000,
        64'h9517b799_3cb050ef,
        64'h08681da5_85930000,
        64'ha5974611_f4f70de3,
        64'h02045703_f6f701e3,
        64'h17fd67c1_01e45703,
        64'hf6e787e3_5fe00713,
        64'hbf95c8cf_f0ef02a4,
        64'h051385ca_595030ef,
        64'h14050513_00009517,
        64'hca2ff0ef_852285a6,
        64'h5a9030ef_14450513,
        64'h00009517_02e79863,
        64'h4d200713_b765d4bf,
        64'he0ef02a4_051321e5,
        64'h85930000_a59721a6,
        64'h06130000_a61721e6,
        64'h86930000_a697f7e9,
        64'h439c22a7_87930000,
        64'ha797c799_439c23a7,
        64'h87930000_a79722f7,
        64'h2b230000_a71747e2,
        64'h04e69463_04300713,
        64'h80826161_79a27942,
        64'h74e26406_60a65900,
        64'h60ef4501_02a40593,
        64'hff89061b_24c78793,
        64'h0000a797_66a24762,
        64'h49f050ef_e43626f7,
        64'h2b230000_a7172765,
        64'h05130000_a51726e5,
        64'h85930000_a5974619,
        64'h47e228d7_9b230000,
        64'ha79704e7_9b6301c1,
        64'h56830450_071300e1,
        64'h0e230234_470300e1,
        64'h0ea301c1_19030224,
        64'h470300e1_0e232781,
        64'h02744703_00e10ea3,
        64'h01c11783_00f10e23,
        64'h02544783_00f10ea3,
        64'h02644703_02444783,
        64'hbdbd22a5_05130000,
        64'h9517b561_21c50513,
        64'h00009517_bd4920e5,
        64'h05130000_9517a06d,
        64'hda5fe0ef_450185a2,
        64'h862602a4_122300a1,
        64'h1e238d5d_05220085,
        64'h579bdb3f_f0ef00f4,
        64'h1e230029_d78300f4,
        64'h1d230009_d78302f4,
        64'h10230224_0513fde4,
        64'h859b01c4_578300f4,
        64'h1f230204_12230204,
        64'h012301a4_578357d0,
        64'h50ef854a_37458593,
        64'h0000a597_461958d0,
        64'h50ef8522_85ca4619,
        64'h10f71b63_3a67d783,
        64'h0000a797_02045703,
        64'h12f71363_3b498993,
        64'h0000a997_3bc7d783,
        64'h0000a797_01e45703,
        64'hb73d40a5_05130000,
        64'h9517f0f5_9ce30880,
        64'h079326f5_88630ff0,
        64'h079326f5_87630890,
        64'h0793b73d_f4f58ae3,
        64'h40050513_00009517,
        64'h06c00793_26f58a63,
        64'h06700793_00b7ef63,
        64'h28f58563_08400793,
        64'hbf91f6f5_8de33ee5,
        64'h05130000_951705e0,
        64'h079328f5_836305c0,
        64'h0793b7bd_f8f58ae3,
        64'h3d850513_00009517,
        64'h03200793_28f58663,
        64'h02f00793_00b7ef63,
        64'h2af58163_03300793,
        64'h04b7e263_2cf58163,
        64'h06200793_b7c93d65,
        64'h05130000_9517faf5,
        64'h96e30290_07932af5,
        64'h85630210_0793bf6d,
        64'hfef580e3_3bc50513,
        64'h00009517_47d916f5,
        64'h896347c5_00b7ed63,
        64'h2cf58163_47f5a429,
        64'h020040ef_fef591e3,
        64'h3a050513_00009517,
        64'h47a118f5_81634799,
        64'ha41503a0_40ef5365,
        64'h05130000_951702f5,
        64'h836339a5_05130000,
        64'h95174789_10f58463,
        64'h478502b7_e3631af5,
        64'h82634791_04b7e563,
        64'h1cf58163_47b108b7,
        64'he76332f5_886302e0,
        64'h07930174_45836ed0,
        64'h50ef4aa5_05130000,
        64'ha5174619_85ca0064,
        64'h09137010_50ef4611,
        64'h082884b2_05e94407,
        64'h99638005_079b0af5,
        64'h0e636dd7_879367a1,
        64'h3cf50463_842e8067,
        64'h8793f44e_f84afc26,
        64'he486e0a2_6785715d,
        64'hbf45943e_93c117c2,
        64'h00f11723_8fd90087,
        64'h979b0087_d71b0489,
        64'h00c15783_753050ef,
        64'h00684609_85a68082,
        64'h61459141_694264e2,
        64'h1542fff5_45137402,
        64'h70a29522_01045513,
        64'h942a9041_14420104,
        64'h551302f0_44634099,
        64'h07bb00a5_893b4401,
        64'h84aaf406_e84aec26,
        64'hf0227179_80824165,
        64'h05130000_9517bf75,
        64'h46050513_00009517,
        64'h84078793_fce608e3,
        64'h46050513_00009517,
        64'h83878713_bfe944e5,
        64'h05130000_95178287,
        64'h879300c7_4963fee6,
        64'h09e34725_05130000,
        64'h95178307_87138082,
        64'hfaf612e3_45450513,
        64'h00009517_81878793,
        64'h00e60a63_45450513,
        64'h00009517_81078713,
        64'h80820141_5ac50513,
        64'h0000a517_60a21820,
        64'h40efe406_5bc50513,
        64'h0000a517_4f458593,
        64'h00009597_9e3d1141,
        64'h7c07879b_77fd04c7,
        64'hc9635025_05130000,
        64'h951787f7_87936785,
        64'hc3ad4825_05130000,
        64'h95178006_079b04c7,
        64'h496306e6_0b634a65,
        64'h05130000_95178087,
        64'h871308a7_4463862a,
        64'h0ce50763_82078713,
        64'h67858082_953e057e,
        64'h450597aa_20000537,
        64'he3089536_00178693,
        64'h00756513_157d631c,
        64'h65870713_0000a717,
        64'h80824000_05378082,
        64'h057e4505_8082853e,
        64'h4785bf99_03840413,
        64'h2a0506a0_60ef856a,
        64'h4581864e_254040ef,
        64'h856285ea_9d3e864e,
        64'h40f989b3_01843d03,
        64'h0337f163_701c0284,
        64'h39830e00_60ef856a,
        64'h85ee864e_27c040ef,
        64'h856686ce_85ea866e,
        64'h80826165_853e6da2,
        64'h6d426ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h694664e6_740670a6,
        64'h478d2aa0_40ef5065,
        64'h05130000_9517864a,
        64'h02bafa63_95ce00b4,
        64'h8db30184_3d03640c,
        64'h04098d63_02043983,
        64'h2d0040ef_855e85d2,
        64'hcbc1741c_09679b63,
        64'h401ca835_478100fa,
        64'h64630384_d783566c,
        64'h8c930000_9c97586c,
        64'h0c130000_9c17546b,
        64'h8b930000_9b974b05,
        64'h4a01942a_84aa892e,
        64'h06eae663_478d9722,
        64'h020ada93_e46ee86a,
        64'hec66f062_f45ef85a,
        64'he0d2e4ce_e8caeca6,
        64'hf4860205_9a93fc56,
        64'h7100f0a2_02f70733,
        64'h71590380_07930385,
        64'h570310e6_97634709,
        64'h00454683_10e69c63,
        64'h478957f7_0713464c,
        64'h47370005_668312b7,
        64'hf4630400_0793bfd5,
        64'h8f8d2505_8082e21c,
        64'h00b7f463_45019181,
        64'h87aa1582_b70d0705,
        64'h27850117_00230006,
        64'h54634186_561b0186,
        64'h161bc519_09757513,
        64'h00054503_00cc0533,
        64'h00074603_bfdd4781,
        64'hbf253cfd_fe97eae3,
        64'h27856782_0dc070ef,
        64'he03e855e_b76500c5,
        64'h80230ff6_761395be,
        64'h082c0007_4603bf6d,
        64'h00c59023_95aa9241,
        64'h16420828_00179593,
        64'h00075603_011d1d63,
        64'hbfd1e190_95aa0828,
        64'h00379593_6310010d,
        64'h1963bf9d_46914821,
        64'h07859752_488967a2,
        64'h67024120_40efe03a,
        64'he43e855a_85d69201,
        64'h1602c190_95aa2601,
        64'h08280027_95934310,
        64'h02dd1963_b79d557d,
        64'hd13d0b00_70ef9936,
        64'h92811682_41b4043b,
        64'h668244a0_40effa07,
        64'h8c23e036_69450513,
        64'h00009517_97ba1098,
        64'h0b079c63_0006881b,
        64'h02e00893_85ba4781,
        64'h083803bd_06bb0d9d,
        64'he56399be_034787b3,
        64'h9381020d_979305b6,
        64'h6b630007_861b4889,
        64'h48214691_4781874e,
        64'h000c8d9b_008cf463,
        64'h00040d9b_4a4040ef,
        64'h6d850513_00009517,
        64'h85ca8082_61697da6,
        64'h7d467ce6_6c0a6baa,
        64'h6b4a6aea_7a0a79aa,
        64'h794a74ea_640e60ae,
        64'h4501e00d_5dcc0c13,
        64'h00008c17_684b8b93,
        64'h00009b97_71cb0b13,
        64'h00009b17_020a5a13,
        64'h001a849b_020d1a13,
        64'h001d1a9b_03acdcbb,
        64'h4cc1000c_956302cc,
        64'hdcbb0400_0c9300e7,
        64'hf6638436_8d3289ae,
        64'h892a0400_0793f4ee,
        64'he162e55e_e95aed56,
        64'hf152fd26_e586f8ea,
        64'hf54ef94a_e1a202c7,
        64'h073b8cba_fce67155,
        64'h5400406f_610576e5,
        64'h05130000_951764a2,
        64'h690285a6_864a60e2,
        64'h644255a0_40ef7665,
        64'h05130000_951785a2,
        64'hc80156a0_40ef8932,
        64'h77050513_00009517,
        64'h85be0785_14590087,
        64'h74630104_5433942a,
        64'h472500d4_14334405,
        64'h03b6869b_02e50533,
        64'h4729c10d_44018d79,
        64'hfff74713_01071733,
        64'h577db7f5_7c450513,
        64'h00009517_85aafab7,
        64'h1ce32705_5bc0406f,
        64'h61057da5_05130000,
        64'h951785aa_690264a2,
        64'h60e26442_e495e04a,
        64'he822ec06_00074483,
        64'he426972e_11017ce5,
        64'h85930000_a5979301,
        64'h1702cf85_00f557b3,
        64'h883e03c6_879b02e8,
        64'h86bb4599_58d94701,
        64'h862ebfa1_7fc50513,
        64'h00009517_85aabf55,
        64'h4401bf51_843a0086,
        64'hf46302f4_5733bf61,
        64'h02e45433_62c0406f,
        64'h61058425_05130000,
        64'ha5176902_64a285ca,
        64'h862660e2_64426460,
        64'h40ef8525_05130000,
        64'ha51785a2_c8016560,
        64'h40ef84b2_85c50513,
        64'h0000a517_943e0014,
        64'h44130324_341302e4,
        64'h743302f4_57b30640,
        64'h07130087_7d630630,
        64'h0713cf39_02f47733,
        64'h46a547a9_0687e263,
        64'h47293e80_0793c815,
        64'h02f555b3_02f57433,
        64'hbf7d2407_87934685,
        64'hb7d9a007_87934681,
        64'h6b00406f_61058a65,
        64'h05130000_a51785aa,
        64'h690264a2_60e26442,
        64'h02091663_e426e822,
        64'hec060007_4903e04a,
        64'h97361101_8cc70713,
        64'h0000b717_3e800793,
        64'h46890ca7_fc633e70,
        64'h079304a7_676323f7,
        64'h8713000f_47b704a7,
        64'h6963862e_9ff78713,
        64'h3b9ad7b7_8082612d,
        64'h450160ee_714040ef,
        64'h90050513_0000a517,
        64'h002cfebf_f0efed86,
        64'h45050c80_0613002c,
        64'h7115f73f_f06f4581,
        64'h862e86b2_80826145,
        64'h69a26942_64e2854a,
        64'h740270a2_306060ef,
        64'h91858593_0000a597,
        64'h00890533_ffd4841b,
        64'h00f44463_ffe4879b,
        64'h9c2972a0_40ef954a,
        64'h94860613_0000a617,
        64'h86ce40a4_85bb0095,
        64'h5d630009_8f63842a,
        64'h748040ef_854a85a6,
        64'h96060613_0000a617,
        64'he1870713_00009717,
        64'h96868693_0000a697,
        64'hc5092226_86930000,
        64'ha6978932_89ae84b6,
        64'hf022f406_e44ee84a,
        64'hec267179_bfdd7c60,
        64'h40ef8562_b7f10905,
        64'h7d0040ef_856600fb,
        64'he7630ff7_f793fe05,
        64'h879b0007_c5830129,
        64'h87b3bf15_04857ee0,
        64'h40ef50a5_05130000,
        64'ha51700f4_5a630009,
        64'h079b4124_093b0070,
        64'h40ef00f4_f913855a,
        64'hff2dcce3_2d850170,
        64'h40ef8552_bfdd01f0,
        64'h40ef8562_b75d0905,
        64'h029040ef_856600fb,
        64'he7630ff7_f793fe05,
        64'h879b0007_c5830129,
        64'h87b3a805_00f97913,
        64'h4d81fffd_4913068d,
        64'h12630530_40efa165,
        64'h05130000_a5170007,
        64'hc5830099_87b30670,
        64'h40ef8552_06d040ef,
        64'h58850513_0000a517,
        64'h02879d63_0009079b,
        64'hff048913_085040ef,
        64'h855ae39d_00f47793,
        64'hc01d8082_61656da2,
        64'h6d426ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h694664e6_740670a6,
        64'h03544163_0004841b,
        64'hfff58d1b_a6cc8c93,
        64'h0000ac97_a7cc0c13,
        64'h0000ac17_06000b93,
        64'ha70b0b13_0000ab17,
        64'h7a0a0a13_0000aa17,
        64'h44818aae_89aae46e,
        64'he8caf0a2_f486e86a,
        64'hec66f062_f45ef85a,
        64'hfc56e0d2_e4ceeca6,
        64'h7159b7cd_105040ef,
        64'hd007a823_0000b797,
        64'ha9850513_0000a517,
        64'h80826151_641260b2,
        64'h85221230_40efa7e5,
        64'h05130000_a517a565,
        64'h85930000_a597860a,
        64'hc10d842a_e01ff0ef,
        64'h85221430_40efa765,
        64'h05130000_a517a765,
        64'h85930000_a597842a,
        64'h00054603_00154683,
        64'h00254703_00354783,
        64'h00454803_00554883,
        64'he222e606_716d8082,
        64'h616569a6_694664e6,
        64'h74064501_70a67f01,
        64'h01138ddf_f0ef86c6,
        64'h85a61808_56326882,
        64'hfc4ff0ef_03e10513,
        64'h863e86c2_85a267c2,
        64'h6822f94f_f0efd64e,
        64'h05210513_85a2864a,
        64'h86ba943e_7fc40413,
        64'h6762747d_97ba8107,
        64'h87931018_678503d0,
        64'h60efd602_e83eec3a,
        64'he4428936_89b2e046,
        64'h05a10513_84aa8101,
        64'h0113e4ce_e8caeca6,
        64'hf0a2f486_71591f70,
        64'h406fb125_05130000,
        64'ha51785aa_80826125,
        64'h7aa27a42_79e26906,
        64'h64a66446_450160e6,
        64'h911a6305_96fff0ef,
        64'h85ce86a6_10084652,
        64'h855ff0ef_460156fd,
        64'h02e10513_85a2821f,
        64'hf0ef0440_06130430,
        64'h06930421_051385a2,
        64'h943e1451_978a020a,
        64'h879312f1_1c233537,
        64'h87936799_12f11b23,
        64'h26378793_77e10d50,
        64'h60ef04f1_06230661,
        64'h05134641_479985ce,
        64'h04f11523_10100793,
        64'h0a1060ef_ca3e04a1,
        64'h05134581_0f000613,
        64'h0fc00793_103060ef,
        64'h000107a3_15410223,
        64'h14f101a3_14510513,
        64'h460585ca_57fd11d0,
        64'h60ef13f1_05134611,
        64'h95beff04_0593978a,
        64'h020a8793_12f10f23,
        64'h479112f1_0ea30370,
        64'h07931410_60ef0141,
        64'h07a31a68_460585ca,
        64'h993e978a_020a8793,
        64'h12f11d23_13500793,
        64'hc83e4a05_fef40913,
        64'h439ccda7_87930000,
        64'hb7971230_60ef8526,
        64'h55fd4619_94beff84,
        64'h0493978a_020a8793,
        64'h747d31b0_40efca02,
        64'h6a85c225_05130000,
        64'ha517911a_89aaf456,
        64'hf852fc4e_e0cae4a6,
        64'he8a2ec86_711d737d,
        64'hb34d3430_40efc0e5,
        64'h05130000_a517bf45,
        64'hc0850513_0000a517,
        64'h95be978a_d0040593,
        64'h35078793_67853670,
        64'h40efc025_05130000,
        64'ha5173730_40efbfe5,
        64'h05130000_a51700fa,
        64'h20234785_de0794e3,
        64'h000a2783_b3fd38f0,
        64'h40efc0a5_05130000,
        64'ha517bbf5_39d040ef,
        64'hc0050513_0000a517,
        64'h95be978a_f0040593,
        64'h35048793_3b5040ef,
        64'hc0850513_0000a517,
        64'h95bee004_0593978a,
        64'h35048793_3cd040ef,
        64'h02f5d5bb_e107879b,
        64'h678502f6_763b02f5,
        64'hf6bb02f5_d63b03c0,
        64'h079304f7_1e230000,
        64'hb7170121_578306f7,
        64'h13230000_b717c2e5,
        64'h05130000_a51755c2,
        64'h01015783_40d040ef,
        64'hc2050513_0000a517,
        64'h01014583_01114603,
        64'h01214683_01314703,
        64'h429040ef_c1c50513,
        64'h0000a517_01814583,
        64'h01914603_01a14683,
        64'h01b14703_445040ef,
        64'h00b14703_0cf71323,
        64'h0000b717_c1c50513,
        64'h0000a517_00814583,
        64'h35215783_0cf71e23,
        64'h0000b717_00914603,
        64'h00a14683_35015783,
        64'h479040ef_c1c50513,
        64'h0000a517_35014583,
        64'h35114603_35214683,
        64'h35314703_303060ef,
        64'h01490593_4611953e,
        64'hcb840513_978a3504,
        64'h87936485_31b060ef,
        64'h0e880109_05934611,
        64'h4b9040ef_c4c50513,
        64'h0000a517_00fa2023,
        64'h47851207_9a63000a,
        64'h2783b321_d00d0023,
        64'h347060ef_9d228562,
        64'h866ab749_cc048513,
        64'hbb39cef4_2023401c,
        64'h00f41023_8fd90087,
        64'h979b0087_d71bce24,
        64'h578300f4_11238fd9,
        64'h0087979b_0087d71b,
        64'hce045783_383060ef,
        64'h4611953e_ce048513,
        64'h978a3507_87936785,
        64'hbfdd855a_4611b395,
        64'h39f060ef_85564611,
        64'hb3bdf00d_00233ad0,
        64'h60ef9d22_953e866a,
        64'hf0048513_978a3507,
        64'h87936785_a00d953e,
        64'h978a3507_87936785,
        64'h4611cd04_85138082,
        64'h3b010113_35013d03,
        64'h35813c83_36013c03,
        64'h36813b83_37013b03,
        64'h37813a83_38013a03,
        64'h38813983_39013903,
        64'h39813483_3a013403,
        64'h3a813083_911a6305,
        64'hcf3ff0ef_0e8885de,
        64'h86ca5672_bd9ff0ef,
        64'h35e10513_85a24601,
        64'h56fdba5f_f0ef3721,
        64'h051385a2_04400613,
        64'h04300693_943ecec4,
        64'h0413978a_350a8793,
        64'h46f11423_35378793,
        64'h679946f1_13232637,
        64'h879377e1_45b060ef,
        64'h36f10e23_39610513,
        64'h85de4799_464136f1,
        64'h1d231010_07934270,
        64'h60efde3e_37a10513,
        64'h45810f00_06131020,
        64'h07934890_60ef4731,
        64'h0d230001_03a346f1,
        64'h0ca347b1_051385a6,
        64'h460557fd_4a3060ef,
        64'h47410a23_47510513,
        64'h461195be_cf440593,
        64'h978a350a_879346f1,
        64'h09a30360_07934c50,
        64'h60ef4741_072346f1,
        64'h05134611_4a1195be,
        64'hcf040593_978a350a,
        64'h879346f1_06a30320,
        64'h07934e90_60efc0d2,
        64'h46c10513_85a64605,
        64'h94becb74_0493c2a6,
        64'h978a350a_879346f1,
        64'h15231350_079300f1,
        64'h03a3478d_4c5060ef,
        64'h854a55fd_4619993e,
        64'hcf840913_978a350a,
        64'h87936bb0_40efde02,
        64'h54e25a52_e3c50513,
        64'h0000a517_53b060ef,
        64'h953e4611_01490593,
        64'hce840513_978a350a,
        64'h87935510_60ef013c,
        64'ha023953e_46110109,
        64'h0593ce44_05134985,
        64'h978a350a_87936a85,
        64'h16079263_000ca783,
        64'h3af59f63_478938f5,
        64'h83634799_24f58363,
        64'h747d4795_00614583,
        64'hf8e79ce3_0ff00713,
        64'h24e78563_03800713,
        64'haac94605_cb648513,
        64'hfae798e3_03500713,
        64'h20e78e63_03300713,
        64'h00f76e63_22e78163,
        64'h03600713_b769e00d,
        64'h00235c90_60ef9d22,
        64'h953e866a_e0048513,
        64'h978a3507_87936785,
        64'hfee794e3_473d22e7,
        64'h83634731_bf4d77f0,
        64'h40ef0625_05130000,
        64'ha51785be_22e78763,
        64'hcc848513_470d2ae7,
        64'h89634705_02f76263,
        64'h22e78f63_471904f7,
        64'h6b6326e7_8b6301a9,
        64'h89bb0589_02a00713,
        64'h29890f07_c7830015,
        64'hcd030139_07b395ca,
        64'h0f098593_9c3a9b3a,
        64'h49818a36_8cb28bae,
        64'hd0048c13_cb848b13,
        64'h970a3507_87139aba,
        64'hcd848a93_970a3507,
        64'h871374fd_678524f7,
        64'h1d634789_00054703,
        64'ha0010020_50eff5e5,
        64'h05130000_a51785aa,
        64'h00e7ea63_892a5800,
        64'h073797aa_d0040023,
        64'hf0040023_e0040023,
        64'hca040b23_ce042023,
        64'hd00007b7_943e747d,
        64'h978a911a_35078793,
        64'h35a13823_35913c23,
        64'h37813023_37713423,
        64'h37613823_37513c23,
        64'h39413023_39313423,
        64'h38913c23_3a113423,
        64'h39213823_3a813023,
        64'h6785737d_c5010113,
        64'hfadff06f_614564e2,
        64'h00e4859b_70a27402,
        64'h852200f4_162347a1,
        64'h6ff060ef_85b64619,
        64'h852266a2_70b060ef,
        64'he436f406_46190519,
        64'h84b2842a_ec26f022,
        64'h71798082_01416402,
        64'h60a28522_fa1ff0ef,
        64'he4064501_85aa8622,
        64'h0005841b_e0221141,
        64'hbfe10505_01173023,
        64'h97369742_0008b883,
        64'h00e588b3_00351713,
        64'h808280c6_b82396be,
        64'h678500f7_47630005,
        64'h071b6805_450102e7,
        64'hc7bb2785_0077e793,
        64'hfff6079b_8007bc23,
        64'h97b64721_67856394,
        64'h31078793_0000b797,
        64'h80826145_740270a2,
        64'h00f41523_fff7c793,
        64'h9fb94107_d71b9fb9,
        64'h93411742_4107579b,
        64'hfed79ce3_9f31ffe7,
        64'hd6030789_470187a2,
        64'h01440693_7c3060ef,
        64'h01040513_002c4611,
        64'h7cf060ef_00c40513,
        64'h00041523_006c4611,
        64'h00f404a3_47c57e50,
        64'h60efec3e_00840513,
        64'h00041323_082c4621,
        64'h47c17f90_60ef0044,
        64'h05130161_05934609,
        64'h006070ef_00f11b23,
        64'hc4360509_084c57fd,
        64'h460900f1_1a238fd9,
        64'h0087979b_0ff77713,
        64'h0087d713_c632842a,
        64'h419c00f5_10230457,
        64'h879b6785_c19c27d1,
        64'hf022f406_7179419c,
        64'h80820005_132300f5,
        64'h122300d5_112300c5,
        64'h10238fd9_0087979b,
        64'h0ff77713_c19c0087,
        64'hd7138ed9_06a20086,
        64'hd71b8e59_27a10622,
        64'h0086571b_419cc19c,
        64'h2785c319_0017f713,
        64'h419cbfcd_fda00513,
        64'h80826121_74a27442,
        64'h70e29782_85a66562,
        64'h701ce509_c39ff0ef,
        64'h842a0830_65a2c105,
        64'hc7dff0ef_84b2e42e,
        64'hf822fc06_f4267139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2655c,
        64'h862686ca_6562e519,
        64'hc75ff0ef_083065a2,
        64'hc115cb7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2615c,
        64'h862686ca_6562e519,
        64'hcb5ff0ef_083065a2,
        64'hc115cf7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hb7e16522_f569cdbf,
        64'hf0ef8526_85ce0030,
        64'hbfc90284_8493c501,
        64'h71d060ef_854a608c,
        64'h2f0050ef_855285ca,
        64'h60908082_61216a42,
        64'h69e27902_74a27442,
        64'h70e24501_00849b63,
        64'h942602f4_043325ea,
        64'h0a130000_aa1789ae,
        64'h892afc06_e852ec4e,
        64'hf04a0280_079302f4,
        64'h043b840d_8c0564e4,
        64'h84930000_b4976564,
        64'h04130000_b417f426,
        64'hf822639c_4f478793,
        64'h0000b797_7139bfdd,
        64'h45018082_61056442,
        64'h60e2fda0_05138302,
        64'h610560e2_65a26442,
        64'h85220003_0e630205,
        64'h3303c919_db9ff0ef,
        64'he42eec06_4108842a,
        64'he8221101_bfc56562,
        64'hf96dd97f_f0ef0830,
        64'h80826145_70a24501,
        64'he50965a2_de1ff0ef,
        64'hf406e42e_7179bfc1,
        64'h5479fcf7_1be30ff0,
        64'h079300c7_c70367a2,
        64'h0d6080ef_6522f565,
        64'h842adcff_f0ef85a6,
        64'h00308522_80826145,
        64'h64e27402_70a28522,
        64'h54351020_80ef31e5,
        64'h05130000_a51700f4,
        64'hcf63445c_3f4050ef,
        64'h32050513_0000a517,
        64'h85a6842a_c11dfda0,
        64'h0413e47f_f0ef84ae,
        64'hf406ec26_f0227179,
        64'h80826145_694264e2,
        64'h740270a2_852213c0,
        64'h80ef6522_42c050ef,
        64'h34850513_0000a517,
        64'h864a608c_ed01842a,
        64'he45ff0ef_84aa85ca,
        64'h0030c11d_fda00413,
        64'he8dff0ef_892eec26,
        64'hf406e84a_f0227179,
        64'hb7d92405_17a080ef,
        64'h652246a0_50ef854e,
        64'h85a20127_896300c7,
        64'hc78367a2_ed09e83f,
        64'hf0ef8526_85a20030,
        64'h80826121_69e27902,
        64'h74a27442_70e200f4,
        64'h496344dc_3a498993,
        64'h0000a997_0ff00913,
        64'h440184aa_cd01eebf,
        64'hf0efec4e_f04af426,
        64'hf822fc06_7139bfd5,
        64'h54798082_61457402,
        64'h70a28522_1e0080ef,
        64'h00f70963_00c54703,
        64'h0ff00793_6562e911,
        64'h842aee7f_f0ef0830,
        64'h65a2c105_fda00413,
        64'hf2dff0ef_e42ef406,
        64'hf0227179_b7c1fda0,
        64'h0513bf65_240521a0,
        64'h80ef4981_652250e0,
        64'h50ef8552_00099563,
        64'h2485cb99_0087c783,
        64'h67a2ed19_f29ff0ef,
        64'h854a85a2_00308082,
        64'h61216a42_69e27902,
        64'h74a27442_70e25535,
        64'he0914501_00f44d63,
        64'h00c92783_264a0a13,
        64'h0000ba17_44014481,
        64'h4985892a_cd31f9bf,
        64'hf0efe852_ec4ef04a,
        64'hf426f822_fc067139,
        64'hbfe54501_80820141,
        64'h60a26108_c509fbbf,
        64'hf0efe406_1141b7f5,
        64'h02870713_fea68de3,
        64'h47148082_853a4701,
        64'h00e79563_97ba02d7,
        64'h87b30280_069302d7,
        64'h87bb878d_8f998c67,
        64'h87930000_c7976294,
        64'h8d070713_0000c717,
        64'h76868693_0000b697,
        64'hb7edfda0_07138302,
        64'h853e85b2_00030563,
        64'h01853303_8082853a,
        64'he21c97b6_470102a7,
        64'h87b30a00_051300b7,
        64'hd963454c_0005cc63,
        64'h5735c285_87ae6914,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h000a2e2e_2e746e65,
        64'h6d6f6d20_61207469,
        64'h61772065_7361656c,
        64'h50202165_6e616972,
        64'h41206d6f_7266206f,
        64'h6c6c6548_ffdff06f,
        64'h10500073_34102373,
        64'h342022f3_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_65a090ef,
        64'hfec5c6e3_02058593,
        64'h0005bc23_0005b823,
        64'h0005b423_0005b023,
        64'h09060613_0000c617,
        64'hb3058593_0000c597,
        64'h30579073_09078793,
        64'h00000797_00078067,
        64'h40b787b3_00d787b3,
        64'h01478793_00000797,
        64'hfcc5cce3_02068693,
        64'h02058593_00e6bc23,
        64'h0185b703_00e6b823,
        64'h0105b703_00e6b423,
        64'h0085b703_00e6b023,
        64'h0005b703_0006b703,
        64'hff810113_01b11113,
        64'h0110011b_fe0e9ae3,
        64'h0085b703_fffe8e93,
        64'h0005b703_240e8e9b,
        64'h000f4eb7_01169693,
        64'hfff6869b_000066b7,
        64'hac560613_0000c617,
        64'hfc058593_00000597,
        64'h000280e7_13050513,
        64'h00000517_11c28293,
        64'h00008297_000280e7,
        64'h0f628293_00008297,
        64'h01111113_fff1011b,
        64'h00006137_11249463,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
