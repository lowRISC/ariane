/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module etherboot (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 6023;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_87fe7094,
        64'h00000000_87fe70d2,
        64'h00000000_00000000,
        64'hffffffff_00000006,
        64'h00000000_87feb5c0,
        64'h00000000_2f7c5c2d,
        64'h00000000_ffffffff,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_cc33aa55,
        64'h00000000_87feb408,
        64'h00006772_615f6473,
        64'h0000646d_635f6473,
        64'h00000000_0c000000,
        64'h00000000_ffffffff,
        64'h00000000_00000000,
        64'h00000000_43000000,
        64'h00000000_004b4d47,
        64'h00004b4d_47545045,
        64'h00000003_0f060301,
        64'haaaaaaaa_aaaaaaaa,
        64'h55555555_55555555,
        64'h5851f42d_4c957f2d,
        64'h10000000_20000000,
        64'h10325476_98badcfe,
        64'hefcdab89_67452301,
        64'h00000002_464c457f,
        64'hcccccccc_cccccccd,
        64'h00000a0d_70617274,
        64'h00000000_000a7473,
        64'h65742065_68636143,
        64'h00000000_00000a74,
        64'h6f6f6220_50544654,
        64'h00000000_00000a74,
        64'h73657420_4d415244,
        64'h00000000_00000a74,
        64'h6f6f6220_49505351,
        64'h00000000_00000000,
        64'h0a746f6f_62204453,
        64'h00000000_0000000a,
        64'h5825203d_20646565,
        64'h73206d6f_646e6152,
        64'h000a5825_2c582520,
        64'h3d20676e_69747465,
        64'h73206863_74697753,
        64'h0000000a_5825203d,
        64'h205d6425_5b707773,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h0a646c25_2e646c25,
        64'h203d2049_5043202c,
        64'h73656c63_79632064,
        64'h6c25202c_736e6f69,
        64'h74637572_74736e69,
        64'h20646c25_202c424b,
        64'h6425203d_20746573,
        64'h5f676e69_6b726f77,
        64'h00000000_00000000,
        64'h0a2e2979_6c6e6f28,
        64'h2032206e_6f697372,
        64'h65762065_736e6563,
        64'h694c2063_696c6275,
        64'h50206c61_72656e65,
        64'h4720554e_47206568,
        64'h74207265_646e7520,
        64'h6465736e_6563694c,
        64'h00000000_0000000a,
        64'h2e6e6f62_617a6143,
        64'h2073656c_72616843,
        64'h20323130_322d3130,
        64'h30322029_43282074,
        64'h68676972_79706f43,
        64'h00000000_0000000a,
        64'h29746962_2d642528,
        64'h20302e33_2e34206e,
        64'h6f697372_65762072,
        64'h65747365_746d656d,
        64'h00000a74_73657420,
        64'h4d415244_206c6174,
        64'h656d2065_7261420a,
        64'h00000a2e_656e6f44,
        64'h00000000_000a6b6f,
        64'h0000203a_73252020,
        64'h00000073_73657264,
        64'h6441206b_63757453,
        64'h00000000_00000a3a,
        64'h00000000_0075252f,
        64'h00752520_706f6f4c,
        64'h00000000_000a7025,
        64'h7830206f_74207025,
        64'h78302073_69206567,
        64'h6e617220_74736574,
        64'h00000000_00082008,
        64'h00000000_00000008,
        64'h08080808_08080808,
        64'h08082020_20202020,
        64'h20202020_20080808,
        64'h08080808_08080808,
        64'h00000000_0000000a,
        64'h2e2e2e74_73657420,
        64'h7478656e_206f7420,
        64'h676e6970_70696b53,
        64'h00000000_000a2e78,
        64'h25783020_74657366,
        64'h666f2074_6120656e,
        64'h696c2073_73657264,
        64'h64612064_61622065,
        64'h6c626973_736f7020,
        64'h3a455255_4c494146,
        64'h00000000_00007525,
        64'h20676e69_74736574,
        64'h00000000_00007525,
        64'h20676e69_74746573,
        64'h00000000_00080808,
        64'h08080808_08080808,
        64'h00000000_00202020,
        64'h20202020_20202020,
        64'h00000000_0000000a,
        64'h7025203d_20327020,
        64'h2c702520_3d203170,
        64'h00000a2e_78257830,
        64'h20746573_66666f20,
        64'h74612078_25783020,
        64'h3d212078_25783020,
        64'h3a455255_4c494146,
        64'h00000000_000a7325,
        64'h206e6f69_74636e75,
        64'h66202c64_2520656e,
        64'h696c202c_73252065,
        64'h6c696620_2c64656c,
        64'h69616620_7325206e,
        64'h6f697472_65737361,
        64'h00000a72_6564616f,
        64'h6c20746f_6f622065,
        64'h67617473_20747372,
        64'h69662064_65736162,
        64'h20746f6f_622d750a,
        64'h00000000_216b7369,
        64'h6420746e_756f6d75,
        64'h206f7420_6c696166,
        64'h00000000_0021656c,
        64'h69662065_736f6c63,
        64'h206f7420_6c696166,
        64'h0000000a_21746f6f,
        64'h62206e65_706f206f,
        64'h74206465_6c696146,
        64'h00000000_00000000,
        64'h6e69622e_746f6f62,
        64'h00000000_00000a79,
        64'h726f6d65_6d206f74,
        64'h6e69206e_69622e74,
        64'h6f6f6220_64616f4c,
        64'h00000000_0000000a,
        64'h21726576_69726420,
        64'h44532074_6e756f6d,
        64'h206f7420_6c696146,
        64'h00000000_0000000a,
        64'h2e2e2e70_25207373,
        64'h65726464_61207461,
        64'h206d6172_676f7270,
        64'h20646564_616f6c20,
        64'h65687420_746f6f42,
        64'h00000000_5c2d2f7c,
        64'h000a7825_203d206c,
        64'h61757463_61202c58,
        64'h25203d20_64657269,
        64'h75716572_206e656c,
        64'h00000000_00000000,
        64'h0a2e6e6f_69746172,
        64'h65706f20_50544654,
        64'h206c6167_656c6c49,
        64'h00000000_000a2e64,
        64'h656c6c61_63207172,
        64'h775f656c_646e6168,
        64'h00000000_00000a2e,
        64'h646e6520_656c6966,
        64'h20657669_65636552,
        64'h00000000_00000000,
        64'h0a64253d_657a6973,
        64'h6b636f6c_62202c22,
        64'h73252220_3a717277,
        64'h00000000_0000002f,
        64'h00000000_000a646c,
        64'h25202e67_6e6f6c20,
        64'h6f6f7420_68746170,
        64'h20747365_75716552,
        64'h00000064_6c252065,
        64'h646f6320_68746977,
        64'h2064656c_69616620,
        64'h64616572_20666c65,
        64'h000a7972_6f6d656d,
        64'h20524444_206f7420,
        64'h666c6520_64616f6c,
        64'h00000000_00000000,
        64'h0a732520_3d202964,
        64'h252c7025_2835646d,
        64'h00000000_0000000a,
        64'h6425203d_20687467,
        64'h6e656c20_656c6946,
        64'h00000000_00636d6d,
        64'h00000029_73252820,
        64'h00006425_203a7325,
        64'h00000000_434d4d65,
        64'h00000000_00004453,
        64'h00000000_00000000,
        64'h0a646e75_6f662074,
        64'h6f6e2064_25206563,
        64'h69766544_20434d4d,
        64'h0000297a_484d3030,
        64'h32282030_30325348,
        64'h00000000_00297a48,
        64'h4d383032_28203430,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282030,
        64'h35524444_20534855,
        64'h00000000_0000297a,
        64'h484d3030_31282030,
        64'h35524453_20534855,
        64'h00000000_00000029,
        64'h7a484d30_35282035,
        64'h32524453_20534855,
        64'h00000000_00000029,
        64'h7a484d35_32282032,
        64'h31524453_20534855,
        64'h00000000_00000029,
        64'h7a484d32_35282032,
        64'h35524444_20434d4d,
        64'h0000297a_484d3235,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000029_7a484d30,
        64'h35282064_65657053,
        64'h20686769_48204453,
        64'h0000297a_484d3632,
        64'h28206465_65705320,
        64'h68676948_20434d4d,
        64'h00000000_00000079,
        64'h63616765_4c204453,
        64'h00000000_00007963,
        64'h6167656c_20434d4d,
        64'h00000064_252e6425,
        64'h00000000_63256325,
        64'h63256325_63256325,
        64'h00000078_34302578,
        64'h34302520_726e5320,
        64'h78363025_206e614d,
        64'h00000000_00000a21,
        64'h646e756f_66206473,
        64'h635f7478_65206f4e,
        64'h00000000_00000000,
        64'h0a65646f_6d206120,
        64'h7463656c_6573206f,
        64'h7420656c_62616e75,
        64'h00000000_00000000,
        64'h0a217463_656c6573,
        64'h20656761_746c6f76,
        64'h206f7420_646e6f70,
        64'h73657220_746f6e20,
        64'h64696420_64726143,
        64'h0000000a_746e6573,
        64'h65727020_64726163,
        64'h206f6e20_3a434d4d,
        64'h00000000_0000000a,
        64'h64656e6f_69746974,
        64'h72617020_79646165,
        64'h726c6120_64726143,
        64'h00000000_000a7367,
        64'h6e697474_65732079,
        64'h74696c69_6261696c,
        64'h65722065_74697277,
        64'h206e6f69_74697472,
        64'h61702064_656c6c6f,
        64'h72746e6f_63207473,
        64'h6f682074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000a29_7525203e,
        64'h20752528_206d756d,
        64'h6978616d_20736465,
        64'h65637865_20657a69,
        64'h73206465_636e6168,
        64'h6e65206c_61746f54,
        64'h00000000_0000000a,
        64'h65747562_69727474,
        64'h61206465_636e6168,
        64'h6e652074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0a64656e,
        64'h67696c61_20657a69,
        64'h73207075_6f726720,
        64'h50572043_4820746f,
        64'h6e206e6f_69746974,
        64'h72617020_69255047,
        64'h0000000a_64656e67,
        64'h696c6120_657a6973,
        64'h2070756f_72672050,
        64'h57204348_20746f6e,
        64'h20616572_61206465,
        64'h636e6168_6e652061,
        64'h74616420_72657355,
        64'h00000a65_7a697320,
        64'h70756f72_67205057,
        64'h20434820_656e6966,
        64'h65642074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_000a676e,
        64'h696e6f69_74697472,
        64'h61702074_726f7070,
        64'h75732074_6f6e2073,
        64'h656f6420_64726143,
        64'h00000000_0000000a,
        64'h61657261_20617461,
        64'h64207265_73752064,
        64'h65636e61_686e6520,
        64'h726f6620_64657269,
        64'h75716572_20342e34,
        64'h203d3e20_434d4d65,
        64'h00000000_000a2978,
        64'h6c257830_2878616d,
        64'h20736465_65637865,
        64'h20786c25_78302072,
        64'h65626d75_6e206b63,
        64'h6f6c6220_3a434d4d,
        64'h00000000_00000a64,
        64'h6d632070_6f747320,
        64'h646e6573_206f7420,
        64'h6c696166_20636d6d,
        64'h00000000_000a7964,
        64'h61657220_64726163,
        64'h20676e69_74696177,
        64'h2074756f_656d6954,
        64'h0000000a_58383025,
        64'h7830203a_726f7272,
        64'h45207375_74617453,
        64'h00000000_65646f6d,
        64'h206e776f_6e6b6e55,
        64'h00000000_00006473,
        64'h5f637369_72776f6c,
        64'h00000078_25782520,
        64'h00000020_3a78250a,
        64'h00000000_0a732574,
        64'h69622d64_25203a68,
        64'h74646957_20737542,
        64'h00000000_0000203a,
        64'h79746963_61706143,
        64'h00000000_00000a73,
        64'h25203a79_74696361,
        64'h70614320_68676948,
        64'h00000a64_25203a64,
        64'h65657053_20737542,
        64'h00000000_00000a20,
        64'h63256325_63256325,
        64'h6325203a_656d614e,
        64'h00000000_00000000,
        64'h0a782520_3a4d454f,
        64'h00000000_0a782520,
        64'h3a444920_72657275,
        64'h74636166_756e614d,
        64'h00000000_000a7325,
        64'h203a6563_69766544,
        64'h00202020_3a434d4d,
        64'h00000000_52444420,
        64'h00000000_00006f4e,
        64'h00000000_00736559,
        64'h0000000a_7825203d,
        64'h2074736f_68202c78,
        64'h25207461_20646574,
        64'h61657263_20636d6d,
        64'h00000000_00000a64,
        64'h25206f74_20646567,
        64'h6e616863_206b7361,
        64'h6d202c64_65747265,
        64'h736e6920_64726143,
        64'h00000000_0000000a,
        64'h6425206f_74206465,
        64'h676e6168_63206b73,
        64'h616d202c_6465766f,
        64'h6d657220_64726143,
        64'h000a7475_6f656d69,
        64'h74207325_203a6473,
        64'h5f637369_72776f6c,
        64'h00726464_615f6573,
        64'h61625f64_73203d3d,
        64'h20657361_625f6473,
        64'h00000000_00000063,
        64'h2e636d6d_5f637369,
        64'h72776f6c_2f637273,
        64'h00000000_00000000,
        64'h66656463_62613938,
        64'h37363534_33323130,
        64'h007f7c5d_5b3f3e3d,
        64'h3c3b3a2e_2c2b2a22,
        64'h00007f7c_5d5b3f3e,
        64'h3d3c3b3a_2c2b2a22,
        64'h0000000a_2e783230,
        64'h253a7832_30253a78,
        64'h3230253a_78323025,
        64'h3a783230_253a7832,
        64'h3025203d_20737365,
        64'h72646461_2043414d,
        64'h00000a78_6c253a78,
        64'h6c25203d_2043414d,
        64'h00000000_00000a78,
        64'h25203d20_5d64255b,
        64'h4d454f20_49505351,
        64'h000a7264_64612043,
        64'h414d2070_75746553,
        64'h0000000a_21747075,
        64'h72726574_6e692064,
        64'h656c646e_61686e75,
        64'h00000000_00000a78,
        64'h25783020_3d206570,
        64'h79745f6f_746f7270,
        64'h00000000_0a297825,
        64'h28206465_74726f70,
        64'h7075736e_75203d20,
        64'h6f746f72_70205049,
        64'h000a5741_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a534c50_4d203d20,
        64'h6f746f72_50205049,
        64'h00000000_000a4554,
        64'h494c5044_55203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505443_53203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a504d4f_43203d20,
        64'h6f746f72_50205049,
        64'h00000000_0000004d,
        64'h00000000_0000000a,
        64'h5041434e_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000a48,
        64'h50544545_42203d20,
        64'h6f746f72_50205049,
        64'h000a5054_4d203d20,
        64'h6f746f72_50205049,
        64'h00000a48_41203d20,
        64'h6f746f72_50205049,
        64'h000a5053_45203d20,
        64'h6f746f72_50205049,
        64'h000a4552_47203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000000,
        64'h0a505653_52203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000036,
        64'h00000000_00000000,
        64'h0a504343_44203d20,
        64'h6f746f72_50205049,
        64'h00000a50_54203d20,
        64'h6f746f72_50205049,
        64'h000a5044_49203d20,
        64'h6f746f72_50205049,
        64'h000a3a73_746e6574,
        64'h6e6f6320_74736574,
        64'h0000000a_3a726564,
        64'h61656820_74736574,
        64'h000a5055_50203d20,
        64'h6f746f72_50205049,
        64'h000a5047_45203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000054,
        64'h00000000_00000000,
        64'h0a504950_49203d20,
        64'h6f746f72_50205049,
        64'h00000000_00000047,
        64'h00006425_2b544553,
        64'h46464f5f_524c5052,
        64'h00000000_3f3f3f3f,
        64'h00000000_00544553,
        64'h46464f5f_524c5052,
        64'h00000000_00544553,
        64'h46464f5f_44414252,
        64'h00000000_00005445,
        64'h5346464f_5f525352,
        64'h00000000_00544553,
        64'h46464f5f_53434652,
        64'h00544553_46464f5f,
        64'h4c525443_4f49444d,
        64'h00000000_00544553,
        64'h46464f5f_53434654,
        64'h00000000_00544553,
        64'h46464f5f_524c5054,
        64'h00000000_54455346,
        64'h464f5f49_4843414d,
        64'h00000000_54455346,
        64'h464f5f4f_4c43414d,
        64'h00000000_000a3b29,
        64'h78257830_2c302c78,
        64'h25287465_736d656d,
        64'h00000000_0a3b2978,
        64'h2578302c_78257830,
        64'h2c782528_6e666c65,
        64'h00000a70_2520726f,
        64'h72726520_7974696e,
        64'h61732072_64646170,
        64'h00000020_3a5d6425,
        64'h5b6e6f69_74636553,
        64'h000a7325_20202020,
        64'h00786c6c_2a302520,
        64'h00003a78_6c383025,
        64'h00732542_69632520,
        64'h00000000_00732573,
        64'h65747942_20756c25,
        64'h0073257a_48632520,
        64'h00000000_646c252e,
        64'h00000000_00756c25,
        64'h00000000_00000000,
        64'h73257a48_20756c25,
        64'h00000000_00007325,
        64'h00000000_00732520,
        64'h3a646c69_7542202c,
        64'h00000000_73257325,
        64'h00000000_00000a0a,
        64'h00000058_32302520,
        64'h00000000_0000002e,
        64'h00000000_00006325,
        64'h00000000_00000020,
        64'h20202020_20202020,
        64'h000a5245_46464f5f,
        64'h50434844_20726f66,
        64'h20676e69_74696157,
        64'h00000a73_25203a73,
        64'h25206563_69766564,
        64'h206e6f20_59524556,
        64'h4f435349_44205043,
        64'h48442064_6e657320,
        64'h74276e64_6c756f43,
        64'h000a5832_30253a58,
        64'h3230253a_58323025,
        64'h3a583230_253a5832,
        64'h30253a58_32302520,
        64'h3a204341_4d207325,
        64'h00000000_30687465,
        64'h00000000_000a2973,
        64'h2528726f_72726570,
        64'h000a5952_45564f43,
        64'h5349445f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_0000000a,
        64'h64252065_646f6370,
        64'h6f205043_48442064,
        64'h656c646e_61686e55,
        64'h00000000_0a642520,
        64'h6e6f6974_706f2064,
        64'h656c646e_61686e75,
        64'h00000000_0000000a,
        64'h73252072_6f727245,
        64'h00000000_00000a64,
        64'h65737566_65722073,
        64'h73657264_64612064,
        64'h65747365_75716552,
        64'h00000000_0000000a,
        64'h4b414e20_50434844,
        64'h00000000_0a444550,
        64'h50494b53_204b4341,
        64'h000a2273_2522203d,
        64'h20656d61_6e74736f,
        64'h4820746e_65696c43,
        64'h00000a22_73252220,
        64'h3d206e69_616d6f44,
        64'h00000000_0000000a,
        64'h7364253a_6d64253a,
        64'h68642520_3d20656d,
        64'h69742065_7361654c,
        64'h000a6425_2e64252e,
        64'h64252e64_2520203a,
        64'h73736572_64646120,
        64'h6b73616d_2074654e,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h61207265_74756f52,
        64'h00000000_00000000,
        64'h0a64252e_64252e64,
        64'h252e6425_20203a73,
        64'h73657264_64412050,
        64'h49207265_76726553,
        64'h0000000a_64252e64,
        64'h252e6425_2e642520,
        64'h203a7373_65726464,
        64'h41205049_20746e65,
        64'h696c4320_50434844,
        64'h00000000_0000000a,
        64'h4b434120_50434844,
        64'h0000000a_54534555,
        64'h5145525f_50434844,
        64'h20676e69_646e6553,
        64'h00000000_00000000,
        64'h0a702520_2c726f72,
        64'h7265206c_616e7265,
        64'h746e6920_70636864,
        64'h00000a29_73252c73,
        64'h25287075_6b6f6f6c,
        64'h000a6563_69766564,
        64'h206e776f_6e6b6e75,
        64'h00000000_203a6425,
        64'h20656369_7665440a,
        64'h00203a64_25206563,
        64'h69766564_2073250a,
        64'h00000000_00203a64,
        64'h25206563_69766544,
        64'h00000000_00000000,
        64'h73736572_6464612d,
        64'h63616d2d_6c61636f,
        64'h6c006874_6469772d,
        64'h6f692d67_65720074,
        64'h66696873_2d676572,
        64'h00737470_75727265,
        64'h746e6900_746e6572,
        64'h61702d74_70757272,
        64'h65746e69_00646565,
        64'h70732d74_6e657272,
        64'h75630076_65646e2c,
        64'h76637369_72007974,
        64'h69726f69_72702d78,
        64'h616d2c76_63736972,
        64'h0073656d_616e2d67,
        64'h65720064_65646e65,
        64'h7478652d_73747075,
        64'h72726574_6e690073,
        64'h65676e61_7200656c,
        64'h646e6168_702c7875,
        64'h6e696c00_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h00100000_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_00000064,
        64'h6e727768_2d637369,
        64'h72776f6c_1b000000,
        64'h0e000000_03000000,
        64'h00003030_30303030,
        64'h30344064_6e727768,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h00800000_00000000,
        64'h00000030_00000000,
        64'h67000000_10000000,
        64'h03000000_00007fe3,
        64'h023e1800_47010000,
        64'h06000000_03000000,
        64'h03000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_00636d6d,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_02000000,
        64'h25010000_04000000,
        64'h03000000_02000000,
        64'h14010000_04000000,
        64'h03000000_00000100,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40636d6d,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h04000000_3a010000,
        64'h04000000_03000000,
        64'h02000000_30010000,
        64'h04000000_03000000,
        64'h01000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h00c20100_06010000,
        64'h04000000_03000000,
        64'h80f0fa02_4b000000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000010_00000000,
        64'h67000000_10000000,
        64'h03000000_00303537,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000000,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'hffff0000_01000000,
        64'hca000000_08000000,
        64'h03000000_00333130,
        64'h2d677562_65642c76,
        64'h63736972_1b000000,
        64'h10000000_03000000,
        64'h00003040_72656c6c,
        64'h6f72746e_6f632d67,
        64'h75626564_01000000,
        64'h02000000_02000000,
        64'hbb000000_04000000,
        64'h03000000_02000000,
        64'hb5000000_04000000,
        64'h03000000_03000000,
        64'hfb000000_04000000,
        64'h03000000_07000000,
        64'he8000000_04000000,
        64'h03000000_00000004,
        64'h00000000_0000000c,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h09000000_01000000,
        64'h0b000000_01000000,
        64'hca000000_10000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00000c00,
        64'h00000000_00000002,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_01000000,
        64'h03000000_01000000,
        64'hca000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6e696c63,
        64'h01000000_c3000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000008_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h01000000_bb000000,
        64'h04000000_03000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00007663_73697200,
        64'h656e6169_7261202c,
        64'h7a687465_1b000000,
        64'h13000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha8060000_59010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'he0060000_38000000,
        64'h39080000_edfe0dd0,
        64'h00000000_fffff9ae,
        64'hfffff974_fffff99c,
        64'hfffff974_fffff98a,
        64'hfffff976_fffff962,
        64'h00000000_64726143,
        64'h2d445320_726f6620,
        64'h746f6f62_2d752064,
        64'h6573696d_696e696d,
        64'h20435349_52776f4c,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00020000_00010000,
        64'h0000c000_00008000,
        64'h00006000_00004000,
        64'h00002000_00001000,
        64'h00000800_00000400,
        64'h00000200_00000100,
        64'h00000080_00000040,
        64'h00000020_00000000,
        64'h0bebc200_0c65d400,
        64'h02faf080_05f5e100,
        64'h02faf080_017d7840,
        64'h03197500_03197500,
        64'h02faf080_018cba80,
        64'h017d7840_017d7840,
        64'h00989680_000f4240,
        64'h000186a0_00002710,
        64'h50463c37_322d2823,
        64'h1e19140f_0d0c0a00,
        64'h00000000_00000000,
        64'h00000000_10000000,
        64'h00000001_00000000,
        64'h20000000_00000002,
        64'h00000000_40000000,
        64'h00000005_00000001,
        64'h20000000_00000006,
        64'h00000001_40000000,
        64'h70000000_00000000,
        64'h70000000_00000002,
        64'h70000000_00000004,
        64'h60000000_00000005,
        64'h30000000_00000001,
        64'h30000000_00000003,
        64'h00000000_40050100,
        64'h40050000_40040500,
        64'h40040401_40040400,
        64'h40040300_40040200,
        64'h40040100_40040000,
        64'h00000000_87feb570,
        64'h00000000_87feb558,
        64'h00000000_87feb540,
        64'h00000000_87feb528,
        64'h00000000_87feb510,
        64'h00000000_87feb4f8,
        64'h00000000_87feb4e0,
        64'h00000000_87feb4c8,
        64'h00000000_87feb4b0,
        64'h00000000_87feb498,
        64'h00000000_87feb488,
        64'h00000000_87feb478,
        64'hffffc9ba_ffffc9b4,
        64'hffffc9ae_ffffc80a,
        64'hffffb998_ffffb998,
        64'hffffb998_ffffb998,
        64'hffffb994_ffffb990,
        64'hffffb990_ffffb96c,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_87fe4d18,
        64'h00000000_87fe4aba,
        64'h00000000_87fe4eaa,
        64'h00646374_65675f63,
        64'h6d6d5f64_72616f62,
        64'h00000002_0000ffff,
        64'h004c4b40_004c4b40,
        64'h00300000_20000000,
        64'h00000000_87fe9e88,
        64'h00000000_87feb160,
        64'h00717269_5f646e65,
        64'h5f617461_645f6473,
        64'h5f637369_72776f6c,
        64'h00000000_00007172,
        64'h695f646d_635f6473,
        64'h5f637369_72776f6c,
        64'h00007172_695f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0067616c,
        64'h665f7470_75727265,
        64'h746e695f_74696177,
        64'h5f637369_72776f6c,
        64'h00000000_646d635f,
        64'h74726174_735f6473,
        64'h5f637369_72776f6c,
        64'h00000000_0000006e,
        64'h655f7172_695f6473,
        64'h00000000_00007475,
        64'h6f656d69_745f6473,
        64'h00000000_0000657a,
        64'h69736b6c_625f6473,
        64'h00000000_00000074,
        64'h6e636b6c_625f6473,
        64'h00000000_00000000,
        64'h74657365_725f6473,
        64'h00000000_74726174,
        64'h735f646d_635f6473,
        64'h00000000_0000676e,
        64'h69747465_735f6473,
        64'h00000000_00007669,
        64'h645f6b6c_635f6473,
        64'h00000000_00000000,
        64'h6e67696c_615f6473,
        64'h00000000_00006465,
        64'h6c5f7465_735f6473,
        64'h5f637369_72776f6c,
        64'h09020b04_0d060f08,
        64'h010a030c_050e0700,
        64'h020f0c09_0603000d,
        64'h0a070401_0e0b0805,
        64'h0c07020d_08030e09,
        64'h040f0a05_000b0601,
        64'heb86d391_2ad7d2bb,
        64'hbd3af235_f7537e82,
        64'h4e0811a1_a3014314,
        64'hfe2ce6e0_6fa87e4f,
        64'h85845dd1_ffeff47d,
        64'h8f0ccc92_655b59c3,
        64'hfc93a039_ab9423a7,
        64'h432aff97_f4292244,
        64'hc4ac5665_1fa27cf8,
        64'he6db99e5_d9d4d039,
        64'h04881d05_d4ef3085,
        64'heaa127fa_289b7ec6,
        64'hbebfbc70_f6bb4b60,
        64'h4bdecfa9_a4beea44,
        64'hfde5380c_6d9d6122,
        64'h8771f681_fffa3942,
        64'h8d2a4c8a_676f02d9,
        64'hfcefa3f8_a9e3e905,
        64'h455a14ed_f4d50d87,
        64'hc33707d6_21e1cde6,
        64'he7d3fbc8_d8a1e681,
        64'h02441453_d62f105d,
        64'he9b6c7aa_265e5a51,
        64'hc040b340_f61e2562,
        64'h49b40821_a679438e,
        64'hfd987193_6b901122,
        64'h895cd7be_ffff5bb1,
        64'h8b44f7af_698098d8,
        64'hfd469501_a8304613,
        64'h4787c62a_f57c0faf,
        64'hc1bdceee_242070db,
        64'he8c7b756_d76aa478,
        64'h02020202_02020202,
        64'h10020202_02020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02010101_01010101,
        64'h10010101_01010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h08101010_10020202,
        64'h02020202_02020202,
        64'h02020202_02020202,
        64'h02424242_42424210,
        64'h10101010_10010101,
        64'h01010101_01010101,
        64'h01010101_01010101,
        64'h01414141_41414110,
        64'h10101010_10100404,
        64'h04040404_04040404,
        64'h10101010_10101010,
        64'h10101010_101010a0,
        64'h08080808_08080808,
        64'h08080808_08080808,
        64'h08082828_28282808,
        64'h08080808_08080808,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hbf5db7bf_f0efd5df,
        64'hb0ef0da5_05130000,
        64'h2517b7e1_c60f80ef,
        64'hd6ffb0ef_0dc50513,
        64'h00002517_bfe9aa3f,
        64'hf0efd81f_b0ef0de5,
        64'h05130000_2517b7f5,
        64'hedbff0ef_8522d95f,
        64'hb0ef0e25_05130000,
        64'h2517a001_941fe0ef,
        64'h8522da9f_b0ef0e65,
        64'h05130000_25178782,
        64'h97ba439c_97ba078a,
        64'h6b070713_00000717,
        64'h02f76463_47190054,
        64'h579b0ff4_7413fd39,
        64'h1be3dd9f_b0ef2581,
        64'h8552688c_0004b823,
        64'hde7fb0ef_86222401,
        64'h25816080_608ce09c,
        64'h09058556_0007c783,
        64'h016907b3_4991126a,
        64'h0a130000_2a17116a,
        64'h8a930000_2a974400,
        64'h04b723ab_0b130000,
        64'h2b174901_be0f80ef,
        64'hfe9416e3_e2bfb0ef,
        64'h0405854a_0004059b,
        64'h639097ce_00341793,
        64'h449513a9_09130000,
        64'h29174400_09b74401,
        64'hfccfe0ef_13c50513,
        64'h00002517_fa6fe0ef,
        64'he05ae456_e852ec4e,
        64'hf04af426_f822fc06,
        64'h7139feef_e06f1fe5,
        64'h05130000_25179e7f,
        64'he06f0141_60a2e85f,
        64'hb06f0141_cec50513,
        64'h00002517_40a005b3,
        64'h60a20005_5c63b7df,
        64'h70eff2a5_05130000,
        64'h0517ea9f_b0efe406,
        64'hcf850513_00002517,
        64'h1141bf69_2441ebdf,
        64'hb0ef855a_ff5492e3,
        64'hec7fb0ef_8552d93f,
        64'hf0ef2485_45890007,
        64'hc50397ce_93811782,
        64'h009407bb_4481ee5f,
        64'hb0ef8552_db1ff0ef,
        64'h852245a1_bf69008b,
        64'hb02304a1_df3ff0ef,
        64'h00c4541b_85d22421,
        64'h80826125_6be27b02,
        64'h7aa27a42_79e26906,
        64'h64a66446_60e60324,
        64'h6763eaab_0b130000,
        64'h2b174ac1_31ca0a13,
        64'h00001a17_4401da3f,
        64'hd0ef002c_92018552,
        64'h16024089_063be3df,
        64'hf0ef002c_05546463,
        64'h0164053b_00998a33,
        64'h0004841b_44000bb7,
        64'hff860a9b_44818932,
        64'h8b2e89aa_f852e8a2,
        64'hec86ec5e_f05af456,
        64'hfc4ee0ca_e4a6711d,
        64'h80826125_7aa27a42,
        64'h79e26906_64a66446,
        64'h60e6f91f_b0eff1e5,
        64'h05130000_2517ff24,
        64'h91e3fa1f_b0ef854e,
        64'he6dff0ef_24854589,
        64'hff87c503_97ba9381,
        64'h10181782_009407bb,
        64'h49213b29_89930000,
        64'h19974481_fcbfb0ef,
        64'h3c050513_00001517,
        64'he9dff0ef_45a1854a,
        64'hfdffb0ef_f6c50513,
        64'h00002517_ff4992e3,
        64'hfeffb0ef_8556ebbf,
        64'hf0ef2985_45890007,
        64'hc50397a6_93811782,
        64'h013407bb_4a213fea,
        64'h8a930000_1a974981,
        64'h816fc0ef_40c50513,
        64'h00001517_ee9ff0ef,
        64'h854a45a1_82afc0ef,
        64'hfb850513_00002517,
        64'hff4991e3_83afc0ef,
        64'h8556f07f_f0ef2985,
        64'h4589ff07_c50397ba,
        64'h93811018_17820134,
        64'h07bb4a21_44ca8a93,
        64'h00001a97_4981864f,
        64'hc0ef45a5_05130000,
        64'h1517f37f_f0ef854a,
        64'h45a1fcd7_99e30785,
        64'h00e60023_00e55733,
        64'h963e0830_00b60023,
        64'h00e9d5b3_00f48633,
        64'h00b60023_00ea55b3,
        64'h0387071b_963e0810,
        64'h02f8073b_46a15861,
        64'h4781f2bf_f0ef454d,
        64'h45894601_89aa0034,
        64'hf39ff0ef_454d8a2a,
        64'h45894601_0034f47f,
        64'hf0eff456_f852fc4e,
        64'hc43aec86_c63e4589,
        64'h454d84ae_842a4601,
        64'h0034e4a6_e8a20587,
        64'he7938f55_0089179b,
        64'h0189571b_30068693,
        64'h00a7893b_6685e0ca,
        64'h004007b7_711da45f,
        64'he06f0141_60a26402,
        64'h00044503_943e3ee7,
        64'h87930000_2797883d,
        64'hfedff0ef_0045551b,
        64'h35fd00b7_d763842a,
        64'h4785e406_e0221141,
        64'hbfc1f618_07850007,
        64'h67039736_00279713,
        64'h80827388_440007b7,
        64'hffe537fd_c3198b09,
        64'h7a984400_06b73e80,
        64'h079300b7_6f630007,
        64'h871b4400_06374781,
        64'h2581f788_440007b7,
        64'h8d510106_161b8d5d,
        64'h0085979b_80822501,
        64'h7b884400_07b78082,
        64'h25016b88_0007b823,
        64'h440007b7_80822501,
        64'h63884400_07b78082,
        64'he3884400_07b79101,
        64'h1502bff1_f5dff0ef,
        64'h4541f63f_f0ef4521,
        64'hf69ff0ef_4511f6ff,
        64'hf0ef4509_f75ff0ef,
        64'h4505f7bf_f0ef4501,
        64'he4061141_bf51c000,
        64'h28f3c020_26f3fac7,
        64'h10e39f0f_c06f47e5,
        64'h05130000_251702a7,
        64'h473302a7_67b302b3,
        64'h45bb02c7_47334000,
        64'h059302a6_87334116,
        64'h86b33e80_0513c000,
        64'h26f38e15_c0202673,
        64'h02b71d63_2705fe08,
        64'h13e397aa_387d0007,
        64'h802397aa_00078023,
        64'h97aa0007_802397aa,
        64'h00078023_40000813,
        64'h87f245a9_01f61e13,
        64'h46814881_470100c5,
        64'h131b4605_80828082,
        64'h614569a2_694264e2,
        64'h740270a2_ff2417e3,
        64'he73ff0ef_24050135,
        64'h85334605_46850084,
        64'h95b34979_01f49993,
        64'h4441a90f_c0ef4485,
        64'h22050513_00002517,
        64'ha9efc0ef_4e450513,
        64'h00002517_aaafc0ef,
        64'h4c050513_00002517,
        64'hab6fc0ef_4a450513,
        64'h00002517_04000593,
        64'hc45fe0ef_e44ee84a,
        64'hec26f022_f4064a65,
        64'h05130000_25177179,
        64'hbf890485_ae2fc0ef,
        64'h27050513_00002517,
        64'hb7d14a89_af2fc0ef,
        64'h4b850513_00002517,
        64'h97828522_95a20049,
        64'h56130019_5593008a,
        64'h3783b10f_c0ef4ce5,
        64'h05130000_2517c985,
        64'h000a3583_02f74c63,
        64'h6722010a_2783b2cf,
        64'hc0ef856e_e129952f,
        64'hf0ef8522_6582b3cf,
        64'hc0ef856a_85e6b44f,
        64'hc0ef8562_b4afc0ef,
        64'h855e85ce_00098663,
        64'hb56fc0ef_855a85a6,
        64'h80826109_6de27d02,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e67906,
        64'h74a68556_744670e6,
        64'hb7efc0ef_54c50513,
        64'h00002517_0299f863,
        64'h058a0a13_00003a17,
        64'h558d8d93_00002d97,
        64'h558d0d13_00002d17,
        64'h550c8c93_00002c97,
        64'h550c0c13_00002c17,
        64'h550b8b93_00002b97,
        64'h550b0b13_00002b17,
        64'h44854a81_e03e0039,
        64'h5793bd0f_c0efe436,
        64'hfc86ec6e_f06af466,
        64'hf862fc5e_e0dae4d6,
        64'he8d2f4a6_55c50513,
        64'h00002517_85aa842a,
        64'h892e962a_f0caf8a2,
        64'hfff58613_89b2ecce,
        64'h71198082_6505bfb1,
        64'h547dbf05_0d85e99f,
        64'he0ef0007_c50397ea,
        64'h8b8d0007_8b1b001b,
        64'h079beadf_e0ef4521,
        64'hef910ba1_033df7b3,
        64'hff9795e3_00d61023,
        64'h92c116c2_078900fb,
        64'h86330006_d6830187,
        64'h86b34781_e28812a7,
        64'hbf230000_37978d41,
        64'h66e29101_14021502,
        64'h8c510106_161b8d5d,
        64'h0105151b_664267a2,
        64'hfe3fd0ef_e42afe9f,
        64'hd0efe82a_feffd0ef,
        64'h842aff5f_d0efec36,
        64'hb7754a05_80826149,
        64'h7da27d42_7ce26c06,
        64'h6ba66b46_6ae67a06,
        64'h79a67946_74e6640a,
        64'h60aa8522_cb2fc0ef,
        64'h62050513_00002517,
        64'h02fa1863_8aa68bca,
        64'h4785ed4d_842aa94f,
        64'hf0ef854a_85a6866e,
        64'h04fd9663_96d6003d,
        64'h96936782_4d8193ed,
        64'h0d130000_3d179c49,
        64'h89934ca1_1dcc0c13,
        64'h00003c17_4b014a09,
        64'h8ba6f85f_e0ef8aca,
        64'he032f46e_e122e506,
        64'hf86afc66_e0e2e4de,
        64'he8daecd6_f0d26985,
        64'h02000513_84ae892a,
        64'hf4cef8ca_fca67175,
        64'hbfb1547d_bf050d85,
        64'hfbbfe0ef_0007c503,
        64'h97ea8b8d_00078b1b,
        64'h001b079b_fcffe0ef,
        64'h4521ef91_0ba1033d,
        64'hf7b3ff97_95e300d6,
        64'h00230ff6_f6930785,
        64'h00fb8633_0006c683,
        64'h018786b3_4781e288,
        64'h24a7bc23_00003797,
        64'h8d4166e2_91011402,
        64'h15028c51_0106161b,
        64'h8d5d0105_151b6642,
        64'h67a2904f_e0efe42a,
        64'h90afe0ef_e82a910f,
        64'he0ef842a_916fe0ef,
        64'hec36b775_4a058082,
        64'h61497da2_7d427ce2,
        64'h6c066ba6_6b466ae6,
        64'h7a0679a6_794674e6,
        64'h640a60aa_8522dd4f,
        64'hc0ef7425_05130000,
        64'h251702fa_18638aa6,
        64'h8bca4785_ed4d842a,
        64'hbb6ff0ef_854a85a6,
        64'h866e04fd_966396d6,
        64'h003d9693_67824d81,
        64'ha60d0d13_00003d17,
        64'h9c498993_4ca12f6c,
        64'h0c130000_3c174b01,
        64'h4a098ba6_8a6ff0ef,
        64'h8acae032_f46ee122,
        64'he506f86a_fc66e0e2,
        64'he4dee8da_ecd6f0d2,
        64'h69850200_051384ae,
        64'h892af4ce_f8cafca6,
        64'h7175b7e9_5b7db749,
        64'h060500b8_3023e30c,
        64'h85d6e111_85e20016,
        64'h75138082_61096de2,
        64'h7d027ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_855a7446,
        64'h70e6e88f_c0ef7ce5,
        64'h05130000_2517fafb,
        64'h90e30400_07932b85,
        64'hfbb41be3_8c562405,
        64'he9318b2a_c72ff0ef,
        64'h854a85ce_6622eb4f,
        64'hc0ef856a_85daebcf,
        64'hc0efe432_855206f6,
        64'h1063974e_00e90833,
        64'h00361713_67824601,
        64'hfffc4a93_edafc0ef,
        64'h856685da_00848b3b,
        64'hee6fc0ef_85524401,
        64'h003b949b_01779c33,
        64'h47854da1_7d4d0d13,
        64'h00002d17_7ccc8c93,
        64'h00002c97_7c4a0a13,
        64'h00002a17_f12fc0ef,
        64'h4b81e032_89aef862,
        64'he0dae4d6_f4a6f8a2,
        64'hfc86ec6e_f06af466,
        64'hfc5ee8d2_ecce7de5,
        64'h05130000_2517892a,
        64'hf0ca7119_bf755dfd,
        64'hbfc5859a_fe080be3,
        64'h85bab761_0605e10c,
        64'he28c85c6_00080363,
        64'h85be008b_ea630016,
        64'h78138082_61096de2,
        64'h7d027ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_856e7446,
        64'h70e6f88f_c0ef8ce5,
        64'h05130000_3517f8f4,
        64'h1be30800_07932405,
        64'hed298daa_d6aff0ef,
        64'h852685ca_6622facf,
        64'hc0ef8566_85a2fb4f,
        64'hc0efe432_854e0546,
        64'h1c6396ca_00d48533,
        64'h00361693_4601fff7,
        64'hc893fff7_43138fd5,
        64'h008d16b3_00fd17b3,
        64'h0024079b_8f5d00ed,
        64'h173300fd_17b3408b,
        64'h07bb408a_873bff4f,
        64'hc0ef8562_85a2ffcf,
        64'hc0ef854e_8dcc8c93,
        64'h00003c97_03f00b93,
        64'h08100b13_4d0507f0,
        64'h0a938e2c_0c130000,
        64'h3c178da9_89930000,
        64'h3997829f_c0ef4401,
        64'h8a32892e_ec6efc86,
        64'hf06af466_f862fc5e,
        64'he0dae4d6_e8d2ecce,
        64'hf0caf8a2_8f450513,
        64'h00003517_84aaf4a6,
        64'h7119b7f1_5dfdbfe5,
        64'he19ce31c_bf610605,
        64'he194e314_008c6663,
        64'h80826109_6de27d02,
        64'h7ca27c42_7be26b06,
        64'h6aa66a46_69e67906,
        64'h74a6856e_744670e6,
        64'h88ffc0ef_9d450513,
        64'h00003517_fb5417e3,
        64'h2405e139_8daae6cf,
        64'hf0ef8526_85ca6622,
        64'h8affc0ef_856a85a2,
        64'h8b7fc0ef_e4328552,
        64'h05661a63_974a00e4,
        64'h85b30036_17134601,
        64'hfff6c693_fff7c793,
        64'h008996b3_00f997b3,
        64'h408b87bb_8e3fc0ef,
        64'h856685a2_8ebfc0ef,
        64'h85520800_0a939ced,
        64'h0d130000_3d1703f0,
        64'h0c134985_07f00b93,
        64'h9d0c8c93_00003c97,
        64'h9c8a0a13_00003a17,
        64'h917fc0ef_44018b32,
        64'h892eec6e_fc86f06a,
        64'hf466f862_fc5ee0da,
        64'he4d6e8d2_eccef0ca,
        64'hf8a29e25_05130000,
        64'h351784aa_f4a67119,
        64'hb7f15dfd_bfe5e298,
        64'he398bf61_0605e28c,
        64'he38c008c_66638082,
        64'h61096de2_7d027ca2,
        64'h7c427be2_6b066aa6,
        64'h6a4669e6_790674a6,
        64'h856e7446_70e697df,
        64'hc0efac25_05130000,
        64'h3517fb54_1be32405,
        64'he1398daa_f5aff0ef,
        64'h852685ca_662299df,
        64'hc0ef856a_85a29a5f,
        64'hc0efe432_85520566,
        64'h1a6397ca_00f486b3,
        64'h00361793_46010089,
        64'h95b300e9_9733408b,
        64'h873b9c9f_c0ef8566,
        64'h85a29d1f_c0ef8552,
        64'h08000a93_ab4d0d13,
        64'h00003d17_03f00c13,
        64'h498507f0_0b93ab6c,
        64'h8c930000_3c97aaea,
        64'h0a130000_3a179fdf,
        64'hc0ef4401_8b32892e,
        64'hec6efc86_f06af466,
        64'hf862fc5e_e0dae4d6,
        64'he8d2ecce_f0caf8a2,
        64'hac850513_00003517,
        64'h84aaf4a6_7119bff1,
        64'h59fdb74d_0605e29c,
        64'he31c8082_61256c42,
        64'h6be27b02_7aa27a42,
        64'h79e26906_64a6854e,
        64'h644660e6_a53fc0ef,
        64'hb9850513_00003517,
        64'hf94c19e3_0c05e91d,
        64'h89aa831f_f0ef8522,
        64'h85a66622_a73fc0ef,
        64'h855e85ce_a7bfc0ef,
        64'he432854a_05561763,
        64'h972600e4_06b30036,
        64'h17134601_8fd9038c,
        64'h17138fd9_030c1713,
        64'h8fd9028c_17138fd9,
        64'h020c1713_8fd9018c,
        64'h17130187_e7b38fd9,
        64'h008c1793_010c1713,
        64'habffc0ef_855a85ce,
        64'h000c099b_acbfc0ef,
        64'h854a1000_0a13baeb,
        64'h8b930000_3b97ba6b,
        64'h0b130000_3b17b9e9,
        64'h09130000_3917aedf,
        64'hc0ef4c01_8ab284ae,
        64'hfc4eec86_e862ec5e,
        64'hf05af456_f852e0ca,
        64'he4a6bb25_05130000,
        64'h3517842a_e8a2711d,
        64'hb7e15d7d_b7790605,
        64'he198e398_872ac291,
        64'h876a0016_7693bf49,
        64'h000b3d03_80826165,
        64'h6d426ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h694664e6_856a7406,
        64'h70a6b51f_c0efc965,
        64'h05130000_3517fb44,
        64'h1ae32405_e5298d2a,
        64'h92fff0ef_852685ca,
        64'h6622b71f_c0ef8566,
        64'h85a2b79f_c0efe432,
        64'h854e0556_1c6397ca,
        64'h00f485b3_00361793,
        64'hfffd4513_4601b95f,
        64'hc0ef8562_85a2000b,
        64'hbd03cba5_00147793,
        64'hba7fc0ef_854e0400,
        64'h0a13c8ac_8c930000,
        64'h3c97c82c_0c130000,
        64'h3c17f8ab_8b930000,
        64'h3b97f8ab_0b130000,
        64'h3b17c8a9_89930000,
        64'h3997bd9f_c0ef4401,
        64'h8ab2892e_e86af486,
        64'hec66f062_f45ef85a,
        64'hfc56e0d2_e4cee8ca,
        64'hf0a2ca25_05130000,
        64'h351784aa_eca67159,
        64'hbfc154fd_bf590605,
        64'he198e398_8726c291,
        64'h87660016_76938082,
        64'h61656ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h64e66946_85267406,
        64'h70a6c39f_c0efd7e5,
        64'h05130000_3517fb54,
        64'h1be32405_e12984aa,
        64'ha17ff0ef_854a85ce,
        64'h6622c59f_c0ef8562,
        64'h85a2c61f_c0efe432,
        64'h85520566_186397ce,
        64'h00f905b3_00361793,
        64'h14fd4601_40900cb3,
        64'hc7ffc0ef_8885855e,
        64'h85a2fff4_4493c8df,
        64'hc0ef8552_04000a93,
        64'hd70c0c13_00003c17,
        64'hd68b8b93_00003b97,
        64'hd60a0a13_00003a17,
        64'hcaffc0ef_44018b32,
        64'h89aeec66_eca6f486,
        64'hf062f45e_f85afc56,
        64'he0d2e4ce_f0a2d765,
        64'h05130000_3517892a,
        64'he8ca7159_bfc90705,
        64'h00a83023_e28800f7,
        64'h0533ab1f_f06f6121,
        64'h863a69e2_854e7902,
        64'h74a270e2_744200c7,
        64'h1c6396ae_00d98833,
        64'h00371693_47018fc5,
        64'h90811782_65a26602,
        64'h14828fc1_8cc90109,
        64'h179b0105_151b891f,
        64'he0ef84aa_897fe0ef,
        64'h892a89df_e0ef842a,
        64'h8a3fe0ef_89aaec4e,
        64'hf04af426_f822fc06,
        64'he032e42e_7139b7f1,
        64'h00e83023_8f690008,
        64'h3703e314_8ee90785,
        64'h6314b29f_f06f6121,
        64'h863e69e2_854e7902,
        64'h74a270e2_744200c7,
        64'h9c63974e_00e58833,
        64'h00379713_47818d5d,
        64'h91011782_65a26602,
        64'h15028fc1_8d450109,
        64'h179b0105_151b909f,
        64'he0ef84aa_90ffe0ef,
        64'h892a915f_e0ef842a,
        64'h91bfe0ef_89aaec4e,
        64'hf04af426_f822fc06,
        64'he032e42e_7139b7f1,
        64'h00e83023_8f490008,
        64'h3703e314_8ec90785,
        64'h6314ba1f_f06f6121,
        64'h863e69e2_854e7902,
        64'h74a270e2_744200c7,
        64'h9c63974e_00e58833,
        64'h00379713_47818d5d,
        64'h91011782_65a26602,
        64'h15028fc1_8d450109,
        64'h179b0105_151b981f,
        64'he0ef84aa_987fe0ef,
        64'h892a98df_e0ef842a,
        64'h993fe0ef_89aaec4e,
        64'hf04af426_f822fc06,
        64'he032e42e_7139b7d1,
        64'h00e83023_02a75733,
        64'h00083703_e31402a6,
        64'hd6b30785_63144505,
        64'he111c21f_f06f6121,
        64'h863e69e2_854e7902,
        64'h74a270e2_744200c7,
        64'h9c63974e_00e58833,
        64'h00379713_47818d5d,
        64'h91011782_65a26602,
        64'h15028fc1_8d450109,
        64'h179b0105_151ba01f,
        64'he0ef84aa_a07fe0ef,
        64'h892aa0df_e0ef842a,
        64'ha13fe0ef_89aaec4e,
        64'hf04af426_f822fc06,
        64'he032e42e_7139b7e1,
        64'h00e83023_02a70733,
        64'h00083703_e31402a6,
        64'h86b30785_6314c9df,
        64'hf06f6121_863e69e2,
        64'h854e7902_74a270e2,
        64'h744200c7_9c63974e,
        64'h00e58833_00379713,
        64'h47818d5d_91011782,
        64'h65a26602_15028fc1,
        64'h8d450109_179b0105,
        64'h151ba7df_e0ef84aa,
        64'ha83fe0ef_892aa89f,
        64'he0ef842a_a8ffe0ef,
        64'h89aaec4e_f04af426,
        64'hf822fc06_e032e42e,
        64'h7139b7f1_00e83023,
        64'h8f090008_3703e314,
        64'h8e890785_6314d15f,
        64'hf06f6121_863e69e2,
        64'h854e7902_74a270e2,
        64'h744200c7_9c63974e,
        64'h00e58833_00379713,
        64'h47818d5d_91011782,
        64'h65a26602_15028fc1,
        64'h8d450109_179b0105,
        64'h151baf5f_e0ef84aa,
        64'hafbfe0ef_892ab01f,
        64'he0ef842a_b07fe0ef,
        64'h89aaec4e_f04af426,
        64'hf822fc06_e032e42e,
        64'h7139b7f1_00e83023,
        64'h8f290008_3703e314,
        64'h8ea90785_6314d8df,
        64'hf06f6121_863e69e2,
        64'h854e7902_74a270e2,
        64'h744200c7_9c63974e,
        64'h00e58833_00379713,
        64'h47818d5d_91011782,
        64'h65a26602_15028fc1,
        64'h8d450109_179b0105,
        64'h151bb6df_e0ef84aa,
        64'hb73fe0ef_892ab79f,
        64'he0ef842a_b7ffe0ef,
        64'h89aaec4e_f04af426,
        64'hf822fc06_e032e42e,
        64'h7139b7ad_0485ab1f,
        64'hf0ef0007_c50397e2,
        64'h0039f793_0985ac1f,
        64'hf0ef4521_ef8100ad,
        64'hb02300ac_b0238d41,
        64'h91011402_150201a4,
        64'h643300a9_6533010d,
        64'h1d1b0105_151b0344,
        64'hf7b3bd5f_e0ef892a,
        64'hbdbfe0ef_8d2abe1f,
        64'he0ef842a_be7fe0ef,
        64'he47ff06f_61657ae2,
        64'h85567b42_64e685da,
        64'h86266da2_6d426ce2,
        64'h7c027ba2_6a0669a6,
        64'h694670a6_74068a4f,
        64'hd0ef2125_05130000,
        64'h35170374_9b6300fb,
        64'h0cb300fa_8db30034,
        64'h979351ac_0c130000,
        64'h3c179c4a_0a134981,
        64'hb53ff0ef_44818bb2,
        64'h8b2ee46e_e86aec66,
        64'he8caf0a2_f486f062,
        64'hf45ef85a_e4ceeca6,
        64'h02000513_8aaa6a05,
        64'hfc56e0d2_7159b751,
        64'h07a10585_80826161,
        64'h6ba26b42_6ae27a02,
        64'h79a27942_74e26406,
        64'h60a6557d_91afd0ef,
        64'h24050513_00003517,
        64'h926fd0ef_21450513,
        64'h00003517_058e02d6,
        64'h0b63fff7_c693c319,
        64'h86be8b05_63900085,
        64'h8733bf6d_07a10705,
        64'h6394e390_fff7c613,
        64'hc299863e_8a850087,
        64'h06b3a0a9_4501964f,
        64'hd0ef2aa5_05130000,
        64'h3517fd44_17e30405,
        64'h03259963_458187a6,
        64'h97efd0ef_855a85de,
        64'h986fd0ef_854e0327,
        64'h18634701_87a6994f,
        64'hd0ef8556_85de0004,
        64'h0b9b9a0f_d0ef854e,
        64'h4a41282b_0b130000,
        64'h3b1727aa_8a930000,
        64'h3a972729_89930000,
        64'h39979c0f_d0ef4401,
        64'h892ee45e_e486e85a,
        64'hec56f052_f44ef84a,
        64'he0a22825_05130000,
        64'h351784aa_fc26715d,
        64'hbf5d0785_a0019ecf,
        64'hd0ef2825_05130000,
        64'h351785a2_86269fcf,
        64'hd0ef26a5_05130000,
        64'h35176090_600c02e8,
        64'h03636098_00043803,
        64'h80826105_450164a2,
        64'h644260e2_00c79863,
        64'h00d50433_00d584b3,
        64'h00379693_4781e426,
        64'he822ec06_1101bbbf,
        64'hf06f8082_45018082,
        64'h45018082_80828082,
        64'h80824509_80824509,
        64'h80824509_bff92605,
        64'h20040413_6622dfff,
        64'hc0efe432_852285b2,
        64'h80826145_450164e2,
        64'h740270a2_00961863,
        64'h00c684bb_842ef406,
        64'hec26f022_71798082,
        64'h45058082_45058082,
        64'h45058082_01418d7d,
        64'h640260a2_95224080,
        64'h07b3f57f_f0efe406,
        64'h952e842a_e0221141,
        64'ha001cbbf_f0ef4505,
        64'habefd0ef_e4062f65,
        64'h05130000_351785aa,
        64'h862e86b2_87361141,
        64'h808202f5_553347a9,
        64'hb0002573_80824501,
        64'h80824501_80820141,
        64'h450160a2_eadfc0ef,
        64'h42000537_afafd0ef,
        64'he40630a5_05130000,
        64'h35171141_80828082,
        64'h61056442_60e28522,
        64'h936ff0ef_45816622,
        64'hc509842a_fd1ff0ef,
        64'he4328532_ec06e822,
        64'h110102b5_06338082,
        64'h953e055e_10d00513,
        64'he3089536_00178693,
        64'h00756513_157d631c,
        64'hdd070713_00004717,
        64'h80824501_80822405,
        64'h0513000f_4537a001,
        64'hd69ff0ef_e4062501,
        64'h11419002_00000023,
        64'hee1ff0ef_8522b781,
        64'h37050513_00003517,
        64'hc5112501_c87fa0ef,
        64'h4501fea5_85930000,
        64'h35974605_bfb93765,
        64'h05130000_3517c511,
        64'h2501b72f_b0efbfe5,
        64'h05130000_4517bb4f,
        64'hd06f0141_21c50513,
        64'h00003517_60a26402,
        64'h408005b3_cf81439c,
        64'he5c78793_00004797,
        64'h00054863_842a8bcf,
        64'h90efe607_a5230000,
        64'h4797e607_ab230000,
        64'h4797e985_05130000,
        64'h0517bf8f_d0ef2465,
        64'h05130000_3517b7e1,
        64'h3c850513_00003517,
        64'hc5112501_d69fa0ef,
        64'hc6850513_00004517,
        64'h3d058593_00003597,
        64'h4605c28f_d0ef3be5,
        64'h05130000_3517c34f,
        64'hd06f0141_60a26402,
        64'h3b050513_00003517,
        64'hc9112501_d47fa0ef,
        64'he022e406_ee450513,
        64'h00004517_0b458593,
        64'h00003597_46051141,
        64'h83020141_d7c58593,
        64'h00002597_60a26402,
        64'h8322f140_25730ff0,
        64'h000f0000_100fc84f,
        64'hd0efe406_3cc50513,
        64'h00003517_842a85aa,
        64'he0221141_bf95f287,
        64'ha3230000_47979c25,
        64'hbf5d2f40_10ef854e,
        64'hde7ff0ef_00094503,
        64'h993e0039_79133f67,
        64'h87930000_37970009,
        64'h099b00c4_591be05f,
        64'hf0ef4521_b775f6f7,
        64'h21230000_47174785,
        64'hcdefd0ef_3fc50513,
        64'h00003517_85a60496,
        64'h75634632_f8a7a023,
        64'h00004797_c50d2501,
        64'hfe3fa0ef_d5450513,
        64'h00004517_85ca8626,
        64'h0074f8f7_2d230000,
        64'h471757fd_80826121,
        64'h69e27902_74a27442,
        64'h70e2faa7_ab230000,
        64'h4797c10d_2501f08f,
        64'hb0efd8a5_05130000,
        64'h451702b7_856384b2,
        64'h842e892a_ec4efc06,
        64'hf04af426_f8227139,
        64'h439cfe27_87930000,
        64'h47978082_610560e2,
        64'he9fff0ef_00914503,
        64'hea7ff0ef_00814503,
        64'hf13ff0ef_ec06002c,
        64'h11018082_61456942,
        64'h64e27402_70a2fe94,
        64'h10e3ec9f_f0ef0091,
        64'h4503ed1f_f0ef3461,
        64'h00814503_f3fff0ef,
        64'h0ff57513_002c0089,
        64'h553354e1_03800413,
        64'h892af406_e84aec26,
        64'hf0227179_80826145,
        64'h694264e2_740270a2,
        64'hfe9410e3_f0bff0ef,
        64'h00914503_f13ff0ef,
        64'h34610081_4503f81f,
        64'hf0ef0ff5_7513002c,
        64'h0089553b_54e14461,
        64'h892af406_e84aec26,
        64'hf0227179_80826105,
        64'h644260e2_f43ff0ef,
        64'h00914503_f4bff0ef,
        64'h00814503_fb7ff0ef,
        64'h0ff47513_002cf5df,
        64'hf0ef0091_4503f65f,
        64'hf0ef0081_4503fd1f,
        64'hf0efec06_8121842a,
        64'h002ce822_11018082,
        64'h00f58023_00e580a3,
        64'h0007c783_00074703,
        64'h97aa973e_811100f5,
        64'h7713f1a7_87930000,
        64'h2797b7f5_0405fa5f,
        64'hf0ef8082_01416402,
        64'h60a2e509_00044503,
        64'h842ae406_e0221141,
        64'h808200e7_88230200,
        64'h071300e7_8423fc70,
        64'h071300e7_8623470d,
        64'h00078223_00e78023,
        64'h476d00e7_8623f800,
        64'h07130007_82234100,
        64'h07b78082_00a70023,
        64'hdfe50207_f7930147,
        64'h47834100_07378082,
        64'h02057513_0147c503,
        64'h410007b7_80820005,
        64'h45038082_00b50023,
        64'h80826105_690264a2,
        64'h644260e2_f47dfa1f,
        64'hf0ef4124_0433854a,
        64'h89260084_f3638922,
        64'h68048493_842ae04a,
        64'hec06e822_009894b7,
        64'he4261101_80826105,
        64'h690264a2_644260e2,
        64'hfe856ee3_f45ff0ef,
        64'h0405944a_02855433,
        64'h24040413_000f4437,
        64'h02a48533_3e2000ef,
        64'h892af63f_f0ef84aa,
        64'he04ae426_e822ec06,
        64'h11018082_02a7d533,
        64'h01419101_15026402,
        64'h60a202f4_07b32407,
        64'h8793000f_47b74140,
        64'h00ef842a_f95ff0ef,
        64'he022e406_11418082,
        64'h610564a2_8d0502a7,
        64'hd5336442_60e29101,
        64'h150202f4_07b33e80,
        64'h07934400_00ef842a,
        64'hfc1ff0ef_84aae426,
        64'he822ec06_11018082,
        64'h45018082_01418d5d,
        64'h91011782_150260a2,
        64'h1007e783_10a7a223,
        64'h10e1a023_27051001,
        64'ha70300e5_7763878e,
        64'h1041e703_504000ef,
        64'he4061141_8082cf1f,
        64'hf06fe225_85930000,
        64'h45974611_cb8103a7,
        64'hd7830000_47978082,
        64'h24010113_22013903,
        64'h22813483_23013403,
        64'h23813083_f63ff0ef,
        64'h8522002c_e90ff0ef,
        64'he802c44a_08282040,
        64'h061385a6_e52ff0ef,
        64'h22113c23_00282180,
        64'h06134581_893284ae,
        64'h842a2321_30232291,
        64'h34232281_3823dc01,
        64'h0113ebff_f06f6145,
        64'h05c170a2_41907402,
        64'hd8bff06f_614570a2,
        64'h65a27402_8522875f,
        64'hd0efe42e_75c50513,
        64'h00003517_842a885f,
        64'hd06f6145_78450513,
        64'h00003517_70a27402,
        64'h02f70a63_478d00d7,
        64'h0e6301e1_570300e1,
        64'h0f230115_c70300e1,
        64'h0fa34689_0105c703,
        64'hf022f406_71798082,
        64'h61056902_64a26442,
        64'h60e2d47f_f06f6105,
        64'h690264a2_60e26442,
        64'h8d7fd0ef_7a450513,
        64'h00003517_0087cf63,
        64'h278d439c_12478793,
        64'h00004797_12f71823,
        64'h00004717_27850007,
        64'hd78313e7_87930000,
        64'h47972400_00ef0200,
        64'h0513d19f_f0ef4515,
        64'h1545d583_00004597,
        64'h256000ef_4535e29f,
        64'hf0ef854a_f5c58593,
        64'h00004597_f6a79323,
        64'h00004797_4611cf3f,
        64'hf0ef17e5_55030000,
        64'h4517f6a7_9d230000,
        64'h4797d07f_f0ef4511,
        64'hda9ff0ef_00448513,
        64'hffc4059b_06a79a63,
        64'h25010024_d783d23f,
        64'hf0ef1ae5_55030000,
        64'h451708a7_95632501,
        64'h0004d783_d39ff0ef,
        64'h84ae450d_892a08c7,
        64'hdf638432_478de04a,
        64'he426ec06_e8221101,
        64'hb7911cf7_1f230000,
        64'h47174785_eafff0ef,
        64'h854efe25_85930000,
        64'h45974611_fea79723,
        64'h00004797_d79ff0ef,
        64'h4501fea7_9d230000,
        64'h4797d87f_f0ef20f7,
        64'h3f230000_471720f7,
        64'h3f230000_47174511,
        64'h07e20810_07939edf,
        64'hd0ef89a5_05130000,
        64'h4517858a_43902367,
        64'h87930000_4797decf,
        64'hf0ef850a_85a2df4f,
        64'hf0ef850a_8b458593,
        64'h00004597_00f70963,
        64'h02f00793_01294703,
        64'hde0ff0ef_850a6865,
        64'h85930000_3597855f,
        64'hf0ef850a_45811000,
        64'h0613b755_26f72e23,
        64'h00004717_20000793,
        64'h80826155_69b26952,
        64'h64f27412_70b2a5df,
        64'hd0ef8e25_05130000,
        64'h451700a4_05b3f1cf,
        64'hf0ef6ca5_05130000,
        64'h3517842a_f2aff0ef,
        64'h852204a7_f2630ff0,
        64'h07939526_f3aff0ef,
        64'h6e850513_00003517,
        64'h84aaf48f_f0ef8522,
        64'h2ca7ac23_00004797,
        64'h04e7ee63_1ff00793,
        64'hfff5071b_e93ff0ef,
        64'h95260505_f6aff0ef,
        64'h852600a4_04b30505,
        64'hf76ff0ef_892eea4a,
        64'hee26f606_852289aa,
        64'he64e0125_8413f222,
        64'h71698082_45018082,
        64'h01416402_60a28522,
        64'h547d0085_0363822f,
        64'ha0ef8432_e406e022,
        64'h114166a0_006f6105,
        64'h64a260e2_6442b0df,
        64'hd06f6105_97450513,
        64'h00004517_40a005b3,
        64'h64a260e2_64420005,
        64'h5e63809f_90efef85,
        64'h05130000_0517b35f,
        64'hd0ef9825_05130000,
        64'h4517b41f_d0ef9765,
        64'h05130000_45178622,
        64'h86aa608c_e2dfc0ef,
        64'h85a26088_b5bfd0ef,
        64'h85a29c11_ec0697e5,
        64'h05130000_45176380,
        64'he8226090_3b448493,
        64'h00004497_e4263c67,
        64'h87930000_47971101,
        64'h80826105_64a26442,
        64'he00c95a6_60e2600c,
        64'ha05ff0ef_ec066008,
        64'h85aa84ae_862ee426,
        64'h3f040413_00004417,
        64'he8221101_80823ef7,
        64'h3f230000_47173ef7,
        64'h3f230000_471707e2,
        64'h08100793_5020006f,
        64'h03050513_014160a2,
        64'h640202a4_753b4529,
        64'hfe7ff0ef_357d02b4,
        64'h55bb45a9_00b7f863,
        64'h47a500a0_4563842e,
        64'he406e022_1141b7c5,
        64'h0505fd07_879b9fb9,
        64'h02f607bb_00b6e763,
        64'hfd07059b_27018082,
        64'h853ee319_00054703,
        64'h462946a5_4781a93f,
        64'hf06f95be_92011602,
        64'h91811582_639c4767,
        64'h87930000_47978082,
        64'h01419141_15421141,
        64'h8d5d0522_0085579b,
        64'hfa5ff06f_4581d7df,
        64'hf06f0141_05054581,
        64'h462960a2_6402f77d,
        64'h8b110007_4703973e,
        64'h00054703_fea47ae3,
        64'h157d8082_0141557d,
        64'h640260a2_e7198b11,
        64'h00074703_973efff5,
        64'h8513fe27_87930000,
        64'h2797fff5_c70300a4,
        64'h05b3951f_f0efe589,
        64'h842ae406_e0221141,
        64'hbfd50789_bff1052a,
        64'h052ab7e9_e01c078d,
        64'h00e69863_04200713,
        64'h0027c683_fce69fe3,
        64'h052a0690_07130017,
        64'hc683fed7_16e306b0,
        64'h069302d7_076304d0,
        64'h06938082_01416402,
        64'h60a202d7_0e630470,
        64'h069300e6_ea6302d7,
        64'h04630007_c70304b0,
        64'h0693601c_f87ff0ef,
        64'h842ee406_e0221141,
        64'hb7e1e008_b7cdfc97,
        64'h879b0ff7_f793fe07,
        64'h079bc609_8a09b7d1,
        64'h96be0505_02d586b3,
        64'hfeb7f4e3_fd07879b,
        64'h00088b63_00467893,
        64'h80826105_85366442,
        64'h60e2ec05_00089863,
        64'h04467893_00064603,
        64'h00f80633_0007079b,
        64'h00054703_0bc80813,
        64'h00002817_468100c1,
        64'h6583e0df_f0efc632,
        64'hec06006c_842ee822,
        64'h1101bfd5_0789bff1,
        64'h052a052a_b7e9e01c,
        64'h078d00e6_98630420,
        64'h07130027_c683fce6,
        64'h9fe3052a_06900713,
        64'h0017c683_fed716e3,
        64'h06b00693_02d70763,
        64'h04d00693_80820141,
        64'h640260a2_02d70e63,
        64'h04700693_00e6ea63,
        64'h02d70463_0007c703,
        64'h04b00693_601cf0df,
        64'hf0ef842e_e406e022,
        64'h11418082_014140a0,
        64'h053360a2_f23ff0ef,
        64'he4060505_1141f2df,
        64'hf06f00e6_846302d0,
        64'h07130005_4683b7e9,
        64'h4501e088_fcf718e3,
        64'h47a9fd27_9be30785,
        64'h8f81cb01_0007c703,
        64'hfe8782e3_67e2f5df,
        64'hf0ef8522_082c892a,
        64'h862e8082_61217902,
        64'h74a27442_70e25529,
        64'he90165a2_b03ff0ef,
        64'h84b2842a_e42e0006,
        64'h3023f04a_fc06f426,
        64'hf8227139_b7e1e008,
        64'hb7cdfc97_879b0ff7,
        64'hf793fe07_079bc609,
        64'h8a09b7d1_96be0505,
        64'h02d586b3_feb7f4e3,
        64'hfd07879b_00088b63,
        64'h00467893_80826105,
        64'h85366442_60e2ec05,
        64'h00089863_04467893,
        64'h00064603_00f80633,
        64'h0007079b_00054703,
        64'h21080813_00002817,
        64'h468100c1_6583f61f,
        64'hf0efc632_ec06006c,
        64'h842ee822_11018082,
        64'hfae78fe3_4741bfed,
        64'h47a98082_c19c47a1,
        64'ha8090509_00e79c63,
        64'h07800713_0ff7f793,
        64'h0207879b_c7098b05,
        64'h00074703_973e25e7,
        64'h07130000_27170015,
        64'h478302f7_1f630300,
        64'h07930005_4703c19c,
        64'h47c1cf95_0447f793,
        64'h0007c783_97ba0025,
        64'h470304d7_17630780,
        64'h06930ff7_77130207,
        64'h071bc689_8a850006,
        64'hc68300e7_86b32a67,
        64'h87930000_27970015,
        64'h470306f7_1e630300,
        64'h07930005_4703e7c9,
        64'h419cb7f1_377d87aa,
        64'hbfa5fef5_1be30785,
        64'hf8b712e3_0007c703,
        64'h00d80a63_00878513,
        64'h0007b803_bfcd367d,
        64'h0785f8b7_1fe30007,
        64'hc703d24d_8a1deb11,
        64'h87aa2701_8edd0036,
        64'h57130207_96938fd9,
        64'h01071793_00b7e733,
        64'h00859793_8e19953a,
        64'h93011702_fed819e3,
        64'h0007869b_0785fcb6,
        64'h9de30007_c68387aa,
        64'h00a7083b_9f1d4721,
        64'hc39d0075_7793b7f5,
        64'h367d0785_feb71ce3,
        64'h0007c703_8082853e,
        64'h4781e601_87aa2601,
        64'h00c7ef63_0ff5f593,
        64'h47c1b7ed_853efeb7,
        64'h0be30015_07930005,
        64'h47038082_450100c5,
        64'h14630ff5_f593962a,
        64'hbfe10405_d17df83f,
        64'hf0ef8522_85ca8626,
        64'h80826145_69a26942,
        64'h64e27402_70a28522,
        64'h44010097_db634089,
        64'h87bb0085_09bbd0df,
        64'hf0ef8522_c8990005,
        64'h049bd19f_f0ef892e,
        64'he44ef406_e84aec26,
        64'h852e842a_f0227179,
        64'hbfc50505_feb78de3,
        64'h00054783_808200c5,
        64'h1363962a_8082853e,
        64'hd3f59f95_07050006,
        64'hc6830007_c78300e5,
        64'h86b300e5_07b3a821,
        64'h478100e6_14634701,
        64'hb7e500b7_00239722,
        64'h0005c583_00e685b3,
        64'h00f80733_fef605e3,
        64'h17fd4781_fff64613,
        64'h86ae8832_80820141,
        64'h640260a2_8522f53f,
        64'hf0ef00a5_e963842a,
        64'he406e022_11418082,
        64'h614564e2_69428526,
        64'h740270a2_00040023,
        64'hf75ff0ef_944a864a,
        64'h8522fff6_091300c5,
        64'h64636582_892ace11,
        64'h84aa6622_dd3ff0ef,
        64'he02ee84a_f406e432,
        64'hec26852e_842af022,
        64'h7179b7e5_01068023,
        64'h078500f7_06b30006,
        64'hc80300f5_86b38082,
        64'h00f61363_478100f5,
        64'h0733963a_95be078e,
        64'h02e78733_57610036,
        64'h5793fed7_65e340f6,
        64'h06b30106_b02307a1,
        64'h00f506b3_0006b803,
        64'h00f586b3_a811471d,
        64'h4781eb9d_872a8b9d,
        64'h00b567b3_04b50463,
        64'hb7f5feb7_8fa30785,
        64'hbfe9fee7_bc2307a1,
        64'h808200c7_9763963e,
        64'h963a97aa_078e02e7,
        64'h87335761_00365793,
        64'h0106ee63_40f88833,
        64'h469d00c5_08b387aa,
        64'hffed8f55_37fd0722,
        64'h0ff5f693_47a1eb05,
        64'h87aa0075_77138082,
        64'h4501b7e5_078900d7,
        64'h80a300e7_80238082,
        64'he3110017_c703ce81,
        64'h0007c683_87aacf99,
        64'h00054783_c11d8082,
        64'h610564a2_85266442,
        64'h60e2e008_05050005,
        64'h0023c501_f73ff0ef,
        64'h8526842a_c891e822,
        64'hec066104_e4261101,
        64'hbfd986a7_b1230000,
        64'h57970505_00050023,
        64'hc7810005_4783c519,
        64'hf9fff0ef_852285a6,
        64'h80826105_64a26442,
        64'h60e28522_44018807,
        64'hb7230000_5797ef81,
        64'h00044783_942afa1f,
        64'hf0ef85a6_8522cc11,
        64'h63808aa7_87930000,
        64'h5797e519_842a84ae,
        64'hec06e426_e8221101,
        64'hbfd587ae_b7e50505,
        64'hfafd0007_c6830785,
        64'hfee68fe3_80824501,
        64'heb190005_4703b7c5,
        64'h07858082_853efa7d,
        64'h00074603_070500d6,
        64'h0863a021_872eca89,
        64'h00074683_00f50733,
        64'h4781bfd5_872eb7d5,
        64'h0785fa7d_00074603,
        64'h0705fed6_0ee38082,
        64'h853eea99_00074683,
        64'h00f50733_4781b7fd,
        64'h07858082_40a78533,
        64'he7010007_c70300b7,
        64'h856387aa_95aa8082,
        64'h61056442_60e24501,
        64'hfe857be3_157d00b7,
        64'h86630005_47830ff5,
        64'hf5939522_65a2fe5f,
        64'hf0efec06_842ae42e,
        64'he8221101_bfcd0785,
        64'h808240a7_8533e701,
        64'h0007c703_87aabfcd,
        64'h0505dffd_808200b7,
        64'h93630005_47830ff5,
        64'hf5938082_4501bfcd,
        64'h0505c399_808200b7,
        64'h93630005_47830ff5,
        64'hf5938082_853efee1,
        64'h0705e399_4187d79b,
        64'h0187979b_40f687bb,
        64'h0007c783_00e587b3,
        64'h0007c683_00e507b3,
        64'ha0154781_00e61463,
        64'h47018082_853ef37d,
        64'h0505e399_4187d79b,
        64'h0187979b_40f707bb,
        64'hfff5c783_00054703,
        64'h05858082_00078023,
        64'hfec799e3_d375fee7,
        64'h8fa30785_fff5c703,
        64'h0585963e_fb7d0017,
        64'h86930007_c70387b6,
        64'h8082e219_87aab7d5,
        64'h87b68082_fb75fee7,
        64'h8fa30785_fff5c703,
        64'h0585eb09_00178693,
        64'h0007c703_87aa8082,
        64'hf76d00e6_80230785,
        64'h00f506b3_00074703,
        64'h00f58733_00c78c63,
        64'h47818082_fb75fee7,
        64'h8fa30785_fff5c703,
        64'h058587aa_80820141,
        64'h640260a2_8d411502,
        64'h9001fd1f_f0ef1402,
        64'h0005041b_fdbff0ef,
        64'he022e406_11418082,
        64'h01412501_640260a2,
        64'h8d410105_151bfe9f,
        64'hf0ef842a_fefff0ef,
        64'he022e406_1141fc3f,
        64'hf06faaa5_05130000,
        64'h55178082_25018d5d,
        64'h00f717bb_40f007bb,
        64'h00f7553b_93ed836d,
        64'h8f3d0127_d713e118,
        64'h97360017_671302d7,
        64'h86b36518_6294611c,
        64'h88068693_00005697,
        64'h1c60106f_80826105,
        64'h690264a2_644260e2,
        64'h8522e99f_f0ef10f4,
        64'h00230247_c7838522,
        64'h0ea42e23_681c18f4,
        64'h34232b87_87930000,
        64'h179718f4_30232c87,
        64'h87930000_179716f4,
        64'h3c238fa7_8793ffff,
        64'hf797e65f_f0ef0405,
        64'h28230325_3023e904,
        64'h10f502a3_47850ef5,
        64'h2c234799_c57c57fd,
        64'hcd21842a_20a010ef,
        64'h45051c00_059384aa,
        64'h892ec7ad_639cc7bd,
        64'h651ccbad_511ccbbd,
        64'h4d5ccfad_44014d1c,
        64'hc1414401_e04ae426,
        64'hec06e822_1101b771,
        64'h60003340_10ef9665,
        64'h05130000_451701a9,
        64'h8863d80f_e0ef8566,
        64'h85e20097_8e63601c,
        64'hd8efe0ef_855e85ca,
        64'h00090663_d9afe0ef,
        64'h638c855a_0fc42603,
        64'h681c8956_0007c363,
        64'h89524c1c_c7914901,
        64'h541cdb8f_e06f6125,
        64'h54850513_00004517,
        64'h6d026ca2_6c426be2,
        64'h7b027aa2_7a4279e2,
        64'h690664a6_60e66446,
        64'h02941563_4d299dec,
        64'h8c930000_4c970005,
        64'h0c1b3fab_8b930000,
        64'h4b973fab_0b130000,
        64'h4b173faa_8a930000,
        64'h4a973faa_0a130000,
        64'h4a1789aa_e0caec86,
        64'he06ae466_e862ec5e,
        64'hf05af456_f852fc4e,
        64'h6080e8a2_c3448493,
        64'h00005497_e4a6711d,
        64'h8082e308_e518e11c,
        64'he7886798_c4c78793,
        64'h00005797_e5088082,
        64'haa07a023_00005797,
        64'he79ce39c_c6478793,
        64'h00005797_b7d56000,
        64'ha8cff0ef_8522c781,
        64'h19a44783_80826105,
        64'h64a26442_60e20094,
        64'h176384be_ec06e426,
        64'h6380e822_c9478793,
        64'h00005797_11018082,
        64'h4388aea7_87930000,
        64'h57978082_0f850513,
        64'h8082c398_0015071b,
        64'h4388b027_87930000,
        64'h5797bfd5_55358082,
        64'h610564a2_644260e2,
        64'he0800f84_0413e501,
        64'hce0ff0ef_842acd09,
        64'hf7dff0ef_84aee822,
        64'hec06e426_1101bfcd,
        64'hf8400513_bfe54501,
        64'h80826105_60e25535,
        64'he97fe06f_610560e2,
        64'h00f70c63_0ff00793,
        64'h08154703_02b70063,
        64'h65a21035_4703c105,
        64'hfbdff0ef_e42eec06,
        64'h11014148_8082853e,
        64'hbfd187b6_00a60463,
        64'h0fc7a603_80820141,
        64'h853e4781_60a2f3cf,
        64'he0efe406_51450513,
        64'h00004517_85aa1141,
        64'h02e79063_6394631c,
        64'hd6070713_00005717,
        64'h80824501_80820141,
        64'h45016402_60a20dc0,
        64'h00ef13e0_00ef02c0,
        64'h0513fc5f_f0ef8522,
        64'h00055563_ac0fe0ef,
        64'h852212a0_00efd8f7,
        64'h29230000_5717842a,
        64'he406e022_47851141,
        64'hef9d439c_da878793,
        64'h00005797_808218b5,
        64'h0d238082_557d8082,
        64'h557d8082_4501c56c,
        64'h8702972a_4318972a,
        64'h8379eea5_05130000,
        64'h35171702_ef056863,
        64'h450d0007_081b377d,
        64'h8b3d01a6_571bf0e5,
        64'h1c634000_073706bb,
        64'ha42306db_a22306fb,
        64'ha02304cb_ae23018b,
        64'ha50345e6_46d647c6,
        64'h4636e805_1763842a,
        64'h90ffe0ef_c4be855e,
        64'h0107979b_008c4601,
        64'h07cbd783_c2be479d,
        64'h04f11023_47a506fb,
        64'h9e2304e1_57830007,
        64'hd663018b_a783ec05,
        64'h1163842a_943fe0ef,
        64'hc2be47d5_855ec4be,
        64'h0107979b_008c4601,
        64'h07cbd783_04f11023,
        64'h478d6ce0_00ef06cb,
        64'h851300ec_4641ef2f,
        64'hf06ffa10_0413bf6d,
        64'h11872583_97528379,
        64'h02079713_fcfc65e3,
        64'h4581bfa1_d171d13f,
        64'he0ef855e_45850b70,
        64'h06130ff6_f693bb35,
        64'hf53d9d9f_e0ef855e,
        64'hc9aff0ef_855e4601,
        64'h18fbae23_08bba223,
        64'h0017b793_17ed088b,
        64'ha583ef8d_1afba823,
        64'h409ce79d_0046f793,
        64'h00892683_f14dfeff,
        64'he0ef855e_408c913f,
        64'he0ef855e_02ebaa23,
        64'h0017b713_41b787b3,
        64'h01a78663_471100d7,
        64'h89634721_400006b7,
        64'h00092783_bfa5fb99,
        64'h10e30931_941fe0ef,
        64'h855e035b_aa2308fb,
        64'ha223180b_ae231a0b,
        64'ha823088b_a783dabf,
        64'he0ef855e_45850b70,
        64'h06134681_c90ddbbf,
        64'he0ef855e_0fb6f693,
        64'h45850b70_06130089,
        64'h4683c3a1_27818ff9,
        64'h00f9f7b3_00092703,
        64'h40dc04f7_19630017,
        64'hb79317ed_00494703,
        64'h409c1000_0db72000,
        64'h0d3715a9_09130000,
        64'h3917bd21_97bfe0ef,
        64'h5e050513_00004517,
        64'hff6498e3_04a1eb99,
        64'h278100f9_f7b300fa,
        64'h97bb409c_1c0c8c93,
        64'h00003c97_4c2d18eb,
        64'h0b130000_3b174a85,
        64'h17848493_00003497,
        64'hdaaff0ef_2981855e,
        64'h00f9f9b3_4601088b,
        64'ha583044b_a783040b,
        64'ha983e6f7_69e34004,
        64'h07b704fb_a02300c7,
        64'he793040b_a783d7dd,
        64'h8b8504db_a0230106,
        64'he693040b_a68304db,
        64'ha0230216_869bc589,
        64'h00c7f593_cd910027,
        64'hf5931abb_a42303f7,
        64'hf5930c46_478304fb,
        64'ha0230016_879b7000,
        64'h06b7b129_6a450513,
        64'h00004517_e611b5f1,
        64'he225ecf7_69e34004,
        64'h07b700f7_78631a0b,
        64'hb6034004_07b704fb,
        64'ha0232785_100007b7,
        64'hb0cd02fb_a4234785,
        64'h00d010ef_8526a39f,
        64'he0ef8a3d_8abd0146,
        64'h561b0106_569b0624,
        64'h85137325_85930000,
        64'h4597074b_a603a59f,
        64'he0ef04d4_85137365,
        64'h85930000_45970186,
        64'hd69b0ff7_77130ff7,
        64'hf7930ff6_f8130106,
        64'hd71b0086_d79b06cb,
        64'hc603077b_c883070b,
        64'ha683a8df_e0effef5,
        64'h36230245_05137565,
        64'h85930000_459784aa,
        64'h06fbc603_074bd683,
        64'h07abd703_02c7d7b3,
        64'hed109201_0a8bb783,
        64'hd11c9fb9_071200e0,
        64'h37338f75_02071613,
        64'h76c19fb5_068e00d0,
        64'h36b38ef9_f0068693,
        64'hff0106b7_9fb5068a,
        64'h00d036b3_8ef90f06,
        64'h8693f0f0_f6b79fb5,
        64'h00f037b3_068600d0,
        64'h36b32781_8ef98ff9,
        64'hccc68693_aaa78793,
        64'hccccd6b7_aaaab7b7,
        64'h08cba703_00050623,
        64'h00051523_4a0000ef,
        64'h855e08fb_a82308fb,
        64'ha6232000_0793c799,
        64'h19cba783_1afbaa23,
        64'h1b0ba783_0adba223,
        64'h0afba023_02d606bb,
        64'h02f757bb_8a8d0106,
        64'hd69b02e6_073b3e80,
        64'h0613c305_03f77713,
        64'h0126d71b_c78d2781,
        64'h8fd18ff9_0186d61b,
        64'h17fd67c1_00cda683,
        64'h08fbae23_0087171b,
        64'h1487a783_97b6078a,
        64'h2e068693_00003697,
        64'h04d61c63_800306b7,
        64'h018ba603_00f6f863,
        64'h8bbd00c7_579b46a5,
        64'h008da703_fda59ee3,
        64'hfefd2e23_8fd98ff5,
        64'h8f510087_d79b8e69,
        64'h0087961b_8f510187,
        64'h971b0187_d61b0d11,
        64'h000d2783_f0068693,
        64'h00ff0537_040d0593,
        64'h66c1bf91_11872583,
        64'h97528379_02079713,
        64'hf6f762e3_4581472d,
        64'hb575def9_8be310bc,
        64'h099181df_f0ef855e,
        64'h84058593_4601180b,
        64'hae23096b_a2231afb,
        64'ha823017d_85b74785,
        64'hf3f537fd_670267a2,
        64'hc521d51f_e0efe03a,
        64'hc93ae556_e16ae43e,
        64'h855e110c_01100400,
        64'h07134791_d5028dea,
        64'hd33a0af1_1023fe0c,
        64'h7d1347b5_6702ed05,
        64'hd7ffe0ef_d53ee03a,
        64'hd33a855e_110c0107,
        64'h979b4601_475507cb,
        64'hd7830af1_10230370,
        64'h0793895f_f0ef855e,
        64'h460118fb_ae2308bb,
        64'ha2230017_b79317ed,
        64'h088ba583_efd91afb,
        64'ha823409c_09b79063,
        64'h8bbd010c_c783e541,
        64'hdcffe0ef_c93ee556,
        64'he166855e_110c0400,
        64'h07930110_d53e00fd,
        64'he7b317c1_2d818100,
        64'h07b7d33e_47d50af1,
        64'h10234799_4d850ae7,
        64'h9d63470d_00e78663,
        64'h4705409c_d41fe0ef,
        64'h855e02fb_aa23001d,
        64'h379340fd_0d331000,
        64'h07b700ed_08634791,
        64'h20000737_00ed0d63,
        64'h47a14000_07370e05,
        64'h19638daa_8bfff0ef,
        64'h855e0015_b59340bd,
        64'h05b31000_05b700fd,
        64'h08634591_200007b7,
        64'h00fd0d63_45a14000,
        64'h07b71207_8e632781,
        64'h01a7f7b3_00f977b3,
        64'h0009ad03_40dc840b,
        64'h0b1b0601_0993017d,
        64'h8b37bf01_04fba023,
        64'h0087e793_040ba783,
        64'hf20750e3_02e79713,
        64'h8fd58ff9_0087d79b,
        64'h0087969b_f0070713,
        64'h674144dc_fbe18b85,
        64'h83a54cdc_e6051de3,
        64'heb7fe0ef_dc3ef84a,
        64'hf426c556_855e010c,
        64'h04000793_1030c33e,
        64'h47d508f1_10234799,
        64'h02098863_39fd0905,
        64'h3ac54995_98811902,
        64'h01000ab7_0ff10493,
        64'h4905bfa9_80030737,
        64'hb7858002_07370007,
        64'h45630307_9713b7bd,
        64'ha007071b_80011737,
        64'hb949df40_0413e15f,
        64'he0efa7a5_05130000,
        64'h5517fef4_93e35ee7,
        64'h87930000_379704a1,
        64'hebc52781_00f977b3,
        64'h00e797bb_47854098,
        64'h0a8583f9_79130207,
        64'h9a934785_00f97933,
        64'hfe0c7c93_60c48493,
        64'h00003497_044ba783,
        64'hf0be0ff1_0c13040b,
        64'ha903639c_21c78793,
        64'h00005797_08f71363,
        64'h800107b7_018ba703,
        64'h04fba023_8fd92000,
        64'h0737040b_a7830007,
        64'h596302d7_971300eb,
        64'hac238001_073708d7,
        64'h0e634689_c7010927,
        64'h0d638b3d_0187d71b,
        64'h04ebac23_8f558f71,
        64'h8ecd0087_571b8de9,
        64'h0087159b_8ecd0187,
        64'h169b0187_559b40d8,
        64'h04fbaa23_27818fd5,
        64'h8ef1f007_06138fd1,
        64'h67410087_569b8e69,
        64'h8fd50087_161b0187,
        64'h179b0187_569b00ff,
        64'h05374098_bd798a9d,
        64'h938100f6_d69b1782,
        64'h8fd901e6_d71b8ff9,
        64'h0027979b_17716705,
        64'hb54508bb_a82300b5,
        64'h15bb89bd_0165d59b,
        64'hbd914004_0737bda9,
        64'h40030737_bd894002,
        64'h0737bb75_842afe09,
        64'h96e339fd_c529844f,
        64'hf0efd05a_ec56e826,
        64'h855e108c_08104b21,
        64'h0a854991_d48206f1,
        64'h10239881_02091a93,
        64'h03300793_0bf10493,
        64'h4905d2ca_ed05874f,
        64'hf0efd4be_d2ca855e,
        64'h0107979b_108c4601,
        64'h07cbd783_06f11023,
        64'h03700793_04fba023,
        64'h27891000_07b75407,
        64'h5963018b_a703e205,
        64'h15e3842a_ff3fe0ef,
        64'h855e00b5_45831130,
        64'h00ef855e_e40510e3,
        64'h842ac94f_f0ef855e,
        64'h08fb80a3_57fd08fb,
        64'haa234785_e4051ce3,
        64'h842a8d8f_f0efc4be,
        64'hc2ca855e_008c0107,
        64'h979b4601_495507cb,
        64'hd78304f1_1023479d,
        64'h8f6ff0ef_c282c4be,
        64'h04e11023_855e008c,
        64'h46010107_979b4711,
        64'h00e78e63_577d04cb,
        64'ha783c215_08fba823,
        64'h00e7f463_20000793,
        64'h090ba703_08fba623,
        64'h0107d463_20000793,
        64'h0afbb823_0e0bb023,
        64'h0c0bbc23_0c0bb823,
        64'h0c0bb423_0c0bb023,
        64'h0a0bbc23_030787b3,
        64'h00d797b3_26890785,
        64'h46a18fd9_0106d79b,
        64'h8f7d003f_07370107,
        64'h979b1407_0f6302cb,
        64'ha703090b_a8231408,
        64'hdd63090b_a62300e5,
        64'h183b8b3d_0107d71b,
        64'h08eba223_08eba423,
        64'h04cba823_180bae23,
        64'h1a0ba823_8a0500c7,
        64'hd61b02c7_073b018b,
        64'ha8834505_0f874703,
        64'h10862603_96529752,
        64'h060a8b3d_7f4a0a13,
        64'h00003a17_8a1d0036,
        64'h571b00eb_ac234007,
        64'h071b4001_0737a029,
        64'h2007071b_40010737,
        64'hbf0506fb_9e234785,
        64'h02fba623_8b8541e7,
        64'hd79b048b_a78300fb,
        64'hac234000_07b7bfe9,
        64'h1f1010ef_06400513,
        64'h08a96fe3_163010ef,
        64'h85260007_cc63048b,
        64'ha783f155_842ab1ef,
        64'hf0ef855e_45853e80,
        64'h09139081_02051493,
        64'h187010ef_4501afef,
        64'hf0ef855e_0407c163,
        64'h180b8c23_048ba783,
        64'h8082615d_6db66d56,
        64'h6cf67c16_7bb67b56,
        64'h7af66a1a_69ba695a,
        64'h64fa741a_70ba8522,
        64'hd55d842a_d99ff0ef,
        64'h855ea031_020ba423,
        64'hf4fd34fd_10050de3,
        64'h842aa88f_f0ef855e,
        64'h008c4601_4495cf81,
        64'h8b851b8b_a7831205,
        64'h0ae3842a_aa2ff0ef,
        64'hc482c2be_855e008c,
        64'h479d4601_04f11023,
        64'h4789e7b5_180b8ca3,
        64'h198bc783_c7b1199b,
        64'hc7832190_10ef4501,
        64'h8baae3b5_4401e6ee,
        64'heaeaeee6_f2e2f6de,
        64'hfadafed6_e352e74e,
        64'heb4aef26_f706f322,
        64'h7161551c_b58584aa,
        64'hb595fa10_04939fcf,
        64'hf0efe325_05130000,
        64'h5517d965_c04ff0ef,
        64'h85224585_bfd118f4,
        64'h0c234785_0007d663,
        64'h443ced09_c1cff0ef,
        64'h85224581_becff0ef,
        64'h852202f5_1f63f920,
        64'h0793b55d_18f40ca3,
        64'h47850604_1e23d45c,
        64'h8b8541e7_d79bc43c,
        64'hcc188001_073700e6,
        64'h85638002_07374c14,
        64'hbf4534b0_10ef3e80,
        64'h05130609_0863397d,
        64'h0007ca63_47b2ed1d,
        64'hb76ff0ef_8522858a,
        64'h4601c43e_0197e7b3,
        64'h01871563_c43e0177,
        64'hf7b3c25a_4bdc0151,
        64'h10234c18_681ce13d,
        64'hb9eff0ef_c402c252,
        64'h01311023_8522858a,
        64'h46014000_0cb78002,
        64'h0c3700ff_8bb74b05,
        64'h02900a93_4a550370,
        64'h09933e90_0913cc1c,
        64'h800207b7_00f71563,
        64'h0aa00793_00c14703,
        64'he911be0f_f0efc23e,
        64'hc43a8522_858a4601,
        64'h47d50aa0_0713e399,
        64'h1aa00713_8ff94bdc,
        64'h00ff8737_681c00f1,
        64'h102347a1_000505a3,
        64'h46d000ef_8522f149,
        64'h84aacdaf_f0ef8522,
        64'hf13ff0ef_85224581,
        64'h4601b5ef_f0ef8522,
        64'hd85c4785_08f42223,
        64'h1a042823_18042e23,
        64'h08842783_f94584aa,
        64'h97826b9c_679c8522,
        64'h681c43b0_10ef7d00,
        64'h0513b8ef_f0ef8522,
        64'h02042c23_02f40823,
        64'h47851af4_2c23478d,
        64'hf93ff0ef_f3e54481,
        64'h541c8082_61097ca2,
        64'h7c427be2_6b066aa6,
        64'h6a4669e6_74a67906,
        64'h85267446_70e6f850,
        64'h0493b98f_f0effb65,
        64'h05130000_55170204,
        64'h2423eb8d_6b9c679c,
        64'h681cc509_f07ff0ef,
        64'h842ac17c_8fd9f466,
        64'hf862fc5e_e0dae4d6,
        64'he8d2ecce_f0caf4a6,
        64'hfc86f8a2_070d4b9c,
        64'h71191000_0737691c,
        64'h80828082_c18ff06f,
        64'h02c50823_dd0c0007,
        64'h859b87ba_00d5f363,
        64'h0007069b_0007859b,
        64'h4f1887ae_00d5f363,
        64'h0007869b_4f5c6918,
        64'he215b7cd_c402fef4,
        64'h14e34785_80826121,
        64'h790274a2_744270e2,
        64'hd26ff0ef_8526858a,
        64'h4601c43e_478900f4,
        64'h1f634791_c24a00f1,
        64'h10234799_ed19d44f,
        64'hf0efc43e_c24a8526,
        64'h858a4601_0107979b,
        64'h4955842e_07c4d783,
        64'h00f11023_03700793,
        64'h04f59263_55294785,
        64'h00f58663_84aa4791,
        64'hf04af822_fc06f426,
        64'h71398082_01416402,
        64'h60a24505_83020141,
        64'h60a26402_85220003,
        64'h07630187_b303679c,
        64'h681c0005_5e63ffdf,
        64'he0ef842a_e406e022,
        64'h1141b325_842ab335,
        64'hdd79842a_941ff0ef,
        64'h85264585_0a700613,
        64'h86cab381_842a953f,
        64'hf0ef8526_458509b0,
        64'h06134685_01279b63,
        64'h0a79c783_d4fb0ee3,
        64'h4785ed19_971ff0ef,
        64'h85264585_09c00613,
        64'h86defdba_18e30c11,
        64'h0ffa7a13_2a0dffac,
        64'h90e30ffa_fa932ca1,
        64'h2a85e139_999ff0ef,
        64'h85260ff6_f6930196,
        64'hd6bb4585_8656000c,
        64'h26834c81_8ad209b0,
        64'h0d934d61_08f00a13,
        64'hff9a10e3_2a05e92d,
        64'h9c5ff0ef_85264585,
        64'h0ff67613_0ff6f693,
        64'hf8ca061b_00dad6bb,
        64'h003a169b_4c8dfdbd,
        64'h1fe32d05_e9458a2a,
        64'h9edff0ef_85264585,
        64'h0ff67613_0ff6f693,
        64'hf88d061b_00dcd6bb,
        64'h003d169b_4d914d01,
        64'h08f4aa23_00a7979b,
        64'h0e09c783_0af987a3,
        64'h4785e579_a21ff0ef,
        64'h85264585_0af00613,
        64'h4685e395_8b850af9,
        64'hc783e20b_05e3b535,
        64'h547ddb8f_f0ef1b65,
        64'h05130000_5517cb89,
        64'h8b8509b9_c783bfd1,
        64'h00f97933_fff7c793,
        64'hb5a939c0_20ef1865,
        64'h05130000_5517ef89,
        64'h8b850a69_c78302d9,
        64'h0263fcb6_14e387b2,
        64'h0ff97913_0127e933,
        64'hc70d4189_591b4187,
        64'hd79b8b05_0189191b,
        64'h0187979b_0027571b,
        64'h00c517bb_c39d8b85,
        64'h0017579b_4b9897d2,
        64'h078e0017_861b4591,
        64'h45054781_0016e913,
        64'hc3990fe6_f9138b89,
        64'hc7198936_0017f713,
        64'h0a79c683_008a4783,
        64'hb5c9e50f_f0ef1ce5,
        64'h05130000_551785ca,
        64'h01267a63_963e09d9,
        64'hc7839e3d_0087979b,
        64'h0106161b_09e9c783,
        64'h09f9c603_ee051ae3,
        64'h842af8af_f0ef8526,
        64'h85ceee06_8de31d65,
        64'h05130000_55178a89,
        64'h000b8963_fa6596e3,
        64'h87ae0611_05210128,
        64'h893b0ffb_fb9300fb,
        64'hebb300be_17bbcb89,
        64'h8b850107_c78397d2,
        64'h078e0208_00630116,
        64'h202302e8_58bbb7f1,
        64'h4b814a81_4c81b7c9,
        64'hed6ff0ef_1f450513,
        64'h00005517_00088d63,
        64'h02e878bb_0017859b,
        64'h00052803_43114e05,
        64'h47818956_866200ca,
        64'h05138c0a_009c9c9b,
        64'he3994b85_02eadabb,
        64'h54dcb761_5429f14f,
        64'hf0ef1fa5_05130000,
        64'h5517cb89_02ecf7bb,
        64'h0005ac83_e79102ea,
        64'hf7bb060a_8063fe09,
        64'hf99302f1_09930045,
        64'haa83db45_1fc50513,
        64'h00005517_0984a703,
        64'h80822a01_01132381,
        64'h3d832401_3d032481,
        64'h3c832501_3c032581,
        64'h3b832601_3b032681,
        64'h3a832701_3a032781,
        64'h39832801_39032881,
        64'h34832901_34032981,
        64'h30838522_f8400413,
        64'hf8eff0ef_22450513,
        64'h00005517_e7b90016,
        64'hf79307e4_c68300e7,
        64'heb632025_05130000,
        64'h55178a2e_8b3284aa,
        64'hbfe78793_3ffc07b7,
        64'h9f3dbff7_879bbffc,
        64'h07b74d18_0ac7ed63,
        64'h478923b1_3c2325a1,
        64'h30232591_34232581,
        64'h38232571_3c232761,
        64'h30232751_34232741,
        64'h38232731_3c232921,
        64'h30232891_34232881,
        64'h38232811_3c23d601,
        64'h01138082_614569a2,
        64'h694264e2_740270a2,
        64'h85220135_05a317a0,
        64'h10ef8526_842a86df,
        64'hf0ef8526_85ca0009,
        64'h1c6300f5_1e63842a,
        64'h57b5c519_cc1ff0ef,
        64'h84aa4585_0b300613,
        64'h8edd892e_9be10079,
        64'hf6930ff5_f9930815,
        64'h4783f022_f406e44e,
        64'he84aec26_7179bfd9,
        64'h84aab755_4685fef7,
        64'h60e354a9_4705ffc5,
        64'h879b8082_24010113,
        64'h22813483_22013903,
        64'h85262301_34032381,
        64'h3083df40_0493e399,
        64'h0b944783_e9159a7f,
        64'hf0ef854a_85a29801,
        64'h01f10413_ed912581,
        64'h99f5ffe4_059be11d,
        64'h84aad3ff_f0ef892a,
        64'h45850b90_0613842e,
        64'hed8554a9_468104b7,
        64'hec6306f5_84634789,
        64'h23213023_22913423,
        64'h22813823_22113c23,
        64'hdc010113_b7655929,
        64'hb7755951_bf451a04,
        64'hb0235f00_20efdd4d,
        64'h1a04b503_892ab75d,
        64'h08f4aa23_02f707bb,
        64'h27852705_8bfd8b7d,
        64'h0057d79b_00a7d71b,
        64'h50fcf3dd_8b850af4,
        64'h47838082_25010113,
        64'h22813983_23013903,
        64'h23813483_854a2401,
        64'h34032481_308308f4,
        64'h80230a74_478308f4,
        64'hac2300a7_979b02e7,
        64'h87bb0dd4_47030e04,
        64'h4783f8dc_07a60d44,
        64'h27830009_8663c799,
        64'h54dc08f4_aa2300a7,
        64'h979b0e04_47830af4,
        64'h07a34785_e141e0bf,
        64'hf0ef8526_45850af0,
        64'h06134685_c6b5e391,
        64'h8bfd09c4_4783c789,
        64'h8b850a04_4783f4fc,
        64'h07a6c319_f4fc54d8,
        64'h9fb90884_47039fb9,
        64'h0087171b_08944703,
        64'h9fb90107_171b0187,
        64'h979b08a4_470308b4,
        64'h4783f8fc_07ce02e7,
        64'h87b30dd4_478302f7,
        64'h07330e04_470397ba,
        64'h08c44703_9fb90087,
        64'h171b0107_979b4685,
        64'h08d44703_08e44783,
        64'h04098f63_fce514e3,
        64'h0621070d_e21c07ce,
        64'h02b787b3_0dd44783,
        64'h02f585b3_0e044583,
        64'h00098c63_4685c391,
        64'h97aeffe7_45839fad,
        64'h0105959b_0087979b,
        64'h00074583_fff74783,
        64'he0fc07c6_468109d4,
        64'h05130a84_4783fcdc,
        64'h07c60c84_86130914,
        64'h07130e24_478306f4,
        64'h8fa309c4_4783c789,
        64'h8b890a04_47830009,
        64'h8a6308f4_80a30b34,
        64'h4783c789_0e244783,
        64'he7810019_f9938b85,
        64'h06f48f23_09b44983,
        64'h0a044783_f8dc00d7,
        64'h73630147_d69307a6,
        64'h80070713_67050d44,
        64'h278300e7_fd63cc98,
        64'h1ff78793_400407b7,
        64'h53b897ba_078a1ee7,
        64'h07130000_47171cf7,
        64'h6d634721_0c044783,
        64'h13d010ef_85a22000,
        64'h06131e05_05631a04,
        64'hb5031aa4_b0237920,
        64'h20ef2000_0513e799,
        64'h1a04b783_1e051a63,
        64'h892ac03f_f0ef84aa,
        64'h85a29801_01f10413,
        64'h1ce7f363_49013ffc,
        64'h07372331_34232291,
        64'h3c232481_30232411,
        64'h34239fb9_23213823,
        64'hbffc07b7_db010113,
        64'h4d18bfcd_fc79347d,
        64'h80826121_74a27442,
        64'h70e2d8bf_f0ef8526,
        64'h3e800593_e919c4df,
        64'hf0ef8526_858a4601,
        64'h440dc432_c23e84aa,
        64'hfc06f426_f82247f5,
        64'h8e5500f1_10230300,
        64'h06b78e55_47997139,
        64'h0106161b_0086969b,
        64'h80826121_6aa26a42,
        64'h69e274a2_79028526,
        64'h744270e2_fc0999e3,
        64'h9aa20287_84339a22,
        64'h408989b3_08c96783,
        64'hfc851ae3_f01ff0ef,
        64'h854a85d6_865286a2,
        64'h844e0089_f3630207,
        64'he4030109_378389a6,
        64'hf96decdf_f0ef854a,
        64'h08c92583_a0894481,
        64'hbd7ff0ef_60450513,
        64'h00005517_00b67a63,
        64'h014485b3_68100005,
        64'h4d638b3f_a0ef8522,
        64'h00b44583_c11d892a,
        64'h4a4010ef_8ab684b2,
        64'h8a2e4148_842ace05,
        64'he456e852_ec4ef04a,
        64'hf426f822_fc067139,
        64'hb7c54401_b7d50004,
        64'h841bb74d_02f6063b,
        64'hbf6147c5_80826125,
        64'h690664a6_644660e6,
        64'h8522c41f_f0ef64e5,
        64'h05130000_5517c11d,
        64'hd4fff0ef_d23ed402,
        64'h854a100c_47f54601,
        64'h02f11023_47b10497,
        64'hf0634785_e529842a,
        64'hd6fff0ef_c83eca26,
        64'hd23a854a_100c4785,
        64'h0030cc3e_e42e4755,
        64'hd432cf31_08c92783,
        64'h260102f1_102302c9,
        64'h270347c9_06d7f663,
        64'h84b6892a_4785e8a2,
        64'hec86e0ca_e4a6711d,
        64'h80824501_bfd54501,
        64'h80826121_74a27442,
        64'h70e2f8ed_34fdc901,
        64'hdc7ff0ef_8522858a,
        64'h46014495_cb918b89,
        64'h1b842783_c11ddddf,
        64'hf0efc23e_842af426,
        64'hfc06f822_858a4601,
        64'h47d5c42e_00f11023,
        64'h47c17139_e7a919c5,
        64'h2783bf6d_f9200513,
        64'hd07ff0ef_6f450513,
        64'h00005517_fc8047e3,
        64'h45018456_b74d8456,
        64'h608020ef_3e800513,
        64'h00805863_fff40a9b,
        64'hfe04c5e3_34fd8082,
        64'h61257b02_7aa27a42,
        64'h79e26906_64a66446,
        64'h60e6fba0_0513d4df,
        64'hf0ef7225_05130000,
        64'h5517c795_0125f7b3,
        64'h05479563_0135f7b3,
        64'hc7891005_f79345b2,
        64'hed15e71f_f0ef855a,
        64'h858a4601_e00a0a13,
        64'he0098993_08090913,
        64'h4495c43e_842e8b2a,
        64'hf456ec86_f05ae4a6,
        64'he8a26a05_6989fdf9,
        64'h49370107_979bf852,
        64'hfc4ee0ca_07c55783,
        64'hc23e47d5_00f11023,
        64'h47b5711d_80826145,
        64'h740270a2_c43c47b2,
        64'he119ec9f_f0ef8522,
        64'h858a4601_c43e8fd9,
        64'h40000737_8fd98f75,
        64'h600006b7_8ff58ff9,
        64'hf8068693_4bdc0080,
        64'h06b74538_691cc195,
        64'h842ac402_c23ef406,
        64'hf0224785_00f11023,
        64'h47857179_80826145,
        64'h740270a2_85226fe0,
        64'h20ef7d00_0513e509,
        64'h842af21f_f0efc202,
        64'hc4020001_1023858a,
        64'h46018522_71c020ef,
        64'hf4063e80_0513842a,
        64'hf0227179_80824501,
        64'hbf654501_fd4559b0,
        64'h10ef0d44_85130d44,
        64'h05934611_fcf715e3,
        64'h0e044783_0e04c703,
        64'hfcf71be3_0c044783,
        64'h0c04c703_fef711e3,
        64'h0dd44783_0dd4c703,
        64'h80822401_01132281,
        64'h34832301_34032381,
        64'h3083fb60_051300f7,
        64'h0d630a04_47830a04,
        64'hc703e909_fadff0ef,
        64'h1a053483_22113c23,
        64'h22913423_85a29801,
        64'h01f10413_22813823,
        64'hdc010113_08e6e063,
        64'h40040737_4d148082,
        64'h616160a6_fd3ff0ef,
        64'hcc3ed402_e486100c,
        64'h20000793_0030e83e,
        64'he42e0785_17824785,
        64'hd23e47d5_02f11023,
        64'h47a1715d_83020007,
        64'hb303679c_691c8082,
        64'h8c850513_00006517,
        64'h80826108_953e8175,
        64'h64878793_00004797,
        64'h150200a7_eb6347ad,
        64'h8082557d_80820141,
        64'h640260a2_45018302,
        64'h014160a2_64028522,
        64'h00030763_0207b303,
        64'h679c681c_00055e63,
        64'hff5ff0ef_842ae406,
        64'he0221141_8082557d,
        64'h8082557d_b7f1659c,
        64'h95aa058e_05e135f1,
        64'hbfe1617c_bff17d5c,
        64'h80826105_45016442,
        64'he90064a2_60e20294,
        64'h54330e70_10ef9081,
        64'h14827540_f55c08c5,
        64'h2483795c_878297b6,
        64'he426e822_ec061101,
        64'h431c9736_00259713,
        64'h6b068693_00004697,
        64'h04b7ec63_479d8082,
        64'h45018302_00030363,
        64'h0087b303_679c691c,
        64'h80826135_645260f2,
        64'h85221570_20ef0808,
        64'h842ae3ff_f0efe436,
        64'heec6eac2_e6bee2ba,
        64'hea22ee06_08081000,
        64'h05931234_862afe36,
        64'hfa32f62e_710d8082,
        64'h616160e2_e69ff0ef,
        64'he436e4c6_e0c2fc3e,
        64'hf83aec06_10000593,
        64'h1014862e_f436f032,
        64'h715d8082_616160e2,
        64'he8dff0ef_e436e4c6,
        64'he0c2fc3e_f83aec06,
        64'h1034f436_715db7f1,
        64'h85220201_03930005,
        64'h059b5010_10ef8522,
        64'h01247433_60000084,
        64'h0b13b5fd_845ad89f,
        64'hf0ef0084_0b130201,
        64'h03930004_4503a809,
        64'hdd1ff0ef_00280201,
        64'h03930005_059be31f,
        64'hf0ef4008_45a94601,
        64'h0016b693_00380084,
        64'h0b13f8b5_0693a811,
        64'h45c10016_36134685,
        64'h00380084_0b13fa85,
        64'h0613f6e5_10e30780,
        64'h071302e5_00630750,
        64'h0713a00d_46014685,
        64'h00380084_0b13f6e5,
        64'h1ee30700_071300a7,
        64'h6c6306e5_0e630730,
        64'h0713b74d_048d0024,
        64'hc5038082_61090007,
        64'h051b6b06_6aa66a46,
        64'h69e67906_74a67446,
        64'h70e6f55d_08f50963,
        64'h06300793_04d50f63,
        64'h05800693_02a6eb63,
        64'h06d50f63_06400693,
        64'h04890014_c5034781,
        64'h00f6f363_46a50ff7,
        64'hf793fd07_879bcb9d,
        64'h0004c783_03551063,
        64'h47810489_05450f63,
        64'h0014c503_bfe1e71f,
        64'hf0ef0201_03930485,
        64'h01350863_04d7ff63,
        64'h93811782_76820017,
        64'h079bc52d_8f1d0004,
        64'hc50377a2_77420209,
        64'h59130300_0a9306c0,
        64'h0a130250_0993f82a,
        64'hf02ef42a_fc3e8436,
        64'h84b2e0da_fc86e4d6,
        64'he8d2ecce_f4a6f8a2,
        64'h597d011c_f0ca7119,
        64'hb7e10117_80230066,
        64'h00230685_00064883,
        64'h0007c303_00d70633,
        64'h97ba9381_178240f8,
        64'h07bbb7d1_feb50fa3,
        64'h0505bf45_00c8063b,
        64'h808200b7_ea630006,
        64'h879bfff5_081b4681,
        64'h0015559b_9d190005,
        64'h00230505_00f50023,
        64'h02d00793_00030763,
        64'h02f6e963_00a606bb,
        64'h03000593_40e0063b,
        64'h8536fcb8_ffe302b8,
        64'hd53bfec6_8fa30685,
        64'h0ff67613_0306061b,
        64'h04ae6a63_0ff57613,
        64'h02b8f53b_0005089b,
        64'h385986ba_4e250ff6,
        64'hf8130410_0693c219,
        64'h06100693_430540a0,
        64'h053be681_00055663,
        64'h4301bfd9_00d70023,
        64'h07850006_c68300f5,
        64'h06b300d3_b8230017,
        64'h06938082_852e0007,
        64'h002300b6_e6630103,
        64'hb7030007_869b4781,
        64'h9d9dfff7_059b00c6,
        64'hf5638e9d_fff70693,
        64'h0003b703_8f999201,
        64'h02059613_0103b783,
        64'h0083b703_80824501,
        64'h80820007_80234505,
        64'h0103b783_00a70023,
        64'h00f3b823_00170793,
        64'h00d7fe63_93811782,
        64'h278540f7_07b30003,
        64'hb6830083_b7830103,
        64'hb7038082_61454501,
        64'h6a0269a2_694264e2,
        64'h740270a2_2f2000ef,
        64'h28050513_00006517,
        64'hfd241de3_302000ef,
        64'h819100f5_f6130405,
        64'h854e0007_c5830084,
        64'h87b33180_00ef8552,
        64'he7810004_059b01f4,
        64'h77932000_0913cd69,
        64'h89930000_6997cd6a,
        64'h0a130000_6a174401,
        64'hed9ff0ef_85264581,
        64'h346000ef_cd450513,
        64'h00006517_fac60613,
        64'h00006617_e789c4e6,
        64'h06130000_6617584c,
        64'h19c42783_daffb0ef,
        64'h2f858593_00006597,
        64'h744813c0_30efcf65,
        64'h05130000_65173840,
        64'h00efcea5_05130000,
        64'h6517c725_85930000,
        64'h6597c789_c8458593,
        64'h00006597_545c3a40,
        64'h00efcfa5_05130000,
        64'h65175c0c_3b2000ef,
        64'h0186561b_0ff6f693,
        64'h0ff77713_0ff67793,
        64'h0106569b_0086571b,
        64'hd0850513_00006517,
        64'h06c44583_58303dc0,
        64'h00ef91c1_15c20085,
        64'hd59bd125_05130000,
        64'h6517546c_3f2000ef,
        64'hd0850513_00006517,
        64'h06f44583_402000ef,
        64'h638cd0a5_05130000,
        64'h6517681c_224010ef,
        64'h842a4bf0_10ef4501,
        64'h479010ef_0001b503,
        64'h1ea030ef_d2450513,
        64'h00006517_84aa0e20,
        64'h30efe052_e44ee84a,
        64'hec26f022_f4062000,
        64'h05137179_7a00006f,
        64'h61054685_60e26622,
        64'h644285a2_501010ef,
        64'he42eec06_4501842a,
        64'he8221101_80820141,
        64'h640260a2_557de391,
        64'h4505703c_1a8030ef,
        64'hcc050513_00006517,
        64'hcb058593_00006597,
        64'h34c00613_b5c68693,
        64'h00005697_02f40263,
        64'h420007b7_e4066380,
        64'he0221141_711c8082,
        64'h25016388_97aa4200,
        64'h07b7050e_f73ff06f,
        64'h42000537_45814609,
        64'h8082b7f9_c45c4785,
        64'hd8f14501_8885bfe9,
        64'h4501c45c_4789c789,
        64'h0024f793_f4040124,
        64'h2423e01c_420007b7,
        64'h80826145_69a26942,
        64'h64e27402_70a2557d,
        64'h1f6030ef_85220009,
        64'h9d635080_00efdce5,
        64'h05130000_65178622,
        64'h85aa89aa_7b3010ef,
        64'hbc050513_00005517,
        64'h85a2c41d_5551842a,
        64'h1dc030ef_892e84b2,
        64'he44ef406_e84aec26,
        64'hf0220480_05137179,
        64'h08b04163_5535b7dd,
        64'h87ca14e1_09a13c20,
        64'h20efe43e_002c4621,
        64'h854e639c_00878913,
        64'hdcd50109_64830009,
        64'h398397a6_67a1bf41,
        64'hb1bff0ef_8522b771,
        64'h00f92623_0009b783,
        64'hdbd98b85_bd856770,
        64'h20ef4505_d8098ce3,
        64'hc43ff0ef_8522484c,
        64'hc85c9bf5_4985485c,
        64'hb4bff0ef_8522ef8d,
        64'h8b850089_27830009,
        64'h09630404_30232ea0,
        64'h30ef855a_85d60ca0,
        64'h0613c526_86930000,
        64'h56970184_8c630404,
        64'h39036004_cc9d4985,
        64'h8889c85c_9bf9485c,
        64'hc85c0027_e793485c,
        64'hcbb5603c_feb690e3,
        64'h0791872a_2685c398,
        64'h8f518361_ff873703,
        64'h01068763_c3900086,
        64'h161bff87_05136310,
        64'h4591480d_468100c9,
        64'h07930189_871308e6,
        64'h9f630037_f693470d,
        64'h02043c23_00492783,
        64'hcba97c1c_368030ef,
        64'h855a85d6_09c00613,
        64'hcb868693_00005697,
        64'h01898c63_03843903,
        64'h00043983_cfb50014,
        64'hf7936600_00efefe5,
        64'h05130000_651785ca,
        64'hd1bff0ef_85ca2901,
        64'h00496913_ff397913,
        64'h85220144_2903c39d,
        64'h0084f793_68a000ef,
        64'hf0050513_00006517,
        64'h85cad45f_f0ef85ca,
        64'h29010089_6913ff39,
        64'h79138522_01442903,
        64'hc39d0044_f793b29f,
        64'hf0ef8522_4581b71f,
        64'hf0ef8522_4581cc5c,
        64'hf9200793_c7817c1c,
        64'h00f76f63_0c893783,
        64'h02093703_14048063,
        64'h24818cfd_4981485c,
        64'h07093483_418030ef,
        64'h855a85d6_0f200613,
        64'h86e60189_09630004,
        64'h3903b711_702000ef,
        64'hf6050513_00006517,
        64'hd5058593_00005597,
        64'h000b9d63_3bfd4200,
        64'h0c378bd2_bd6100c4,
        64'he493bd85_458030ef,
        64'hf7050513_00006517,
        64'hf6058593_00006597,
        64'h14900613_d6c68693,
        64'h00005697_b7654701,
        64'h47812585_e31c9746,
        64'h93818375_17821702,
        64'h00be873b_8fd98fe9,
        64'h01076733_0087d79b,
        64'h01c87833_0087981b,
        64'h01076733_0187971b,
        64'h0187d81b_f2e50067,
        64'h036316fd_06052781,
        64'h0107e7b3_01e8183b,
        64'h07050037_1f1b0006,
        64'h4803ec06_89e36e89,
        64'hf0050513_00ff0e37,
        64'h43114701_47814581,
        64'h63900107_e6836541,
        64'h00043883_603cee07,
        64'h9be38b85_449cdf5f,
        64'hf0ef8522_488cdb9f,
        64'hf0efe024_852244cc,
        64'h80826165_45016ce2,
        64'h7c027ba2_7b427ae2,
        64'h6a0669a6_694664e6,
        64'h740670a6_efe9485c,
        64'h040b0b13_00006b17,
        64'h030a8a93_00006a97,
        64'hebbff0ef_25810015,
        64'he593e7ac_8c930000,
        64'h5c978522_0d89b583,
        64'hcdbff0ef_85224585,
        64'he9bff0ef_85222405,
        64'h8593000f_45b7d31f,
        64'hf0ef8522_45814605,
        64'h46854705_cffff0ef,
        64'h85224581_cc7ff0ef,
        64'h852285a6_c8bff0ef,
        64'h681a0a13_85220009,
        64'h5583c55f_f0ef0098,
        64'h9a378522_00892583,
        64'hbe3ff0ef_85224581,
        64'hd73ff0ef_85224581,
        64'h46054681_47050144,
        64'he4931607_86638b85,
        64'h008a2783_000a0963,
        64'h8cdd0324_3c234c1c,
        64'h4485e391_448d8b89,
        64'hc7090017_f7134481,
        64'h00492783_16f99a63,
        64'h04043a03_420007b7,
        64'h00043983_bf7ff0ef,
        64'h45856008_0e049c63,
        64'h6f6020ef_00c90513,
        64'h45814611_d01ce030,
        64'h84b2892e_0005d783,
        64'h020408a3_ec66f062,
        64'hf45ef85a_fc56e0d2,
        64'he4cef486_e8caeca6,
        64'h7100f0a2_71598082,
        64'h61056902_64a26442,
        64'h60e2c844_04993c23,
        64'h64c030ef_16450513,
        64'h00006517_15458593,
        64'h00006597_07600613,
        64'hf5068693_00005697,
        64'h02f90263_84ae842a,
        64'h420007b7_ec06e426,
        64'he8220005_3903e04a,
        64'h11018082_610564a2,
        64'h644260e2_e4246920,
        64'h30ef1aa5_05130000,
        64'h651719a5_85930000,
        64'h659706f0_0613f866,
        64'h86930000_569702f4,
        64'h026384ae_420007b7,
        64'hec06e426_6100e822,
        64'h11018082_610564a2,
        64'h644260e2_e0a09051,
        64'h14526d60_30ef1ee5,
        64'h05130000_65171de5,
        64'h85930000_65970680,
        64'h0613fba6_86930000,
        64'h569702f4_8263842e,
        64'h420007b7_ec06e822,
        64'h6104e426_11018082,
        64'h610564a2_644260e2,
        64'hfc809041_144271a0,
        64'h30ef2325_05130000,
        64'h65172225_85930000,
        64'h65970610_0613fee6,
        64'h86930000_569702f4,
        64'h8263842e_420007b7,
        64'hec06e822_6104e426,
        64'h1101d4df_f06f0141,
        64'h458160a2_64026008,
        64'hf23ff0ef_46054685,
        64'h47054581_8522ef1f,
        64'hf0ef4581_8522f39f,
        64'hf0ef842a_45810405,
        64'h30230205_3c234605,
        64'h46814705_e022e406,
        64'h11418082_01414501,
        64'h640260a2_d97ff0ef,
        64'h45816008_f67ff0ef,
        64'h45814605_46854705,
        64'h8522f35f_f0ef4581,
        64'h8522f7df_f0efe406,
        64'h45818522_46054681,
        64'h47057100_e0221141,
        64'h80826121_69e27902,
        64'h74a27442_70e20289,
        64'hb8238c45_88a10124,
        64'h64330034_949b8c59,
        64'h00497913_0029191b,
        64'h8b058809_0014141b,
        64'h67227fe0_30efe43a,
        64'h31850513_00006517,
        64'h30858593_00006597,
        64'h05a00613_0c468693,
        64'h00005697_02f98463,
        64'h84368932_84ae4200,
        64'h07b7fc06_f04af426,
        64'hf8220005_3983ec4e,
        64'h71398082_610564a2,
        64'h644260e2_f40404b0,
        64'h30ef3625_05130000,
        64'h65173525_85930000,
        64'h65970530_06130fe6,
        64'h86930000_569702f4,
        64'h026384ae_420007b7,
        64'hec06e426_6100e822,
        64'h11018082_610564a2,
        64'h644260e2_f00408b0,
        64'h30ef3a25_05130000,
        64'h65173925_85930000,
        64'h659704c0_061312e6,
        64'h86930000_569702f4,
        64'h026384ae_420007b7,
        64'hec06e426_6100e822,
        64'h11018082_610564a2,
        64'h644260e2_ec809001,
        64'h14020cf0_30ef3e65,
        64'h05130000_65173d65,
        64'h85930000_65970450,
        64'h0613fc26_86930000,
        64'h769702f4_8263842e,
        64'h420007b7_ec06e822,
        64'h6104e426_11018082,
        64'h610564a2_644260e2,
        64'he8809001_14021130,
        64'h30ef42a5_05130000,
        64'h651741a5_85930000,
        64'h659703e0_061300e6,
        64'h86930000_769702f4,
        64'h8263842e_420007b7,
        64'hec06e822_6104e426,
        64'h11018082_610564a2,
        64'h644260e2_e4041530,
        64'h30ef46a5_05130000,
        64'h651745a5_85930000,
        64'h65970360_06131e66,
        64'h86930000_569702f4,
        64'h026384ae_420007b7,
        64'hec06e426_6100e822,
        64'h11018082_610564a2,
        64'h644260e2_e0041930,
        64'h30ef4aa5_05130000,
        64'h651749a5_85930000,
        64'h659702f0_06132166,
        64'h86930000_569702f4,
        64'h026384ae_420007b7,
        64'hec06e426_6100e822,
        64'h11018082_610564a2,
        64'h644260e2_fc241d30,
        64'h30ef4ea5_05130000,
        64'h65174da5_85930000,
        64'h65970880_061323e6,
        64'h86930000_569702f5,
        64'h026384ae_842a4200,
        64'h07b7ec06_e426e822,
        64'h11018082_556dbfe5,
        64'h0007ac23_80824501,
        64'hcf980200_071300d7,
        64'h17634691_00d70d63,
        64'h711c46a1_59588082,
        64'h6149640a_60aaf83f,
        64'hf0ef0808_f01ff0ef,
        64'h0808e85f_f0ef0808,
        64'h85a26622_f71ff0ef,
        64'he42ee506_0808842a,
        64'he1227175_80826105,
        64'h31050513_00007517,
        64'h60e2fca7_1de3fef6,
        64'h8fa3fec6_8f230007,
        64'hc78397ae_00064603,
        64'h8bbd962e_0047d613,
        64'h07050689_0007c783,
        64'h00e107b3_45415765,
        64'h85930000_659734e6,
        64'h86930000_76974701,
        64'h3e5020ef_ec06850a,
        64'h46410505_05931101,
        64'h8082e13c_b8078793,
        64'h00000797_ed3c639c,
        64'h14078793_00007797,
        64'he93c0405_3423639c,
        64'h14878793_00007797,
        64'h80826145_69a26942,
        64'h64e27402_70a2fd24,
        64'hfde34501_97828522,
        64'h603cfc1c_078e643c,
        64'h0124f563_3f3020ef,
        64'h95224581_92011602,
        64'h0006091b_40a9863b,
        64'h449d0400_099300e7,
        64'h802397a2_f8000713,
        64'h00178513_e84af406,
        64'he44eec26_842a03f7,
        64'hf793f022_7179653c,
        64'h80826161_6ba26b42,
        64'h6ae27a02_79a27942,
        64'h74e26406_60a6b7c9,
        64'h97824401_852660bc,
        64'h01741763_99d64159,
        64'h09334a70_20ef0144,
        64'h043b8656_00848533,
        64'h85ce020a_da93020a,
        64'h1a930009_0a1b00f9,
        64'h74639381_17820007,
        64'h8a1b408b_07bb0400,
        64'h0b930400_0b13e53c,
        64'h893289ae_84aa97b2,
        64'h03f7f413_ec56f052,
        64'he486e45e_e85af44e,
        64'hf84afc26_e0a2715d,
        64'h653c8082_61056922,
        64'h64c2cd70_cd34c97c,
        64'h05052823_00c8863b,
        64'h00d306bb_00fe07bb,
        64'h010e883b_6462f3ff,
        64'h1de300e5_87bb0005,
        64'h869b0003_861b0f91,
        64'h8f5d0157_171b00b7,
        64'h579b9f3d_00774733,
        64'h9fa18f4d_fff74713,
        64'h0007081b_00b385bb,
        64'h40809fa1_8dd50115,
        64'hd59b94aa_00f5969b,
        64'h048a9db5_ffc2a403,
        64'h8db902c1_0075e5b3,
        64'hfff7c593_023fc483,
        64'h9ead00c7_03bb00c3,
        64'he633400c_9ead0166,
        64'h561b00a6_139b0082,
        64'ha5839e2d_8e3d8e59,
        64'hfff6c613_9db100f8,
        64'h073b0107_683301a8,
        64'h581b0003_a5839e2d,
        64'h0068171b_0107083b,
        64'h0042a583_9f2d942a,
        64'h040a418c_95aa058a,
        64'h93aa038a_020fc583,
        64'h9f2d022f_c403021f,
        64'hc3830002_a70300d7,
        64'h45b38f5d_fff64713,
        64'h49028293_00005297,
        64'hf45f17e3_00e407bb,
        64'h0004069b_0005861b,
        64'h02918f5d_0177171b,
        64'h0097579b_9f3d8f21,
        64'h9fa58f2d_0007081b,
        64'h00d5843b_8ec10009,
        64'h24830106_d69b9fa5,
        64'h0106941b_992a9ea1,
        64'h090a8ead_00e7c6b3,
        64'hffc3a483_9c3500c7,
        64'h05bb03c1_8e4d0156,
        64'h561b0132_c90300b6,
        64'h159b4080_9e2d9ea1,
        64'h94aa8db9_048a00f8,
        64'h073b0083_a4039e21,
        64'h01076833_01c8581b,
        64'h0048171b_0122c483,
        64'h0107083b_40809e21,
        64'h94aa048a_0043a403,
        64'h9f210112_c4839f25,
        64'h400000c5_c4b3942a,
        64'h040a00d7_c5b30003,
        64'ha7030102_c40350e3,
        64'h83930000_539782fe,
        64'h598f8f93_00005f97,
        64'hf25f1ee3_00e407bb,
        64'h0004069b_0003861b,
        64'h0005881b_8f5d0147,
        64'h171b00c7_579b9f3d,
        64'h00774733_8f6d0083,
        64'hc7339fb9_00d3843b,
        64'h8ec14098_0126d69b,
        64'h9fb900e6_941b94aa,
        64'h048affcf_a7039eb9,
        64'h0fc18ead_ffff4483,
        64'h8efd0075_c6b30f11,
        64'h9f3500c5_83bb00c3,
        64'he6334018_9eb90176,
        64'h561b0096_139b008f,
        64'ha7039e39_8e3d8e75,
        64'h00b7c633_9f3100f8,
        64'h05bb0105_e8330003,
        64'ha70301b8_581b9e39,
        64'h0058159b_0105883b,
        64'h004fa703_9db9942a,
        64'h040a4318_972a070a,
        64'h93aa038a_000f4703,
        64'h9db9002f_4403001f,
        64'h4383000f_a58300b6,
        64'hc7338df1_00d7c5b3,
        64'h67828293_00005297,
        64'h5b0f8f93_00005f97,
        64'h678f0f13_00005f17,
        64'hf45f17e3_00e387bb,
        64'h0003869b_0005881b,
        64'h0f418f5d_0167171b,
        64'h00a7579b_9f3d8f2d,
        64'h9fa10077_77338f2d,
        64'h0007061b_00d703bb,
        64'hffcfa403_9fa100d3,
        64'he6b30116_969b00f6,
        64'hd39b0076_86bb8ebd,
        64'h00cf2403_8ef900b7,
        64'hc6b300d3_83bb00c5,
        64'h873b0083_83bb8e59,
        64'h0146561b_00c6171b,
        64'h9e39008f_23838e35,
        64'h8e6d00f6_c6339f31,
        64'h00f805bb_0077073b,
        64'h0105e833_0198581b,
        64'h0078159b_0105883b,
        64'h004f2703_ff4fa383,
        64'h9db90075_85bb0fc1,
        64'h008fa403_000f2583,
        64'h000fa383_00b64733,
        64'h8dfd00c6_c5b3636f,
        64'h8f930000_5f978876,
        64'h87f2869a_86460405,
        64'h02938f2a_e44ae826,
        64'hec221101_05c52883,
        64'h05852303_05452e03,
        64'h05052e83_bf81842a,
        64'hbdd100e7_85a34721,
        64'h6786a8df_d0ef082c,
        64'h462d6506_ab7fd0ef,
        64'h45810200_06136506,
        64'hf8350005_041ba19f,
        64'he0ef1028_d3c10181,
        64'h478302f5_1b634791,
        64'hb7710005_041b8b2f,
        64'he0ef00f5_02234785,
        64'h752200f5_00235795,
        64'hb7c50785_00c68023,
        64'h96be0834_b77df0f7,
        64'h13e30e50_07930181,
        64'h470300d7_79630007,
        64'h869b0200_06134729,
        64'h93810206_1793f8f6,
        64'he9e30007_069b00d5,
        64'h80230705_95ba082c,
        64'hfe6702e3_b7ddffc8,
        64'h1be30008_05630005,
        64'hc8030585_80826125,
        64'h644660e6_85224419,
        64'hfeb045e3_4185d59b,
        64'h0185959b_a8310006,
        64'h8e1bada5_85930000,
        64'h759792c1_16c23681,
        64'h0108ec63_03085813,
        64'h1842f9f6_881b92c1,
        64'h03059693_0017061b,
        64'h0006c583_00e506b3,
        64'h432d48e5_4701fec6,
        64'h86e30006_c68396aa,
        64'h92810207_1693fff7,
        64'h871bb77d_87bab745,
        64'h2785a0e9_00e78ca3,
        64'h00078ba3_00078b23,
        64'h04600713_00e78c23,
        64'h02100713_6786bb1f,
        64'hd0ef082c_462dc7e5,
        64'h65060181_47831005,
        64'h15632501_ac3fe0ef,
        64'h10284585_e0450005,
        64'h041bbccf_e0efda02,
        64'h10284581_ebb10200,
        64'h0613eb29_00074703,
        64'h972a9301_02079713,
        64'h47810001_0c236522,
        64'he4710005_041beddf,
        64'hd0efec86_e8a21028,
        64'h002c4605_e42a711d,
        64'hb7d5842a_bf550004,
        64'h802300f5_15634791,
        64'h80826125_690664a6,
        64'h644660e6_852200a9,
        64'h2023c15f_d0ef953e,
        64'h03478793_02700793,
        64'h00e68463_00054683,
        64'h04300793_470d6562,
        64'he0150005_041be63f,
        64'hd0ef510c_65620209,
        64'h0a63fec7_83e3177d,
        64'h0007c783_97a69381,
        64'h17820007_869bfff6,
        64'h879bce89_00070023,
        64'h02000613_46ad00b4,
        64'h8713c8df_d0ef8526,
        64'h462d75c2_e93d2501,
        64'hb97fe0ef_08284585,
        64'he5592501_c9efe0ef,
        64'hd2020828_4581c4b9,
        64'he0510005_041bf95f,
        64'hd0efec86_e8a20828,
        64'h4601002c_893284ae,
        64'he42ae0ca_e4a6711d,
        64'h80826125_644660e6,
        64'h2501acef_e0ef00f5,
        64'h02234785_00e78ca3,
        64'h0087571b_00e78c23,
        64'h00445703_00e78ba3,
        64'h0087571b_00e78b23,
        64'h75220064_5703cb85,
        64'h6786eb95_0207f793,
        64'h00b7c783_451967a6,
        64'he1292501_99dfe0ef,
        64'he4be1028_083c65a2,
        64'he9292501_80afe0ef,
        64'hec861028_002c4605,
        64'h842ee42a_e8a2711d,
        64'hbfcd47a1_8082614d,
        64'h853e64ea_740a70aa,
        64'h0005079b_b48fe0ef,
        64'h6506e791_0005079b,
        64'he18fe0ef_008800f7,
        64'h022306d7_07a34785,
        64'h06f704a3_0086d69b,
        64'h0106d69b_0087d79b,
        64'h0107d79b_0107979b,
        64'h06f70423_0107d79b,
        64'h06f70723_0107969b,
        64'h57d602f6_9c630557,
        64'h468302e0_07936706,
        64'hefa90005_079bfbbf,
        64'hd0ef8522_c1bd4789,
        64'h0005059b_ca4fe0ef,
        64'h85220005_059bf25f,
        64'hd0ef85a6_00044503,
        64'h06f70763_57d64736,
        64'hcbb58bc1_00b4c783,
        64'h00f40223_478500f4,
        64'h85a30207_e7936406,
        64'h02814783_df7fd0ef,
        64'h00d48513_02a10593,
        64'h464d648a_ebdd0005,
        64'h079bdcbf_e0ef10a8,
        64'h0ce79263_4711cbf1,
        64'h0005079b_a9dfe0ef,
        64'h10a86582_0c054c63,
        64'h47adefdf_d0ef850a,
        64'he33fd0ef_10a8008c,
        64'h02800613_e3ffd0ef,
        64'h102805ad_46550e05,
        64'h8d634791_65e61007,
        64'h11630207_77134799,
        64'h00b7c703_77861007,
        64'h99630005_079bae7f,
        64'he0eff0be_083cf4be,
        64'h008865a2_67861207,
        64'h95630005_079b95cf,
        64'he0efed26_f122f506,
        64'h0088002c_4605e02e,
        64'he42a7171_80826165,
        64'h64e67406_70a62501,
        64'hc94fe0ef_00f50223,
        64'h47850087_05a38c3d,
        64'h02747413_8c658cbd,
        64'h752200b7_4783c30d,
        64'h6706e39d_0207f793,
        64'h00b7c783_451967a6,
        64'he9152501_b55fe0ef,
        64'he4be1028_083c65a2,
        64'he1312501_9c2fe0ef,
        64'hf4861028_4605002c,
        64'h843284ae_e42aeca6,
        64'hf0a27159_b7c54421,
        64'h8082614d_6d466ce6,
        64'h7c067ba6_7b467ae6,
        64'h6a0a69aa_694a64ea,
        64'h740a70aa_8522f2bf,
        64'he0ef85a6_7522441d,
        64'hb7498c6a_0ffbfb93,
        64'hf53fd0ef_3bfd855a,
        64'h45812000_0613ec09,
        64'h0005041b_8d4fe0ef,
        64'h01950223_03852823,
        64'h001c0d1b_7522a82d,
        64'h0005041b_d50fe0ef,
        64'h00f50223_47850127,
        64'h8aa30157_8a230137,
        64'h8da30147_8d2300e7,
        64'h8ca30007_8ba30007,
        64'h8b230460_071300e7,
        64'h8c230210_071300e7,
        64'h85a37522_47416786,
        64'he8350005_041bf5ff,
        64'he0ef1028_040b9963,
        64'h4c850027_4b8306f4,
        64'h04a306d4_07a30087,
        64'hd79b0086_d69b0107,
        64'hd79b0106_d69b0107,
        64'h979b06f4_04230107,
        64'hd79b0107_969b06f4,
        64'h07234781_00f69363,
        64'h571400d6_166357d2,
        64'h00074603_468d0574,
        64'h0aa37722_ff7fd0ef,
        64'h05440513_85da0524,
        64'h04a30554_04230534,
        64'h07a30544_07230404,
        64'h05a30404_05230374,
        64'h0a230200_061304f4,
        64'h06a30089_591b0089,
        64'hd99b0460_07930ff4,
        64'hfa1304f4_062302e0,
        64'h0b930109_591b0210,
        64'h07930109_d99b02f4,
        64'h0fa30109_191b0104,
        64'h999b0ff9_7a9347c1,
        64'h87afe0ef_855a0200,
        64'h0593462d_886fe0ef,
        64'h855a0005_0c1b4581,
        64'h20000613_03440b13,
        64'hf60fe0ef_85220104,
        64'hd91b85a6_74221604,
        64'h12630005_041ba8cf,
        64'he0ef16f4_88634405,
        64'h57fd16f4_8c634409,
        64'h75224785_18048063,
        64'h0005049b_b33fe0ef,
        64'h45817522_18079d63,
        64'h0207f793_00b7c783,
        64'h441967a6_1af41563,
        64'h47911c04_07630005,
        64'h041bd53f_e0efe4be,
        64'h1028083c_65a21c04,
        64'h12630005_041bbc4f,
        64'he0efe8ea_ece6f0e2,
        64'hf4def8da_fcd6e152,
        64'he54ee94a_ed26f506,
        64'hf1221028_002c4605,
        64'he42a7171_b7edf551,
        64'h250191ef_f0ef85a2,
        64'h7502bf61_2501f12f,
        64'he0ef7502_e411f155,
        64'h25019e3f_e0ef1008,
        64'hfaf518e3_4791d94d,
        64'h2501838f_f0ef00a8,
        64'h4581f161_2501941f,
        64'he0efcaa2_00a84589,
        64'h952fe0ef_00a8100c,
        64'h02800613_fc878de3,
        64'h01492783_c89d88c1,
        64'hcc0d0005_041baccf,
        64'he0ef0009_45037902,
        64'h80826149_794674e6,
        64'h640a60aa_451dcb81,
        64'h0014f793_00b5c483,
        64'hc59975e2_eb890207,
        64'hf79300b7_c7834519,
        64'h6786e105_2501e27f,
        64'he0efe0be_1008081c,
        64'h65a2e905_2501c94f,
        64'he0eff8ca_fca6e122,
        64'he5061008_002c4605,
        64'he42a7175_b7b100f4,
        64'h0523fbf7_f79300a4,
        64'h4783f55d_250171e0,
        64'h40ef0304_05930017,
        64'hc5034685_4c50601c,
        64'hdba50407_f79300a4,
        64'h4783fcf9_6ae34d1c,
        64'h6008fcf9_00e34509,
        64'h4785b769_449db7e1,
        64'h2501a1ef_f0ef85ca,
        64'h6008f979_2501b25f,
        64'he0ef167d_10000637,
        64'h4c0cb7dd_450502f9,
        64'h146357fd_0005091b,
        64'h941fe0ef_4c0cbf7d,
        64'h84aa00a4_05a3c539,
        64'h00042a23_2501a5af,
        64'hf0ef484c_ef016008,
        64'h00f40523_c8180207,
        64'he793fed7_72e34814,
        64'h4458cf39_0027f713,
        64'h00a44783_80826105,
        64'h64a26902_85266442,
        64'h60e20007_849bcb91,
        64'h00b44783_e4910005,
        64'h049bbb8f_e0ef842a,
        64'he04aec06_e426e822,
        64'h1101bfad_8a2abfbd,
        64'h4a09b749_4a05b7c5,
        64'h39f10911_2485e111,
        64'h65820155_75332501,
        64'haa2fe0ef_e02e854a,
        64'hb745fc0c_94e33cfd,
        64'h39f90909_2485e391,
        64'h8fd90087_979b0009,
        64'h47030019_4783038b,
        64'h91632000_09930344,
        64'h091385ce_e9212501,
        64'hd04fe0ef_0015899b,
        64'h85220009_9e631afd,
        64'h4c094481_49814901,
        64'h10000ab7_504cb74d,
        64'h009b2023_00f402a3,
        64'h0017e793_c8040054,
        64'h4783fef9_63e32905,
        64'h4c1c2485_e1110955,
        64'h08630935_08632501,
        64'ha49fe0ef_852285ca,
        64'h4a8559fd_44814909,
        64'h02fb9f63_47850004,
        64'h4b838082_61656ce2,
        64'h7c027ba2_7b427ae2,
        64'h6a0669a6_694664e6,
        64'h85527406_70a600fb,
        64'h202302f7_6263ffec,
        64'h871b481c_01842c83,
        64'h6000000a_1c630005,
        64'h0a1be70f_e0efec66,
        64'hf062f45e_fc56e4ce,
        64'he8caeca6_f486e0d2,
        64'h8522002c_46018b2e,
        64'he42af85a_8432f0a2,
        64'h7159bfcd_44198082,
        64'h616564e6_740670a6,
        64'h8522c00f_e0ef1028,
        64'h85a6c489_cf816786,
        64'he8010005_041b85ef,
        64'hf0efe4be_1028083c,
        64'h65a2e00d_0005041b,
        64'hecefe0ef_f486f0a2,
        64'h1028002c_460184ae,
        64'he42aeca6_7159bf65,
        64'h84aad16d_bf7d0004,
        64'h2a2300f5_16634791,
        64'h2501f77f_e0ef8522,
        64'h4581c58f_e0ef8522,
        64'h85ca0004_2a2302f5,
        64'h13634791_2501b34f,
        64'hf0ef8522_45810224,
        64'h30238082_614564e2,
        64'h69428526_740270a2,
        64'h0005049b_c4ffe0ef,
        64'h85224581_00091f63,
        64'he8890005_049bd8cf,
        64'he0ef892e_842af406,
        64'he84aec26_f0227179,
        64'h80820141_640260a2,
        64'h00043023_e1192501,
        64'hdaefe0ef_842ae406,
        64'he0221141_b7c1fcf5,
        64'h01e34791_bfdd4525,
        64'h80826121_744270e2,
        64'hf971fcf5_0be34791,
        64'h2501cadf_e0ef00f4,
        64'h14230067_d7838522,
        64'h458167e2_c448e24f,
        64'he0ef0007_c50367e2,
        64'ha02d0004_30234515,
        64'he7898bc1_00b5c783,
        64'hcd996c0c_e5292501,
        64'h968ff0ef_f01c101c,
        64'he01c8522_65a267e2,
        64'he1152501_fdafe0ef,
        64'h0828002c_4601842a,
        64'hc52de42e_f822fc06,
        64'h7139b7bd_c45c0137,
        64'h87bb4134_84bbcc0c,
        64'h445cfaf5_fae34f9c,
        64'h601cfaba_fee3fd45,
        64'h88e30005_059bc3ff,
        64'he0efbf69_84cee599,
        64'h0005059b_fcbfe0ef,
        64'hcb818b89_600800a4,
        64'h4783b765_cc0cc84c,
        64'hb5ed4905_00f405a3,
        64'h478500f5_976357fd,
        64'hbded4909_00f405a3,
        64'h478900f5_97634785,
        64'h0005059b_802ff0ef,
        64'he595484c_bfb19ca9,
        64'h0094d49b_cd112501,
        64'hc79fe0ef_6008d7b5,
        64'h1ff4f793_c45c9fa5,
        64'h445c0499_ea634a85,
        64'h5a7dd1c1_9c9dc45c,
        64'h27814c0c_8ff94130,
        64'h07bb02c6_ed630337,
        64'h563b0336_d6bbfff4,
        64'h869b377d_c7290097,
        64'h999b0025_47836008,
        64'hbf59cc44_ed352501,
        64'h2ef040ef_85ce0017,
        64'hc5038626_4685601c,
        64'h00f40523_fbf7f793,
        64'h00a44783_ed512501,
        64'h341040ef_0017c503,
        64'h85ce4685_601cc385,
        64'h0407f793_03040993,
        64'h00a44783_fc960ee3,
        64'h4c50d3e5_1ff7f793,
        64'h445c4481_bf7d00f4,
        64'h05230207_e79300a4,
        64'h4783c81c_fcf778e3,
        64'h4818445c_e4bd0004,
        64'h26234458_84bae391,
        64'h8b8900a4_47830097,
        64'h77634818_80826121,
        64'h6aa26a42_69e27902,
        64'h74a2854a_744270e2,
        64'h0007891b_cf8900b4,
        64'h47830009_17630005,
        64'h091bfa8f_e0ef84ae,
        64'h842ae456_e852ec4e,
        64'hfc06f04a_f426f822,
        64'h7139b721_fe9465e3,
        64'hfee78fa3_24050785,
        64'h00074703_97369281,
        64'h02041693_67220789,
        64'hbdf54545_b7e900e6,
        64'h0023fc97_4703972a,
        64'h10889301_17020007,
        64'h059bfff5_871bb7e1,
        64'h2785bf19_9c3d0126,
        64'h0023fff7_c793e989,
        64'h963a9301_02069713,
        64'h662236fd_86a285be,
        64'h04e46063_0037871b,
        64'he705fc97_47039736,
        64'h10949301_02079713,
        64'h4781f48f_e0ef1828,
        64'h100cb761_4509f6e5,
        64'h12e367a2_4711dd61,
        64'h2501a86f_f0ef1828,
        64'h45810135_0e632501,
        64'h897fe0ef_0007c503,
        64'h65c677e2_e1052501,
        64'he46ff0ef_18284581,
        64'hf9512501_f4ffe0ef,
        64'h18284581_c2aa8bdf,
        64'he0ef0007_c50365c6,
        64'h77e2f55d_2501e6cf,
        64'hf0ef1828_4581fd4d,
        64'h2501f75f_e0ef1828,
        64'h45858082_614979a6,
        64'h794674e6_640a60aa,
        64'h00078023_078d00e7,
        64'h812302f0_07130e94,
        64'h156300e7_80a303a0,
        64'h071300e7_80230307,
        64'h071b5227_47030000,
        64'h8717e505_67a24501,
        64'h04099163_4996c2be,
        64'h4bdc02f0_09138426,
        64'h77e2ecbe_081ce521,
        64'h2501ab9f_e0ef1828,
        64'h002c4601_84ae0005,
        64'h0023f4ce_f8cae122,
        64'he506e42a_fca67175,
        64'hbfd94415_fcf41ee3,
        64'h4791b7c5_c8c8965f,
        64'he0ef0004_c50374a2,
        64'hcb998bc1_00b5c783,
        64'h80826165_64e67406,
        64'h70a68522_cbd85752,
        64'h77a2e991_6586e41d,
        64'h0005041b_cb4ff0ef,
        64'he4be1028_083c65a2,
        64'hec190005_041bb25f,
        64'he0efeca6_f486f0a2,
        64'h1028002c_4601e42a,
        64'h7159bfe5_452d8082,
        64'h610560e2_45015ca7,
        64'h8b230000_87970005,
        64'h4a63945f_e0efec06,
        64'h0028e42a_11018082,
        64'h01416402_60a20004,
        64'h3023e119_25019b5f,
        64'he0ef8522_e9012501,
        64'hf01ff0ef_842ae406,
        64'he0221141_80820141,
        64'h640260a2_4505ea3f,
        64'he06f0141_60a26402,
        64'h00f50223_478500f4,
        64'h0523fdf7_f7936008,
        64'h00a44783_000789a3,
        64'h00078923_00e78ca3,
        64'h00d78da3_04600713,
        64'h0086d69b_00e78c23,
        64'h02100713_0106d69b,
        64'h00e78aa3_0087571b,
        64'h0107571b_0107171b,
        64'h00e78a23_0107571b,
        64'h0107169b_00e78d23,
        64'h00078ba3_00078b23,
        64'h485800e7_8fa300d7,
        64'h8f230187_571b0107,
        64'h569b00d7_8ea300e7,
        64'h8e230086_d69b0106,
        64'hd69b0107_169b4818,
        64'h00e785a3_02076713,
        64'h00b7c703_741ce155,
        64'h2501b5ff_e0ef6008,
        64'h500c00f4_0523fbf7,
        64'hf79300a4_4783ed4d,
        64'h25016ab0_40ef0304,
        64'h05930017_c5034685,
        64'h4c50601c_c3950407,
        64'hf793cf61_0207f713,
        64'h00a44783_e16d2501,
        64'hab7fe0ef_842ae406,
        64'he0221141_bd15499d,
        64'hb5f1c81c_bf4100f4,
        64'h05230407_e79300a4,
        64'h47839b5f_e0ef9522,
        64'h85d28626_03050513,
        64'h0007049b_01277463,
        64'h40ab873b_1ff57513,
        64'h0009049b_444801b4,
        64'h2e23fd01_25016ed0,
        64'h40ef85da_46850017,
        64'hc50300d7_7a634458,
        64'h481400c7_0e634c58,
        64'hbdc900fa_a0239fa5,
        64'h000aa783_c45c9fa5,
        64'h4099093b_445c9a3e,
        64'h93810204_97930094,
        64'h949b00f4_0523fbf7,
        64'hf79300a4_4783a29f,
        64'he0ef855a_95d22000,
        64'h06139181_15820097,
        64'h959b0297_f26341b5,
        64'h87bb4c4c_f1492501,
        64'h789040ef_85d286a6,
        64'h0017c503_41a684bb,
        64'h00e6f463_0104873b,
        64'h0099549b_0027c683,
        64'h072c7a63_67a28db2,
        64'h00a8063b_000d081b,
        64'hd1592501_964ff0ef,
        64'he43e853e_4c0c601c,
        64'h00f40523_fbf7f793,
        64'h00a44783_f9692501,
        64'h7d9040ef_85da0017,
        64'hc5034685_4c50601c,
        64'hc38d0407_f79300a4,
        64'h4783c85c_e311cc1c,
        64'h4858bf89_498500f4,
        64'h05a34785_01979763,
        64'hb78500f4_05230207,
        64'he79300a4_478312f7,
        64'h6b634818_445cf3fd,
        64'h0005079b_d6aff0ef,
        64'h4c0cb749_498900f4,
        64'h05a34789_02e79863,
        64'h4705cb91_4581485c,
        64'hef01040d_1a630ffd,
        64'h7d1301a7_fd3337fd,
        64'h00254783_00975d1b,
        64'h60081407_94631ff7,
        64'h77930409_04634458,
        64'h5cfd0304_0b131ff0,
        64'h0c132000_0b9304f7,
        64'h6e630127_873b445c,
        64'h1a078263_8b8900a4,
        64'h47838082_61096de2,
        64'h7d027ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_854e7446,
        64'h70e60007_899bc39d,
        64'h00b44783_00099763,
        64'h0005099b_ca3fe0ef,
        64'h8ab68932_8a2e842a,
        64'h0006a023_ec6ef06a,
        64'hf466f862_fc5ee0da,
        64'hf4a6fc86_e4d6e8d2,
        64'heccef0ca_f8a27119,
        64'hb585499d_bf9dbb1f,
        64'he0ef8552_95a28626,
        64'h03058593_0007049b,
        64'h01277463_40bb873b,
        64'h1ff5f593_0009049b,
        64'h444c01b4_2e23f10d,
        64'h25010e80_50ef85da,
        64'h0017c503_86424685,
        64'h601c00f4_0523fbf7,
        64'hf7936822_00a44783,
        64'hf1312501_13c050ef,
        64'he44285da_46850017,
        64'hc503c30d_04077713,
        64'h00a44703_05060163,
        64'h4c50bf39_00faa023,
        64'h9fa5000a_a783c45c,
        64'h9fa54099_093b445c,
        64'h9a3e9381_02049793,
        64'h0094949b_c3ffe0ef,
        64'h955285da_20000613,
        64'h91011502_0097951b,
        64'h0097fc63_41b507bb,
        64'h4c48c385_0407f793,
        64'h00a44783_f9452501,
        64'h176050ef_85d28642,
        64'h86a60017_c50341a6,
        64'h84bb00e6_f46300c4,
        64'h873b0099_549b0027,
        64'hc683072c_7a6367a2,
        64'h8dc200a6_083b000d,
        64'h061bd579_2501b86f,
        64'hf0efe43e_853e4c0c,
        64'h601ccc08_b7954985,
        64'h00f405a3_47850195,
        64'h1763b7e5_2501bc6f,
        64'hf0ef4c0c_bfb54989,
        64'h00f405a3_478900a7,
        64'hec634785_4848eb11,
        64'h020d1963_0ffd7d13,
        64'h01a7fd33_37fd0025,
        64'h47830097_5d1b6008,
        64'h12079163_1ff77793,
        64'h4458fa09_0ae35cfd,
        64'h03040b13_1ff00c13,
        64'h20000b93_0006091b,
        64'h00f67463_893e40f9,
        64'h07bb445c_01042903,
        64'h16078c63_8b8500a4,
        64'h47838082_61096de2,
        64'h7d027ca2_7c427be2,
        64'h6b066aa6_6a4669e6,
        64'h790674a6_854e7446,
        64'h70e60007_899bc39d,
        64'h662200b4_47830009,
        64'h98630005_099be85f,
        64'he0ef8ab6_e4328a2e,
        64'h842a0006_a023ec6e,
        64'hf06af466_f862fc5e,
        64'he0daf0ca_f4a6fc86,
        64'he4d6e8d2_eccef8a2,
        64'h7119bdd1_4525bf51,
        64'hec079ee3_451d8b85,
        64'hfa0900e3_00297913,
        64'hee0716e3_0107f713,
        64'h451100b4_4783ee05,
        64'h1de3bdf5_450100f4,
        64'h94230124_b0230004,
        64'hae230004_a623c888,
        64'h00695783_daffe0ef,
        64'h01c40513_c8c8f35f,
        64'he0ef0009_45030004,
        64'h85a3d09c_01348523,
        64'hf4800309_278385a2,
        64'h79220209_e993c399,
        64'h0089f793_f1392501,
        64'h80cff0ef_01252623,
        64'h85d6397d_7522fd21,
        64'h2501e1ff_f0ef030a,
        64'h2a838552_85ca0209,
        64'h036300fa_02230005,
        64'h091b0004_0aa30004,
        64'h0a230004_0da30004,
        64'h0d234785_f9bfe0ef,
        64'h85a2000a_45030004,
        64'h0fa30004_0f230004,
        64'h0ea30004_0e230004,
        64'h05a300e4_0c230004,
        64'h0ba30004_0b2300e4,
        64'h08230004_07a30004,
        64'h072300f4_0ca300f4,
        64'h08a30210_07130460,
        64'h07937a22_0089e993,
        64'h6406a021_08090a63,
        64'h00897913_fff94521,
        64'h00497793_f3fd8bc5,
        64'h451d00b4_47838082,
        64'h61496ae6_7a0679a6,
        64'h794674e6_640a60aa,
        64'hc9052501_e7dff0ef,
        64'h102800f5_17634791,
        64'hc1151007_8e6301f9,
        64'h799301c9_77934519,
        64'he011e119_64062501,
        64'hb61ff0ef_e4be1028,
        64'h083c65a2_e91d2501,
        64'h9ceff0ef_1028002c,
        64'h8a7984aa_89320005,
        64'h30231605_0c63e42e,
        64'hecd6f0d2_f4cef8ca,
        64'hfca6e122_e5067175,
        64'hbfe5452d_80826121,
        64'h70e22501_a02ff0ef,
        64'h0828080c_460100f6,
        64'h18634785_cb114501,
        64'he39897aa_00070023,
        64'hc3196762_00070023,
        64'hc3196622_631800a7,
        64'h8733050e_cb478793,
        64'h00009797_04054263,
        64'h832ff0ef_f42ee432,
        64'he82efc06_1028ec2a,
        64'h71398082_4509bf4d,
        64'h4505bf5d_4509bf65,
        64'hfaf4e7e3_0004891b,
        64'h4c1c00f4_02a30017,
        64'he7930054_4783c81c,
        64'h27850137_8a63481c,
        64'hfd712501_8abff0ef,
        64'h852285ca_46010334,
        64'h8c630344_8c638082,
        64'h61456a02_69a26942,
        64'h64e27402_70a24501,
        64'he8910005_049bed6f,
        64'hf0ef8522_85ca59fd,
        64'h4a0506f5_f063892e,
        64'h842ae052_e44eec26,
        64'hf406e84a_f0227179,
        64'h4d1c08b7_f0634785,
        64'h80826105_64a28526,
        64'h644260e2_00e78223,
        64'h4705601c_80eff0ef,
        64'h462d6c08_700c838f,
        64'hf0ef4581_02000613,
        64'h6c08e085_0005049b,
        64'ha34ff0ef_6008484c,
        64'he49d0005_049bfa9f,
        64'hf0ef842a_ec06e426,
        64'he8221101_80826105,
        64'h64a26442_60e2451d,
        64'h00f51363_4791dd79,
        64'h2501bb7f_f0ef8522,
        64'h4585cb99_00978d63,
        64'h0007c783_6c1ced09,
        64'h2501a7ef_f0ef6008,
        64'h484c0e50_0493e50d,
        64'h250187df_f0ef842a,
        64'he426ec06_e8224581,
        64'h1101bfe5_4511b7cd,
        64'h00042a23_d9452501,
        64'hbfdff0ef_85224581,
        64'h80826145_69a26942,
        64'h64e27402_70a24501,
        64'h00979a63_0017b793,
        64'h17e18bfd_03378063,
        64'h03270263_03f7f793,
        64'h00b7c783_c3210007,
        64'hc7036c1c_e1292501,
        64'haecff0ef_6008a0b1,
        64'hc90de199_484c49bd,
        64'h0e500913_451184ae,
        64'hf406842a_e44ee84a,
        64'hec26f022_7179bdc1,
        64'h0ff77713_0017e793,
        64'h3701eca8_efe30ff5,
        64'h7513f9f7_051beea8,
        64'hf3e30ff5_7513fbf7,
        64'h051bb575_4519ef07,
        64'h19e30008_06630005,
        64'h48030c25_05130000,
        64'h85170005_4c634185,
        64'h551b0187_151b02b6,
        64'hf263fd37_0ae3f357,
        64'h09e3f347_0be3f2e3,
        64'h7de30007_47039722,
        64'h93011702_0017061b,
        64'h873245ad_46a10ff7,
        64'hf7930027_979b0565,
        64'h9a63b5a1_c4c8ae4f,
        64'hf0ef0007_c503609c,
        64'hdbe58bc1_00b5c783,
        64'h6c8cfbe5_8b91b705,
        64'h4515f315_bfd94511,
        64'hb72d4501_e6070ae3,
        64'h0004bc23_0004a623,
        64'hcb990207_f7930047,
        64'hf713f4e5_13e34711,
        64'hc51500b7_c783709c,
        64'hf1279de3_b7c50106,
        64'h6613fed7_14e34685,
        64'h0037f713_bded00c9,
        64'h05a30086_661300e7,
        64'h94634711_8bb10ff7,
        64'hf7930027_979b0165,
        64'h9f6300e9_00234715,
        64'h00e69563_0e500713,
        64'h00094683_c6e54601,
        64'h00e57363_46119432,
        64'h02000513_92011602,
        64'ha8652685_00e50023,
        64'h954a9101_02069513,
        64'h0027e793_a2110505,
        64'ha8c948e5_02000313,
        64'h478145a1_47014681,
        64'hb78d0240_0793943a,
        64'h12f6e763_02000693,
        64'hf75787e3_b7b54709,
        64'hb73d0405_80826121,
        64'h6b026aa2_6a4269e2,
        64'h790274a2_744270e2,
        64'h0004bc23_2501a81f,
        64'hf0ef8526_4581bf35,
        64'hc55c4bdc_611ca0e1,
        64'hdd5d2501_df9ff0ef,
        64'h85264581_0cd60a63,
        64'hfff64603_0006c683,
        64'h00f58633_078500f7,
        64'h06b3708c_ef898ba1,
        64'h00b74783_12078063,
        64'h00074783_6c981005,
        64'h11632501_ce0ff0ef,
        64'h608848cc_492d1005,
        64'h19632501_adfff0ef,
        64'h85264581_00f905a3,
        64'h02000793_943a0947,
        64'h9b63470d_1d378963,
        64'h00244783_00f900a3,
        64'h02e00793_0b379463,
        64'h00144783_01390023,
        64'h0d379663_00044783,
        64'hb42ff0ef_854a0200,
        64'h0593462d_0204b903,
        64'h0d578463_0d478663,
        64'h00044783_4b2102e0,
        64'h099305c0_0a9302f0,
        64'h0a130ce7_f06347fd,
        64'h00044703_0004a623,
        64'h04050ce7_946305c0,
        64'h071300e7_8663842e,
        64'h84aa02f0_07130005,
        64'hc783e05a_e456e852,
        64'hec4ef04a_fc06f426,
        64'hf8227139_b7e9db1c,
        64'h27855b1c_2a856018,
        64'hf1412501_d24ff0ef,
        64'h01450223_b7b9c848,
        64'ha89ff0ef_85a6c804,
        64'h6008d91c_415787bb,
        64'h591c00fa_ed630025,
        64'h47836008_4a0502aa,
        64'h2823aabf_f0ef8552,
        64'h85a60004_3a03bf0f,
        64'hf0ef0345_05134581,
        64'h20000613_6008f579,
        64'h2501de0f_f0ef6008,
        64'hfcf48de3_57fdfcf4,
        64'h8be34785_d4bd451d,
        64'h0005049b_e83ff0ef,
        64'h480cf60a_0ee306f4,
        64'he0634d1c_6008b761,
        64'h450500f4_946357fd,
        64'hbf494509_0097e463,
        64'h47850005_049bb2ff,
        64'hf0effc0a_9fe30157,
        64'hfab337fd_00495a9b,
        64'h00254783_bf5d4501,
        64'hec1c97ce_03478793,
        64'h01241523_0996601c,
        64'hfcf775e3_0009071b,
        64'h00855783_e18dc85c,
        64'h61082785_480c0009,
        64'h9d63842a_8a2e00f9,
        64'h7993d7ed_495c8082,
        64'h61216aa2_6a4269e2,
        64'h790274a2_744270e2,
        64'h4511eb99_93c1e456,
        64'he852ec4e_f4260309,
        64'h17932905_f822fc06,
        64'h00a55903_f04a7139,
        64'hb795547d_f6f514e3,
        64'h4785dd61_2501dbdf,
        64'hf0ef8526_85ce8622,
        64'hbfb500f4_82a30017,
        64'he7930054_c783c89c,
        64'h37fdf8e7_88e3577d,
        64'hc4c0489c_02099063,
        64'he9052501_debff0ef,
        64'h852685a2_167d1000,
        64'h0637b7cd_fd241de3,
        64'hfb450ae3_05550a63,
        64'hc9012501_c0dff0ef,
        64'h852685a2_4409b7e9,
        64'h4401012a_646300f4,
        64'h67632405_4c9c5afd,
        64'h4a05844a_fef461e3,
        64'h894e4c9c_08f40263,
        64'h57fd8082_61216aa2,
        64'h6a4269e2_790274a2,
        64'h744270e2_85224405,
        64'h0087ed63_47850005,
        64'h041bc5bf_f0efa815,
        64'h490502f9_6d634d1c,
        64'h00090563_00c52903,
        64'he99189ae_84aae456,
        64'he852f04a_f822fc06,
        64'hec4ef426_7139bf79,
        64'h012a81a3_00fa8123,
        64'h0189591b_0109579b,
        64'h00fa80a3_0087d79b,
        64'h03240a23_0107d79b,
        64'h94260109_179b2901,
        64'h01256933_8d71f000,
        64'h06372501_d96ff0ef,
        64'h85569aa6_03440a93,
        64'h1fc47413_0024141b,
        64'hf80a16e3_00050a1b,
        64'hfdcff0ef_9dbd0075,
        64'hd59b515c_bf790134,
        64'h82230324_0aa30089,
        64'h591b0109_591b0109,
        64'h191b0324_0a239426,
        64'h1fe47413_0014141b,
        64'hfc0a12e3_00050a1b,
        64'h815ff0ef_9dbd0085,
        64'hd59b515c_b7e90127,
        64'he9339bc1_00f97913,
        64'h0089591b_0347c783,
        64'h015487b3_80826121,
        64'h6aa26a42_69e27902,
        64'h74a28552_744270e2,
        64'h00f48223_4785032a,
        64'h8a239aa6_0ff97913,
        64'h0049591b_c40d1ffa,
        64'hfa93000a_1f630005,
        64'h0a1b86ff_f0ef9dbd,
        64'h8526009a_d59b50dc,
        64'h00f48223_478502f9,
        64'h8a2399a6_0ff7f793,
        64'h8fd98ff5_0049179b,
        64'h00f7f713_16c16685,
        64'h0347c783_013487b3,
        64'hcc191ff9_f9930ff9,
        64'h77930019_8a9b8805,
        64'h060a1663_00050a1b,
        64'h8bdff0ef_9dbd0099,
        64'hd59b00b9_89bb515c,
        64'h0015d99b_09379463,
        64'h0ee78863_470d0ae7,
        64'h8f63842e_89324709,
        64'h00054783_0af5f063,
        64'h4a0984aa_4d1c0ab9,
        64'hf5634a09_4985e456,
        64'hf04af426_f822fc06,
        64'he852ec4e_71398082,
        64'h610564a2_85266442,
        64'h60e200e7_82234705,
        64'h601c00e7_80235715,
        64'h6c1cf3cf_f0ef4581,
        64'h02000613_6c08ec99,
        64'h0005049b_939ff0ef,
        64'h6008484c_e4950005,
        64'h049bf35f_f0ef842a,
        64'hec06e426_e8221101,
        64'h00a55583_b7954505,
        64'hbfc14134_043bf6f4,
        64'hf7e34f9c_00093783,
        64'hf69afce3_01448c63,
        64'h0005049b_e75ff0ef,
        64'hbf7d2501_e5dff0ef,
        64'h01347663_85a60009,
        64'h35030992_4a855a7d,
        64'h0027c983_84bab75d,
        64'h45010089_3c23943e,
        64'h03478793_0416883d,
        64'h00093783_00f92a23,
        64'h9fa90044_579bd171,
        64'h00992823_5788fce4,
        64'h77e30087_d703eb0d,
        64'h579800e6_9463470d,
        64'h0007c683_e0a9842e,
        64'hfee4f4e3_4f98611c,
        64'h80826121_6aa26a42,
        64'h69e27902_74a27442,
        64'h70e24509_00f49c63,
        64'h892a4785_00b51523,
        64'he456e852_ec4ef822,
        64'hfc06f04a_4544f426,
        64'h71398082_853e4785,
        64'hbfb90245_57931512,
        64'hffaff0ef_954a0345,
        64'h05131fc5_75130024,
        64'h151bf93d_2501a3bf,
        64'hf0ef9dbd_0075d59b,
        64'h515cb761_8fc90087,
        64'h979b0349_45030359,
        64'h47839922_1fe47413,
        64'h0014141b_f1452501,
        64'ha65ff0ef_9dbd0085,
        64'hd59b515c_bf4d93d1,
        64'h17d2bf65_8391c019,
        64'h8fc50087_979b8805,
        64'h03494783_994e1ff9,
        64'hf993f579_2501a93f,
        64'hf0ef0344_c483854a,
        64'h9dbd94ca_1ff4f493,
        64'h0099d59b_0014899b,
        64'h02492783_80826145,
        64'h853e69a2_694264e2,
        64'h740270a2_57fdc911,
        64'h2501ac7f_f0ef9dbd,
        64'h0094d59b_9cad515c,
        64'h0015d49b_00f71e63,
        64'h08d70d63_468d06d7,
        64'h0b63842e_46890005,
        64'h470302e5_f963892a,
        64'he44eec26_f022f406,
        64'he84a7179_4d180eb7,
        64'hf5634785_80824501,
        64'h80829d3d_02b787bb,
        64'h55480025_478300e7,
        64'hf9633779_85beffe5,
        64'h879b4d18_80826105,
        64'h64a26442_60e200a0,
        64'h35332501_671050ef,
        64'h45814601_00144503,
        64'h000402a3_67d050ef,
        64'h85a64685_d81022f4,
        64'h01a322e4_012320d4,
        64'h0ca320d4_0c230187,
        64'hd79b0107_d71b2605,
        64'h22e400a3_22f40023,
        64'h07200693_00144503,
        64'h0087571b_0107571b,
        64'h0107971b_501020e4,
        64'h0f23445c_20f40fa3,
        64'h0187d79b_0107d71b,
        64'h20e40ea3_20f40e23,
        64'h0087571b_0107571b,
        64'h0107971b_20e40d23,
        64'h02e40ba3_04100713,
        64'h481c20f4_0da302f4,
        64'h0b230610_079302f4,
        64'h0aa302f4_0a230520,
        64'h079322f4_09a3faa0,
        64'h079322f4_09230550,
        64'h07939fdf_f0ef8526,
        64'h45812000_06130344,
        64'h04930af7_1b634785,
        64'h00544703_0cf71063,
        64'h478d0004_4703ed69,
        64'h2501c01f_f0ef842a,
        64'he426ec06_e8221101,
        64'hbdcd9cbd_0017d79b,
        64'h88850297_87bb478d,
        64'hb7090014_949b00f9,
        64'h15634789_d41c9fb5,
        64'he00a84e3_b545a19f,
        64'hf0ef0544_0513b5b1,
        64'h0005099b_a27ff0ef,
        64'h05840513_b3514781,
        64'h00042a23_01240023,
        64'h00f41323_7cf71723,
        64'h00009717_93c117c2,
        64'h27857dc7_d7830000,
        64'h9797c448_a57ff0ef,
        64'h22040513_c808a61f,
        64'hf0ef21c4_051300f5,
        64'h1c632727_87932501,
        64'h614177b7_a77ff0ef,
        64'h21840513_02f51763,
        64'h25278793_25014161,
        64'h57b7a8df_f0ef0344,
        64'h051304e7_9263a557,
        64'h07134107_d79b776d,
        64'h0107979b_8fd90087,
        64'h979b0004_02a32324,
        64'h47032334_4783e13d,
        64'h2501ce7f_f0ef8522,
        64'h001a059b_06e79b63,
        64'h47054107_d79b0107,
        64'h979b8fd9_0087979b,
        64'h06444703_06544783,
        64'h08f91963_478d00f4,
        64'h02a3f800_0793c45c,
        64'hc81c57fd_ee99e6e3,
        64'h0094d49b_1ff4849b,
        64'h0024949b_d408b09f,
        64'hf0ef0604_0513f00a,
        64'h93e310e9_1163470d,
        64'hd05c0344_2023cc04,
        64'hd4580147_87bb2489,
        64'h0147073b_090900b9,
        64'h39331955_694100b6,
        64'h77634905_16556605,
        64'hf3266ce3_84ae0326,
        64'h55bb40c5_063bf4c5,
        64'h63e38732_00d7063b,
        64'h9f3d004a_d71b2781,
        64'h033486bb_dfa98fd9,
        64'h0087979b_25010424,
        64'h47030434_47831405,
        64'h0e638d5d_0085151b,
        64'h04744783_04844503,
        64'hffbd00fa_f7930154,
        64'h142300fa_eab3008a,
        64'h9a9b0454_47830464,
        64'h4a83ffc1_00f977b3,
        64'hfff9079b_2901fa09,
        64'h03e30124_01230414,
        64'h4903faf7_69e30ff7,
        64'hf7930094_01a3fff4,
        64'h879b4705_01342e23,
        64'h04444483_29811a09,
        64'h876300f9_e9b30089,
        64'h999b04a4_478304b4,
        64'h4983fee7_91e32000,
        64'h07134107_d79b0107,
        64'h979b8fd9_0087979b,
        64'h03f44703_04044783,
        64'hb78547b5_c1194a01,
        64'hf6e505e3_4785470d,
        64'hbf8500e5_19634785,
        64'h470dfe99_15e30491,
        64'hc10dea1f_f0ef8522,
        64'h85d2000a_07634509,
        64'h0004aa03_01048913,
        64'hff2a14e3_09910941,
        64'h00a9a023_2501c51f,
        64'hf0ef854a_c7894501,
        64'hffc94783_89a623a4,
        64'h0a131fa4_0913848a,
        64'h04f51a63_4785ee5f,
        64'hf0ef8522_4581f571,
        64'h89110009_0463fb79,
        64'h478d0015_77131360,
        64'h60ef00a4_00a30004,
        64'h00230ff4_f5138082,
        64'h6161853e_6ae27a02,
        64'h79a27942_74e26406,
        64'h60a647a9_c1118911,
        64'h00090563_e3850015,
        64'h77932220_60ef0014,
        64'h4503c79d_00044783,
        64'h0089b023_c01547b1,
        64'h84aa6380_97baa567,
        64'h87930000_a7970035,
        64'h17130205_4e6347ad,
        64'hddbff0ef_8932852e,
        64'h89aa0005_3023ec56,
        64'hf052fc26_e0a2e486,
        64'hf44ef84a_715dbfcd,
        64'h450d8082_61056902,
        64'h64a26442_60e200a0,
        64'h35338d05_01257533,
        64'h2501d25f_f0ef0864,
        64'h05130097_8c634501,
        64'h0127f7b3_14650493,
        64'h00544537_fff50913,
        64'h01000537_0005079b,
        64'hd4bff0ef_06a40513,
        64'h02e79f63_a5570713,
        64'h4107d79b_776d0107,
        64'h979b8fd9_0087979b,
        64'h45092324_47032334,
        64'h4783e52d_2501fa3f,
        64'hf0ef842a_d91c0005,
        64'h022357fd_e04ae426,
        64'hec06e822_11018082,
        64'h61056902_64a26442,
        64'h60e28522_0324a823,
        64'h597d4405_c1192501,
        64'h2d6060ef_03448593,
        64'h864a4685_0014c503,
        64'hec190005_041bfddf,
        64'hf0ef892e_84aa02b7,
        64'h87634401_e04ae426,
        64'hec06e822_1101591c,
        64'h80824501_f8dff06f,
        64'hc3990045_4783b7f9,
        64'h4505b7e5_397d34e0,
        64'h60ef85ce_86269cbd,
        64'h46850014_45034c5c,
        64'hff2a74e3_4a050034,
        64'h49038082_61456a02,
        64'h69a26942_64e27402,
        64'h70a24501_00e7eb63,
        64'h40f487bb_00040223,
        64'h4c58505c_e1312501,
        64'h390060ef_85ce8626,
        64'h46850015_4503842a,
        64'h03450993_e052e84a,
        64'hf4065904_e44eec26,
        64'hf0227179_8082853e,
        64'h27818fd5_0107979b,
        64'h8fd10087_179b0145,
        64'hc6030155_c70300e5,
        64'h1d630006_879b8edd,
        64'h0087979b_470d01a5,
        64'hc68301b5_c7838082,
        64'h45258082_014160a2,
        64'h4525c391_45010015,
        64'h77934020_60ef0017,
        64'hc503e406_114102e6,
        64'h90630085_57030067,
        64'hd683c70d_0007c703,
        64'hcb85611c_c915bfd5,
        64'hc5074703_0000a717,
        64'h8082853a_e11c0006,
        64'h871b0789_00b66663,
        64'h0ff6f593_fd06869b,
        64'h577d4605_0007c683,
        64'hb7dd0705_a00d577d,
        64'h00d70663_00178693,
        64'h00c69863_02d5fc63,
        64'h00074683_03a00613,
        64'h02000593_cf99873e,
        64'h611c8082_61056902,
        64'h64a26442_60e20004,
        64'h002300f4_93238fd9,
        64'h0087979b_01694703,
        64'h01794783_00f49223,
        64'h8fd90087_979b0189,
        64'h47030199_4783c088,
        64'hf4bff0ef_00f58423,
        64'h84ae01c9_051300b9,
        64'h4783fcd7_9be30785,
        64'h040500e4_00230405,
        64'h01140023_01031563,
        64'h0007831b_0e500713,
        64'h00a71463_02c70063,
        64'h00074703_00f90733,
        64'h46ad02e0_08934821,
        64'h45150200_06134781,
        64'h01853903_cfb50095,
        64'h8413e04a_e426ec06,
        64'he8221101_495cbfc5,
        64'hfeb50fa3_05058082,
        64'h00f61363_0005079b,
        64'h9e29b7d5_00d70023,
        64'h078500f5_07330007,
        64'h468300f5_87338082,
        64'h00e61363_0007871b,
        64'h47818082_25018d5d,
        64'h05628fd9_07c20035,
        64'h45030025_47838f5d,
        64'h07a20005_47030015,
        64'h4783b7d9_14fdb7e9,
        64'hba7ff0ef_bfc1710a,
        64'h84937c90_50ef4501,
        64'hdff154fd_000a2783,
        64'hbfc5bc1f_f0effc07,
        64'h5de30337_97138309,
        64'h37830207_45630337,
        64'h97138309_37835a0b,
        64'h0493ed1f_e0ef8522,
        64'he78d0009_a783e4a9,
        64'hd807ac23_0000a797,
        64'hda07a223_0000a797,
        64'hda07a823_0000a797,
        64'hda07a423_0000a797,
        64'hda079a23_0000a797,
        64'hdcf70ea3_0000a717,
        64'h00544783_def70423,
        64'h0000a717_00444783,
        64'hdef709a3_0000a717,
        64'h00344783_def70f23,
        64'h0000a717_43001937,
        64'h00262b37_00244783,
        64'he0f708a3_0000a717,
        64'h6a89e02a_0a130000,
        64'haa170014_4783e2f7,
        64'h03230000_a717e0e9,
        64'h89930000_a9974481,
        64'h00044783_e3440413,
        64'h0000a417_09b030ef,
        64'h06050513_00009517,
        64'he485c583_0000a597,
        64'he5164603_0000a617,
        64'he5a6c683_0000a697,
        64'he6584803_0000a817,
        64'he6c7c783_0000a797,
        64'he7374703_0000a717,
        64'h0d7030ef_08c50513,
        64'h00009517_80e7b423,
        64'he05ae456_e852ec4e,
        64'hf04af426_f822fc06,
        64'h8f4d91c1_15c20080,
        64'h07377139_8087b583,
        64'h8007b603_430017b7,
        64'hbf81fd24_1ee31150,
        64'h30ef00c7_80230ff6,
        64'h761300c4_d6330286,
        64'h061b0405_854e0004,
        64'h059b0144_07b3028a,
        64'h863b4919_0d498993,
        64'h00009997_ee4a0a13,
        64'h0000aa17_5ae14401,
        64'h80826161_6ae27a02,
        64'h79a27942_74e282f6,
        64'hb42347a1_640660a6,
        64'h8086b783_8006b783,
        64'h80f6b423_93c180a6,
        64'hb02317c2_91014300,
        64'h16b78fd9_15020ff7,
        64'h77138ff1_83210087,
        64'h179bf006_06130100,
        64'h06374722_f31ff0ef,
        64'h451200f0_50ef0028,
        64'hf4858593_0000a597,
        64'h460901f0_50ef0048,
        64'hf5a58593_0000a597,
        64'h4611f6a7_83a30000,
        64'ha797fe05_6513893d,
        64'h027070ef_f6f70c23,
        64'h0000a717_5791f8f7,
        64'h00a30000_a717578d,
        64'hf8f70523_0000a717,
        64'h5789f8f7_09a30000,
        64'ha7175785_f8f70e23,
        64'h0000a717_57b9ecc5,
        64'hc3110107_9713fff4,
        64'hc7932110_30ef19e5,
        64'h05130000_951784aa,
        64'h099070ef_ec56f052,
        64'hf44ef84a_e0a2fc26,
        64'he486c63e_04b00513,
        64'h45854601_00740207,
        64'h879b0700_07b7715d,
        64'h80822501_8d5d8d79,
        64'h00ff0737_0085151b,
        64'h8fd98f75_0085571b,
        64'hf0068693_8fd966c1,
        64'h0185579b_0185171b,
        64'h80829141_15428d5d,
        64'h05220085_579b8082,
        64'h614564e2_740270a2,
        64'h85228e0f_f0ef02e5,
        64'h05130000_a5170450,
        64'h06930267_57030000,
        64'ha7170228_88930000,
        64'ha89785a6_862247b2,
        64'h0007a803_03c78793,
        64'h0000a797_129050ef,
        64'hf4060068_08458593,
        64'h0000a597_461184ae,
        64'h8432ec26_f0227179,
        64'hbfc14785_ec3ff0ef,
        64'h80826105_64a26442,
        64'h60e2c3c0_0c2007b7,
        64'h2ef030ef_26450513,
        64'h00009517_e7990206,
        64'hc1630337_16938304,
        64'hb7034300_14b74781,
        64'h2401ec06_e42643c0,
        64'he8220c20_07b71101,
        64'h80826101_01135f81,
        64'h34838526_60013403,
        64'h60813083_8287b823,
        64'h430017b7_0405a9bf,
        64'hf0ef8626_fef845e3,
        64'h0006881b_ff063c23,
        64'h06210685_00083803,
        64'h983a0036_98139742,
        64'h85b24681_4037d79b,
        64'h43000837_860a2785,
        64'h0077e793_37ed02d5,
        64'h1e638066_86936685,
        64'hc6918005_069b0001,
        64'h550300d1_00230086,
        64'hd69b0106_d69b0106,
        64'h969b00d1_00a345d4,
        64'h95ba070e_9f318006,
        64'h871b7007_76130084,
        64'h171beb3d_431814e7,
        64'h07130000_a717c349,
        64'h27018f71_fff74713,
        64'h00c5163b_10100513,
        64'h8a1d0905_6c63ffc7,
        64'h849b5f20_0513fee7,
        64'h881b2781_60113423,
        64'h5e913c23_639c97ae,
        64'h430005b7_9fad8406,
        64'h879b0387_f5930034,
        64'h179b6685_8387b703,
        64'h00f67413_26016081,
        64'h30239f01_01138307,
        64'hb6034300_17b7bba5,
        64'h46014210_30ef37e5,
        64'h05130000_951785aa,
        64'hb36900f4_16236080,
        64'h079300f4_1f230024,
        64'hd78300f4_1e230004,
        64'hd78302f4_142301e4,
        64'h578302f4_132302a0,
        64'h061301c4_57832cb0,
        64'h50ef8522_85ca4619,
        64'h2d5050ef_00640513,
        64'h21858593_0000a597,
        64'h46192e70_50ef854e,
        64'h22858593_0000a597,
        64'h46192f70_50ef854a,
        64'h85ce4619_00f59a23,
        64'h01658993_02058913,
        64'h20000793_eaf719e3,
        64'h26a7d783_0000a797,
        64'h0285d703_ecf711e3,
        64'h27848493_0000a497,
        64'h2807d783_0000a797,
        64'h0265d703_b1e93f65,
        64'h05130000_9517b9d1,
        64'h3e850513_00009517,
        64'hb9f93c25_05130000,
        64'h9517b1e5_3ac50513,
        64'h00009517_b9cd39e5,
        64'h05130000_9517b9f5,
        64'h38050513_00009517,
        64'hb31937a5_05130000,
        64'h9517bb01_36450513,
        64'h00009517_bb293565,
        64'h05130000_9517b315,
        64'h34050513_00009517,
        64'hb33d33a5_05130000,
        64'h9517b799_3a9050ef,
        64'h08683025_85930000,
        64'ha5974611_f4f70de3,
        64'h02045703_f6f701e3,
        64'h17fd67c1_01e45703,
        64'hf6e787e3_5fe00713,
        64'hbf95cb4f_f0ef02a4,
        64'h051385ca_573030ef,
        64'h36050513_00009517,
        64'hccaff0ef_852285a6,
        64'h587030ef_36450513,
        64'h00009517_02e79863,
        64'h4d200713_b765d73f,
        64'he0ef02a4_05133465,
        64'h85930000_a5973426,
        64'h06130000_a6173466,
        64'h86930000_a697f7e9,
        64'h439c3527_87930000,
        64'ha797c799_439c3627,
        64'h87930000_a79734f7,
        64'h2f230000_a71747e2,
        64'h04e69463_04300713,
        64'h80826161_79a27942,
        64'h74e26406_60a65a00,
        64'h60ef4501_02a40593,
        64'hff89061b_37478793,
        64'h0000a797_66a24762,
        64'h47d050ef_e43638f7,
        64'h2f230000_a71739e5,
        64'h05130000_a5173965,
        64'h85930000_a5974619,
        64'h47e23ad7_9f230000,
        64'ha79704e7_9b6301c1,
        64'h56830450_071300e1,
        64'h0e230234_470300e1,
        64'h0ea301c1_19030224,
        64'h470300e1_0e232781,
        64'h02744703_00e10ea3,
        64'h01c11783_00f10e23,
        64'h02544783_00f10ea3,
        64'h02644703_02444783,
        64'hbdbd44a5_05130000,
        64'h9517b561_43c50513,
        64'h00009517_bd4942e5,
        64'h05130000_9517a06d,
        64'hdcdfe0ef_450185a2,
        64'h862602a4_122300a1,
        64'h1e238d5d_05220085,
        64'h579bdb3f_f0ef00f4,
        64'h1e230029_d78300f4,
        64'h1d230009_d78302f4,
        64'h10230224_0513fde4,
        64'h859b01c4_578300f4,
        64'h1f230204_12230204,
        64'h012301a4_578355b0,
        64'h50ef854a_49c58593,
        64'h0000a597_461956b0,
        64'h50ef8522_85ca4619,
        64'h10f71b63_4ce7d783,
        64'h0000a797_02045703,
        64'h12f71363_4dc98993,
        64'h0000a997_4e47d783,
        64'h0000a797_01e45703,
        64'hb73d62a5_05130000,
        64'h9517f0f5_9ce30880,
        64'h079326f5_88630ff0,
        64'h079326f5_87630890,
        64'h0793b73d_f4f58ae3,
        64'h62050513_00009517,
        64'h06c00793_26f58a63,
        64'h06700793_00b7ef63,
        64'h28f58563_08400793,
        64'hbf91f6f5_8de360e5,
        64'h05130000_951705e0,
        64'h079328f5_836305c0,
        64'h0793b7bd_f8f58ae3,
        64'h5f850513_00009517,
        64'h03200793_28f58663,
        64'h02f00793_00b7ef63,
        64'h2af58163_03300793,
        64'h04b7e263_2cf58163,
        64'h06200793_b7c95f65,
        64'h05130000_9517faf5,
        64'h96e30290_07932af5,
        64'h85630210_0793bf6d,
        64'hfef580e3_5dc50513,
        64'h00009517_47d916f5,
        64'h896347c5_00b7ed63,
        64'h2cf58163_47f5a429,
        64'h7ff030ef_fef591e3,
        64'h5c050513_00009517,
        64'h47a118f5_81634799,
        64'ha4150180_40ef7565,
        64'h05130000_951702f5,
        64'h83635ba5_05130000,
        64'h95174789_10f58463,
        64'h478502b7_e3631af5,
        64'h82634791_04b7e563,
        64'h1cf58163_47b108b7,
        64'he76332f5_886302e0,
        64'h07930174_45836cb0,
        64'h50ef5d25_05130000,
        64'ha5174619_85ca0064,
        64'h09136df0_50ef4611,
        64'h082884b2_05e94407,
        64'h99638005_079b0af5,
        64'h0e636dd7_879367a1,
        64'h3cf50463_842e8067,
        64'h8793f44e_f84afc26,
        64'he486e0a2_6785715d,
        64'hbf45943e_93c117c2,
        64'h00f11723_8fd90087,
        64'h979b0087_d71b0489,
        64'h00c15783_731050ef,
        64'h00684609_85a68082,
        64'h61459141_694264e2,
        64'h1542fff5_45137402,
        64'h70a29522_01045513,
        64'h942a9041_14420104,
        64'h551302f0_44634099,
        64'h07bb00a5_893b4401,
        64'h84aaf406_e84aec26,
        64'hf0227179_80826365,
        64'h05130000_9517bf75,
        64'h68050513_00009517,
        64'h84078793_fce608e3,
        64'h68050513_00009517,
        64'h83878713_bfe966e5,
        64'h05130000_95178287,
        64'h879300c7_4963fee6,
        64'h09e36925_05130000,
        64'h95178307_87138082,
        64'hfaf612e3_67450513,
        64'h00009517_81878793,
        64'h00e60a63_67450513,
        64'h00009517_81078713,
        64'h80820141_6d450513,
        64'h0000a517_60a21600,
        64'h40efe406_6e450513,
        64'h0000a517_71458593,
        64'h00009597_9e3d1141,
        64'h7c07879b_77fd04c7,
        64'hc9637225_05130000,
        64'h951787f7_87936785,
        64'hc3ad6a25_05130000,
        64'h95178006_079b04c7,
        64'h496306e6_0b636c65,
        64'h05130000_95178087,
        64'h871308a7_4463862a,
        64'h0ce50763_82078713,
        64'h67858082_953e057e,
        64'h450597aa_20000537,
        64'he3089536_00178693,
        64'h00756513_157d631c,
        64'h78070713_0000a717,
        64'h80824000_05378082,
        64'h057e4505_bfb12405,
        64'h03e060ef_854a4581,
        64'h86262280_40ef855e,
        64'h85ca993e_86268c9d,
        64'h79020097_ff6377a2,
        64'h74c29982_85260009,
        64'h061b45c2_24a040ef,
        64'h856a86ca_85a66642,
        64'h8082612d_6d0a6caa,
        64'h6c4a6bea_7b0a7aaa,
        64'h7a4a79ea_690e64ae,
        64'h644e60ee_55752740,
        64'h40ef71a5_05130000,
        64'h951785a6_0397e863,
        64'h018487b3_74820409,
        64'h08637922_292040ef,
        64'h855a85a2_cfbd77c2,
        64'h09579263_47a29982,
        64'h9dbd0028_03800613,
        64'h7786028a_05bba091,
        64'h656600f4_64630781,
        64'h578377ad_0d130000,
        64'h9d170800_0cb78000,
        64'h0c377a2b_8b930000,
        64'h9b9776ab_0b130000,
        64'h9b174a85_03800a13,
        64'h440106e7_9d635579,
        64'h83e107e2_631868e7,
        64'h07130000_a7176786,
        64'h9982e16a_e566e962,
        64'hed5ef15a_f556f952,
        64'he1cae5a6_e9a2ed86,
        64'h00884581_89aa0400,
        64'h0613fd4e_7115bfd5,
        64'h8f8d2505_8082e21c,
        64'h00b7f463_45019181,
        64'h87aa1582_b70d0705,
        64'h27850117_00230006,
        64'h54634186_561b0186,
        64'h161bc519_09757513,
        64'h00054503_00cc0533,
        64'h00074603_bfdd4781,
        64'hbf253cfd_fe97eae3,
        64'h27856782_136070ef,
        64'he03e855e_b76500c5,
        64'h80230ff6_761395be,
        64'h082c0007_4603bf6d,
        64'h00c59023_95aa9241,
        64'h16420828_00179593,
        64'h00075603_011d1d63,
        64'hbfd1e190_95aa0828,
        64'h00379593_6310010d,
        64'h1963bf9d_46914821,
        64'h07859752_488967a2,
        64'h67023c80_40efe03a,
        64'he43e855a_85d69201,
        64'h1602c190_95aa2601,
        64'h08280027_95934310,
        64'h02dd1963_b79d557d,
        64'hd13d10a0_70ef9936,
        64'h92811682_41b4043b,
        64'h66824000_40effa07,
        64'h8c23e036_89450513,
        64'h0000a517_97ba1098,
        64'h0b079c63_0006881b,
        64'h02e00893_85ba4781,
        64'h083803bd_06bb0d9d,
        64'he56399be_034787b3,
        64'h9381020d_979305b6,
        64'h6b630007_861b4889,
        64'h48214691_4781874e,
        64'h000c8d9b_008cf463,
        64'h00040d9b_45a040ef,
        64'h8d850513_0000a517,
        64'h85ca8082_61697da6,
        64'h7d467ce6_6c0a6baa,
        64'h6b4a6aea_7a0a79aa,
        64'h794a74ea_640e60ae,
        64'h4501e00d_7dcc0c13,
        64'h00008c17_884b8b93,
        64'h0000ab97_91cb0b13,
        64'h0000ab17_020a5a13,
        64'h001a849b_020d1a13,
        64'h001d1a9b_03acdcbb,
        64'h4cc1000c_956302cc,
        64'hdcbb0400_0c9300e7,
        64'hf6638436_8d3289ae,
        64'h892a0400_0793f4ee,
        64'he162e55e_e95aed56,
        64'hf152fd26_e586f8ea,
        64'hf54ef94a_e1a202c7,
        64'h073b8cba_fce67155,
        64'h4f60406f_610596e5,
        64'h05130000_a51764a2,
        64'h690285a6_864a60e2,
        64'h64425100_40ef9665,
        64'h05130000_a51785a2,
        64'hc8015200_40ef8932,
        64'h97050513_0000a517,
        64'h85be0785_14590087,
        64'h74630104_5433942a,
        64'h472500d4_14334405,
        64'h03b6869b_02e50533,
        64'h4729c10d_44018d79,
        64'hfff74713_01071733,
        64'h577db7f5_9c450513,
        64'h0000a517_85aafab7,
        64'h1ce32705_5720406f,
        64'h61059da5_05130000,
        64'ha51785aa_690264a2,
        64'h60e26442_e495e04a,
        64'he822ec06_00074483,
        64'he426972e_11019765,
        64'h85930000_b5979301,
        64'h1702cf85_00f557b3,
        64'h883e03c6_879b02e8,
        64'h86bb4599_58d94701,
        64'h862ebfa1_9fc50513,
        64'h0000a517_85aabf55,
        64'h4401bf51_843a0086,
        64'hf46302f4_5733bf61,
        64'h02e45433_5e20406f,
        64'h6105a425_05130000,
        64'ha5176902_64a285ca,
        64'h862660e2_64425fc0,
        64'h40efa525_05130000,
        64'ha51785a2_c80160c0,
        64'h40ef84b2_a5c50513,
        64'h0000a517_943e0014,
        64'h44130324_341302e4,
        64'h743302f4_57b30640,
        64'h07130087_7d630630,
        64'h0713cf39_02f47733,
        64'h46a547a9_0687e263,
        64'h47293e80_0793c815,
        64'h02f555b3_02f57433,
        64'hbf7d2407_87934685,
        64'hb7d9a007_87934681,
        64'h6660406f_6105aa65,
        64'h05130000_a51785aa,
        64'h690264a2_60e26442,
        64'h02091663_e426e822,
        64'hec060007_4903e04a,
        64'h97361101_a7470713,
        64'h0000b717_3e800793,
        64'h46890ca7_fc633e70,
        64'h079304a7_676323f7,
        64'h8713000f_47b704a7,
        64'h6963862e_9ff78713,
        64'h3b9ad7b7_8082612d,
        64'h450160ee_6ca040ef,
        64'hb0050513_0000a517,
        64'h002cfebf_f0efed86,
        64'h45050c80_0613002c,
        64'h7115f73f_f06f4581,
        64'h862e86b2_80826145,
        64'h69a26942_64e2854a,
        64'h740270a2_2bc060ef,
        64'hb1858593_0000a597,
        64'h00890533_ffd4841b,
        64'h00f44463_ffe4879b,
        64'h9c296e00_40ef954a,
        64'hb4860613_0000a617,
        64'h86ce40a4_85bb0095,
        64'h5d630009_8f63842a,
        64'h6fe040ef_854a85a6,
        64'hb6060613_0000a617,
        64'h01870713_00009717,
        64'hb6868693_0000a697,
        64'hc5093ba6_86930000,
        64'ha6978932_89ae84b6,
        64'hf022f406_e44ee84a,
        64'hec267179_bfdd77c0,
        64'h40ef8562_b7f10905,
        64'h786040ef_856600fb,
        64'he7630ff7_f793fe05,
        64'h879b0007_c5830129,
        64'h87b3bf15_04857a40,
        64'h40ef7325_05130000,
        64'ha51700f4_5a630009,
        64'h079b4124_093b7bc0,
        64'h40ef00f4_f913855a,
        64'hff2dcce3_2d857cc0,
        64'h40ef8552_bfdd7d40,
        64'h40ef8562_b75d0905,
        64'h7de040ef_856600fb,
        64'he7630ff7_f793fe05,
        64'h879b0007_c5830129,
        64'h87b3a805_00f97913,
        64'h4d81fffd_4913068d,
        64'h12630090_40efc165,
        64'h05130000_a5170007,
        64'hc5830099_87b301d0,
        64'h40ef8552_023040ef,
        64'h7b050513_0000a517,
        64'h02879d63_0009079b,
        64'hff048913_03b040ef,
        64'h855ae39d_00f47793,
        64'hc01d8082_61656da2,
        64'h6d426ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h694664e6_740670a6,
        64'h03544163_0004841b,
        64'hfff58d1b_c6cc8c93,
        64'h0000ac97_c7cc0c13,
        64'h0000ac17_06000b93,
        64'hc70b0b13_0000ab17,
        64'h940a0a13_0000ba17,
        64'h44818aae_89aae46e,
        64'he8caf0a2_f486e86a,
        64'hec66f062_f45ef85a,
        64'hfc56e0d2_e4ceeca6,
        64'h7159b7cd_0bb040ef,
        64'he007a823_0000b797,
        64'hc9850513_0000a517,
        64'h80826151_641260b2,
        64'h85220d90_40efc7e5,
        64'h05130000_a517c565,
        64'h85930000_a597860a,
        64'hc10d842a_e01ff0ef,
        64'h85220f90_40efc765,
        64'h05130000_a517c765,
        64'h85930000_a597842a,
        64'h00054603_00154683,
        64'h00254703_00354783,
        64'h00454803_00554883,
        64'he222e606_716d8082,
        64'h616569a6_694664e6,
        64'h74064501_70a67f01,
        64'h01138ddf_f0ef86c6,
        64'h85a61808_56326882,
        64'hfc4ff0ef_03e10513,
        64'h863e86c2_85a267c2,
        64'h6822f94f_f0efd64e,
        64'h05210513_85a2864a,
        64'h86ba943e_7fc40413,
        64'h6762747d_97ba8107,
        64'h87931018_67857f20,
        64'h60efd602_e83eec3a,
        64'he4428936_89b2e046,
        64'h05a10513_84aa8101,
        64'h0113e4ce_e8caeca6,
        64'hf0a2f486_71591ad0,
        64'h406fd125_05130000,
        64'ha51785aa_80826125,
        64'h7aa27a42_79e26906,
        64'h64a66446_450160e6,
        64'h911a6305_96fff0ef,
        64'h85ce86a6_10084652,
        64'h855ff0ef_460156fd,
        64'h02e10513_85a2821f,
        64'hf0ef0440_06130430,
        64'h06930421_051385a2,
        64'h943e1451_978a020a,
        64'h879312f1_1c233537,
        64'h87936799_12f11b23,
        64'h26378793_77e108b0,
        64'h60ef04f1_06230661,
        64'h05134641_479985ce,
        64'h04f11523_10100793,
        64'h057060ef_ca3e04a1,
        64'h05134581_0f000613,
        64'h0fc00793_0b9060ef,
        64'h000107a3_15410223,
        64'h14f101a3_14510513,
        64'h460585ca_57fd0d30,
        64'h60ef13f1_05134611,
        64'h95beff04_0593978a,
        64'h020a8793_12f10f23,
        64'h479112f1_0ea30370,
        64'h07930f70_60ef0141,
        64'h07a31a68_460585ca,
        64'h993e978a_020a8793,
        64'h12f11d23_13500793,
        64'hc83e4a05_fef40913,
        64'h439ce827_87930000,
        64'hb7970d90_60ef8526,
        64'h55fd4619_94beff84,
        64'h0493978a_020a8793,
        64'h747d2d10_40efca02,
        64'h6a85e225_05130000,
        64'ha517911a_89aaf456,
        64'hf852fc4e_e0cae4a6,
        64'he8a2ec86_711d737d,
        64'hb34d2f90_40efe0e5,
        64'h05130000_a517bf45,
        64'he0850513_0000a517,
        64'h95be978a_d0040593,
        64'h35078793_678531d0,
        64'h40efe025_05130000,
        64'ha5173290_40efdfe5,
        64'h05130000_a51700fa,
        64'h20234785_de0794e3,
        64'h000a2783_b3fd3450,
        64'h40efe0a5_05130000,
        64'ha517bbf5_353040ef,
        64'he0050513_0000a517,
        64'h95be978a_f0040593,
        64'h35048793_36b040ef,
        64'he0850513_0000a517,
        64'h95bee004_0593978a,
        64'h35048793_383040ef,
        64'h02f5d5bb_e107879b,
        64'h678502f6_763b02f5,
        64'hf6bb02f5_d63b03c0,
        64'h079314f7_1e230000,
        64'hb7170121_578316f7,
        64'h13230000_b717e2e5,
        64'h05130000_a51755c2,
        64'h01015783_3c3040ef,
        64'he2050513_0000a517,
        64'h01014583_01114603,
        64'h01214683_01314703,
        64'h3df040ef_e1c50513,
        64'h0000a517_01814583,
        64'h01914603_01a14683,
        64'h01b14703_3fb040ef,
        64'h00b14703_1cf71323,
        64'h0000b717_e1c50513,
        64'h0000a517_00814583,
        64'h35215783_1cf71e23,
        64'h0000b717_00914603,
        64'h00a14683_35015783,
        64'h42f040ef_e1c50513,
        64'h0000a517_35014583,
        64'h35114603_35214683,
        64'h35314703_2b9060ef,
        64'h01490593_4611953e,
        64'hcb840513_978a3504,
        64'h87936485_2d1060ef,
        64'h0e880109_05934611,
        64'h46f040ef_e4c50513,
        64'h0000a517_00fa2023,
        64'h47851207_9a63000a,
        64'h2783b321_d00d0023,
        64'h2fd060ef_9d228562,
        64'h866ab749_cc048513,
        64'hbb39cef4_2023401c,
        64'h00f41023_8fd90087,
        64'h979b0087_d71bce24,
        64'h578300f4_11238fd9,
        64'h0087979b_0087d71b,
        64'hce045783_339060ef,
        64'h4611953e_ce048513,
        64'h978a3507_87936785,
        64'hbfdd855a_4611b395,
        64'h355060ef_85564611,
        64'hb3bdf00d_00233630,
        64'h60ef9d22_953e866a,
        64'hf0048513_978a3507,
        64'h87936785_a00d953e,
        64'h978a3507_87936785,
        64'h4611cd04_85138082,
        64'h3b010113_35013d03,
        64'h35813c83_36013c03,
        64'h36813b83_37013b03,
        64'h37813a83_38013a03,
        64'h38813983_39013903,
        64'h39813483_3a013403,
        64'h3a813083_911a6305,
        64'hcf3ff0ef_0e8885de,
        64'h86ca5672_bd9ff0ef,
        64'h35e10513_85a24601,
        64'h56fdba5f_f0ef3721,
        64'h051385a2_04400613,
        64'h04300693_943ecec4,
        64'h0413978a_350a8793,
        64'h46f11423_35378793,
        64'h679946f1_13232637,
        64'h879377e1_411060ef,
        64'h36f10e23_39610513,
        64'h85de4799_464136f1,
        64'h1d231010_07933dd0,
        64'h60efde3e_37a10513,
        64'h45810f00_06131020,
        64'h079343f0_60ef4731,
        64'h0d230001_03a346f1,
        64'h0ca347b1_051385a6,
        64'h460557fd_459060ef,
        64'h47410a23_47510513,
        64'h461195be_cf440593,
        64'h978a350a_879346f1,
        64'h09a30360_079347b0,
        64'h60ef4741_072346f1,
        64'h05134611_4a1195be,
        64'hcf040593_978a350a,
        64'h879346f1_06a30320,
        64'h079349f0_60efc0d2,
        64'h46c10513_85a64605,
        64'h94becb74_0493c2a6,
        64'h978a350a_879346f1,
        64'h15231350_079300f1,
        64'h03a3478d_47b060ef,
        64'h854a55fd_4619993e,
        64'hcf840913_978a350a,
        64'h87936710_40efde02,
        64'h54e25a52_03c50513,
        64'h0000a517_4f1060ef,
        64'h953e4611_01490593,
        64'hce840513_978a350a,
        64'h87935070_60ef013c,
        64'ha023953e_46110109,
        64'h0593ce44_05134985,
        64'h978a350a_87936a85,
        64'h16079263_000ca783,
        64'h3af59f63_478938f5,
        64'h83634799_24f58363,
        64'h747d4795_00614583,
        64'hf8e79ce3_0ff00713,
        64'h24e78563_03800713,
        64'haac94605_cb648513,
        64'hfae798e3_03500713,
        64'h20e78e63_03300713,
        64'h00f76e63_22e78163,
        64'h03600713_b769e00d,
        64'h002357f0_60ef9d22,
        64'h953e866a_e0048513,
        64'h978a3507_87936785,
        64'hfee794e3_473d22e7,
        64'h83634731_bf4d7350,
        64'h40ef2625_05130000,
        64'ha51785be_22e78763,
        64'hcc848513_470d2ae7,
        64'h89634705_02f76263,
        64'h22e78f63_471904f7,
        64'h6b6326e7_8b6301a9,
        64'h89bb0589_02a00713,
        64'h29890f07_c7830015,
        64'hcd030139_07b395ca,
        64'h0f098593_9c3a9b3a,
        64'h49818a36_8cb28bae,
        64'hd0048c13_cb848b13,
        64'h970a3507_87139aba,
        64'hcd848a93_970a3507,
        64'h871374fd_678524f7,
        64'h1d634789_00054703,
        64'ha0017b90_40ef15e5,
        64'h05130000_a51785aa,
        64'h00e7ea63_892a5800,
        64'h073797aa_d0040023,
        64'hf0040023_e0040023,
        64'hca040b23_ce042023,
        64'hd00007b7_943e747d,
        64'h978a911a_35078793,
        64'h35a13823_35913c23,
        64'h37813023_37713423,
        64'h37613823_37513c23,
        64'h39413023_39313423,
        64'h38913c23_3a113423,
        64'h39213823_3a813023,
        64'h6785737d_c5010113,
        64'hfadff06f_614564e2,
        64'h00e4859b_70a27402,
        64'h852200f4_162347a1,
        64'h6b5060ef_85b64619,
        64'h852266a2_6c1060ef,
        64'he436f406_46190519,
        64'h84b2842a_ec26f022,
        64'h71798082_01416402,
        64'h60a28522_fa1ff0ef,
        64'he4064501_85aa8622,
        64'h0005841b_e0221141,
        64'hbfe10505_01173023,
        64'h97369742_0008b883,
        64'h00e588b3_00351713,
        64'h808280c6_b82396be,
        64'h678500f7_47630005,
        64'h071b6805_450102e7,
        64'hc7bb2785_0077e793,
        64'hfff6079b_8007bc23,
        64'h97b64721_67856394,
        64'h4b878793_0000b797,
        64'h80826145_740270a2,
        64'h00f41523_fff7c793,
        64'h9fb94107_d71b9fb9,
        64'h93411742_4107579b,
        64'hfed79ce3_9f31ffe7,
        64'hd6030789_470187a2,
        64'h01440693_779060ef,
        64'h01040513_002c4611,
        64'h785060ef_00c40513,
        64'h00041523_006c4611,
        64'h00f404a3_47c579b0,
        64'h60efec3e_00840513,
        64'h00041323_082c4621,
        64'h47c17af0_60ef0044,
        64'h05130161_05934609,
        64'h7bd060ef_00f11b23,
        64'hc4360509_084c57fd,
        64'h460900f1_1a238fd9,
        64'h0087979b_0ff77713,
        64'h0087d713_c632842a,
        64'h419c00f5_10230457,
        64'h879b6785_c19c27d1,
        64'hf022f406_7179419c,
        64'h80820005_132300f5,
        64'h122300d5_112300c5,
        64'h10238fd9_0087979b,
        64'h0ff77713_c19c0087,
        64'hd7138ed9_06a20086,
        64'hd71b8e59_27a10622,
        64'h0086571b_419cc19c,
        64'h2785c319_0017f713,
        64'h419cbfcd_fda00513,
        64'h80826121_74a27442,
        64'h70e29782_85a66562,
        64'h701ce509_c39ff0ef,
        64'h842a0830_65a2c105,
        64'hc7dff0ef_84b2e42e,
        64'hf822fc06_f4267139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2655c,
        64'h862686ca_6562e519,
        64'hc75ff0ef_083065a2,
        64'hc115cb7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hbfc5fda0_05138082,
        64'h61217902_74a27442,
        64'h70e29782_85a2615c,
        64'h862686ca_6562e519,
        64'hcb5ff0ef_083065a2,
        64'hc115cf7f_f0ef893a,
        64'h84b68432_e42efc06,
        64'hf04af426_f8227139,
        64'hb7e16522_f569cdbf,
        64'hf0ef8526_85ce0030,
        64'hbfc90284_8493c501,
        64'h6d3060ef_854a608c,
        64'h2a6050ef_855285ca,
        64'h60908082_61216a42,
        64'h69e27902_74a27442,
        64'h70e24501_00849b63,
        64'h942602f4_043345ea,
        64'h0a130000_aa1789ae,
        64'h892afc06_e852ec4e,
        64'hf04a0280_079302f4,
        64'h043b840d_8c0574e4,
        64'h84930000_b4977564,
        64'h04130000_b417f426,
        64'hf822639c_69478793,
        64'h0000b797_7139bfdd,
        64'h45018082_61056442,
        64'h60e2fda0_05138302,
        64'h610560e2_65a26442,
        64'h85220003_0e630205,
        64'h3303c919_db9ff0ef,
        64'he42eec06_4108842a,
        64'he8221101_bfc56562,
        64'hf96dd97f_f0ef0830,
        64'h80826145_70a24501,
        64'he50965a2_de1ff0ef,
        64'hf406e42e_7179bfc1,
        64'h5479fcf7_1be30ff0,
        64'h079300c7_c70367a2,
        64'h130080ef_6522f565,
        64'h842adcff_f0ef85a6,
        64'h00308522_80826145,
        64'h64e27402_70a28522,
        64'h543515c0_80ef51e5,
        64'h05130000_a51700f4,
        64'hcf63445c_3aa050ef,
        64'h52050513_0000a517,
        64'h85a6842a_c11dfda0,
        64'h0413e47f_f0ef84ae,
        64'hf406ec26_f0227179,
        64'h80826145_694264e2,
        64'h740270a2_85221960,
        64'h80ef6522_3e2050ef,
        64'h54850513_0000a517,
        64'h864a608c_ed01842a,
        64'he45ff0ef_84aa85ca,
        64'h0030c11d_fda00413,
        64'he8dff0ef_892eec26,
        64'hf406e84a_f0227179,
        64'hb7d92405_1d4080ef,
        64'h65224200_50ef854e,
        64'h85a20127_896300c7,
        64'hc78367a2_ed09e83f,
        64'hf0ef8526_85a20030,
        64'h80826121_69e27902,
        64'h74a27442_70e200f4,
        64'h496344dc_5a498993,
        64'h0000a997_0ff00913,
        64'h440184aa_cd01eebf,
        64'hf0efec4e_f04af426,
        64'hf822fc06_7139bfd5,
        64'h54798082_61457402,
        64'h70a28522_23a080ef,
        64'h00f70963_00c54703,
        64'h0ff00793_6562e911,
        64'h842aee7f_f0ef0830,
        64'h65a2c105_fda00413,
        64'hf2dff0ef_e42ef406,
        64'hf0227179_b7c1fda0,
        64'h0513bf65_24052740,
        64'h80ef4981_65224c40,
        64'h50ef8552_00099563,
        64'h2485cb99_0087c783,
        64'h67a2ed19_f29ff0ef,
        64'h854a85a2_00308082,
        64'h61216a42_69e27902,
        64'h74a27442_70e25535,
        64'he0914501_00f44d63,
        64'h00c92783_48ca0a13,
        64'h0000ba17_44014481,
        64'h4985892a_cd31f9bf,
        64'hf0efe852_ec4ef04a,
        64'hf426f822_fc067139,
        64'hbfe54501_80820141,
        64'h60a26108_c509fbbf,
        64'hf0efe406_1141b7f5,
        64'h02870713_fea68de3,
        64'h47148082_853a4701,
        64'h00e79563_97ba02d7,
        64'h87b30280_069302d7,
        64'h87bb878d_8f999c67,
        64'h87930000_c7976294,
        64'h9d070713_0000c717,
        64'h90868693_0000c697,
        64'hb7edfda0_07138302,
        64'h853e85b2_00030563,
        64'h01853303_8082853a,
        64'he21c97b6_470102a7,
        64'h87b30a00_051300b7,
        64'hd963454c_0005cc63,
        64'h5735c285_87ae6914,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h000a2e2e_2e746e65,
        64'h6d6f6d20_61207469,
        64'h61772065_7361656c,
        64'h50202165_6e616972,
        64'h41206d6f_7266206f,
        64'h6c6c6548_ffdff06f,
        64'h10500073_34102373,
        64'h342022f3_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_03f090ef,
        64'hfec5c6e3_02058593,
        64'h0005bc23_0005b823,
        64'h0005b423_0005b023,
        64'h3b860613_0000c617,
        64'hc2058593_0000c597,
        64'h30579073_09078793,
        64'h00000797_00078067,
        64'h40b787b3_00d787b3,
        64'h01478793_00000797,
        64'hfcc5cce3_02068693,
        64'h02058593_00e6bc23,
        64'h0185b703_00e6b823,
        64'h0105b703_00e6b423,
        64'h0085b703_00e6b023,
        64'h0005b703_0006b703,
        64'hff810113_01b11113,
        64'h0110011b_fe0e9ae3,
        64'h0085b703_fffe8e93,
        64'h0005b703_240e8e9b,
        64'h000f4eb7_01169693,
        64'h3ff6869b_000046b7,
        64'hbb560613_0000c617,
        64'hfb058593_00000597,
        64'h000280e7_13050513,
        64'h00000517_0f428293,
        64'h00008297_000280e7,
        64'h0ce28293_00008297,
        64'h01111113_3ff1011b,
        64'h00004137_fe0e9ee3,
        64'hfffe8e93_710e8e9b,
        64'h00002eb7_11249c63,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
