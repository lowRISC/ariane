/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'h011111133ff1011b0000413711249463, /*    1 */
128'h00008297000280e70922829300008297, /*    2 */
128'h000280e713050513000005170b828293, /*    3 */
128'ha1c606130000c617fc05859300000597, /*    4 */
128'h000f4eb7011696933ff6869b000046b7, /*    5 */
128'h0085b703fffe8e930005b703240e8e9b, /*    6 */
128'hff81011301b111130110011bfe0e9ae3, /*    7 */
128'h0085b70300e6b0230005b7030006b703, /*    8 */
128'h0185b70300e6b8230105b70300e6b423, /*    9 */
128'hfcc5cce3020686930205859300e6bc23, /*   10 */
128'h40b787b300d787b30147879300000797, /*   11 */
128'h30579073090787930000079700078067, /*   12 */
128'h1c8606130000c617a30585930000c597, /*   13 */
128'h0005bc230005b8230005b4230005b023, /*   14 */
128'h020004b769a090effec5c6e302058593, /*   15 */
128'h02000937004484930124a02300100913, /*   16 */
128'h3440297310500073ff24c6e34009091b, /*   17 */
128'hf1402973020004b7fe090ae300897913, /*   18 */
128'h0004a903000920230099093300291913, /*   19 */
128'h4009091b0200093700448493fe091ee3, /*   20 */
128'h1050007334102373342022f3ff24c6e3, /*   21 */
128'h41206d6f7266206f6c6c6548ffdff06f, /*   22 */
128'h617720657361656c502021656e616972, /*   23 */
128'h000a2e2e2e746e656d6f6d2061207469, /*   24 */
128'h00000000000000000000000000000000, /*   25 */
128'h00000000000000000000000000000000, /*   26 */
128'h00000000000000000000000000000000, /*   27 */
128'h00000000000000000000000000000000, /*   28 */
128'h00000000000000000000000000000000, /*   29 */
128'h00000000000000000000000000000000, /*   30 */
128'h00000000000000000000000000000000, /*   31 */
128'hd963454c0005cc635735c28587ae6914, /*   32 */
128'he21c97b6470102a787b30a00051300b7, /*   33 */
128'h853e85b200030563018533038082853a, /*   34 */
128'h6f8686930000b697b7edfda007138302, /*   35 */
128'h87930000c7976294824707130000c717, /*   36 */
128'h87b30280069302d787bb878d8f9981a7, /*   37 */
128'h47148082853a470100e7956397ba02d7, /*   38 */
128'hf0efe4061141b7f502870713fea68de3, /*   39 */
128'hbfe545018082014160a26108c509fbbf, /*   40 */
128'hf0efe852ec4ef04af426f822fc067139, /*   41 */
128'h0000ba17440144814985892acd31f9bf, /*   42 */
128'hc091553500f44d6300c9278327ca0a13, /*   43 */
128'h61216a4269e2790274a2744270e24501, /*   44 */
128'h67a2ed19f29ff0ef854a85a200308082, /*   45 */
128'h50ef8552000995632485cb990087c783, /*   46 */
128'h0513bf652405228080ef498165224a60, /*   47 */
128'hf2dff0efe42ef406f0227179b7c1fda0, /*   48 */
128'h842aee7ff0ef083065a2c105fda00413, /*   49 */
128'h00f7096300c547030ff007936562e911, /*   50 */
128'h547980826145740270a285221ee080ef, /*   51 */
128'hf0efec4ef04af426f822fc067139bfd5, /*   52 */
128'h0000a9970ff00913440184aacd01eebf, /*   53 */
128'h74a2744270e200f4496344dc39498993, /*   54 */
128'hf0ef852685a200308082612169e27902, /*   55 */
128'h85a20127896300c7c78367a2ed09e83f, /*   56 */
128'hb7d92405188080ef6522402050ef854e, /*   57 */
128'he8dff0ef892eec26f406e84af0227179, /*   58 */
128'he45ff0ef84aa85ca0030c11dfda00413, /*   59 */
128'h338505130000a517864a608ced01842a, /*   60 */
128'h740270a2852214a080ef65223c4050ef, /*   61 */
128'hf406ec26f022717980826145694264e2, /*   62 */
128'h85a6842ac11dfda00413e47ff0ef84ae, /*   63 */
128'hcf63445c38c050ef310505130000a517, /*   64 */
128'h5435110080ef30e505130000a51700f4, /*   65 */
128'h003085228082614564e2740270a28522, /*   66 */
128'h0e4080ef6522f565842adcfff0ef85a6, /*   67 */
128'h5479fcf71be30ff0079300c7c70367a2, /*   68 */
128'he50965a2de1ff0eff406e42e7179bfc1, /*   69 */
128'hf96dd97ff0ef08308082614570a24501, /*   70 */
128'he42eec064108842ae8221101bfc56562, /*   71 */
128'h852200030e6302053303c919db9ff0ef, /*   72 */
128'h60e2fda005138302610560e265a26442, /*   73 */
128'h0000b7977139bfdd4501808261056442, /*   74 */
128'h04130000b417f426f822639c48478793, /*   75 */
128'h043b840d8c055a2484930000b4975aa4, /*   76 */
128'h892afc06e852ec4ef04a0280079302f4, /*   77 */
128'h942602f4043324ea0a130000aa1789ae, /*   78 */
128'h69e2790274a2744270e2450100849b63, /*   79 */
128'h288050ef855285ca6090808261216a42, /*   80 */
128'hbfc902848493c501695060ef854a608c, /*   81 */
128'hb7e16522f569cdbff0ef852685ce0030, /*   82 */
128'h84b68432e42efc06f04af426f8227139, /*   83 */
128'hcb5ff0ef083065a2c115cf7ff0ef893a, /*   84 */
128'h70e2978285a2615c862686ca6562e519, /*   85 */
128'hbfc5fda0051380826121790274a27442, /*   86 */
128'h84b68432e42efc06f04af426f8227139, /*   87 */
128'hc75ff0ef083065a2c115cb7ff0ef893a, /*   88 */
128'h70e2978285a2655c862686ca6562e519, /*   89 */
128'hbfc5fda0051380826121790274a27442, /*   90 */
128'hc7dff0ef84b2e42ef822fc06f4267139, /*   91 */
128'h701ce509c39ff0ef842a083065a2c105, /*   92 */
128'h8082612174a2744270e2978285a66562, /*   93 */
128'h2785c3190017f713419cbfcdfda00513, /*   94 */
128'hd71b8e5927a106220086571b419cc19c, /*   95 */
128'h0ff77713c19c0087d7138ed906a20086, /*   96 */
128'h122300d5112300c510238fd90087979b, /*   97 */
128'hf022f4067179419c80820005132300f5, /*   98 */
128'h419c00f510230457879b6785c19c27d1, /*   99 */
128'h0087979b0ff777130087d713c632842a, /*  100 */
128'hc4360509084c57fd460900f11a238fd9, /*  101 */
128'h0513016105934609783060ef00f11b23, /*  102 */
128'h00041323082c462147c1775060ef0044, /*  103 */
128'h00f404a347c5761060efec3e00840513, /*  104 */
128'h74b060ef00c4051300041523006c4611, /*  105 */
128'h0144069373f060ef01040513002c4611, /*  106 */
128'hfed79ce39f31ffe7d6030789470187a2, /*  107 */
128'h9fb94107d71b9fb9934117424107579b, /*  108 */
128'h80826145740270a200f41523fff7c793, /*  109 */
128'h97ba46a167856398338787930000b797, /*  110 */
128'hc7bb27850077e793fff6079b8007bc23, /*  111 */
128'h3823973e678500f547636805450102d7, /*  112 */
128'h010686bb0035169b0005b883808280c7, /*  113 */
128'he0221141bff105a125050116b02396ba, /*  114 */
128'hfa5ff0efe406450185aa86220005841b, /*  115 */
128'hec26f022717980820141640260a28522, /*  116 */
128'h68b060efe436f4064619051984b2842a, /*  117 */
128'h162347a167f060ef85b64619852266a2, /*  118 */
128'h614564e200e4859b70a27402852200f4, /*  119 */
128'h3a8130236785737dc5010113fadff06f, /*  120 */
128'h3931342338913c233a11342339213823, /*  121 */
128'h377134233761382337513c2339413023, /*  122 */
128'h3507879335a1382335913c2337813023, /*  123 */
128'hce042023d00007b7943e747d978a911a, /*  124 */
128'hd0040023f0040023e0040023ca040b23, /*  125 */
128'ha51785aa00e7ea63892a5800073797aa, /*  126 */
128'h00054703a00179f040eff52505130000, /*  127 */
128'h970a3507871374fd678526f711634789, /*  128 */
128'hcb848b13970a350787139abacd848a93, /*  129 */
128'h9c3a9b3a49818a368cb28baed0048c13, /*  130 */
128'hc7830015cd03013907b395ca0f098593, /*  131 */
128'h869b01a989bb058902a0071329890f07, /*  132 */
128'h24e78163471904f76b6326e78d630007, /*  133 */
128'hcc848513470d2ae78963470502f76263, /*  134 */
128'h40ef052505130000a51785b622e78963, /*  135 */
128'hfee794e3473d22e785634731b77d7170, /*  136 */
128'h953e866ae0048513978a350787936785, /*  137 */
128'h03600713b759e00d0023545060ef9d22, /*  138 */
128'h22e780630330071300f76e6322e78363, /*  139 */
128'haad94605cb648513fae798e303500713, /*  140 */
128'hf8e79ce30ff0071324e7856303800713, /*  141 */
128'h24e781630007859b747d471500614783, /*  142 */
128'h000ca7833ae79d63470938e781634719, /*  143 */
128'h05134985978a350a87936a8516079263, /*  144 */
128'h60ef013ca023953e461101090593ce44, /*  145 */
128'h01490593ce840513978a350a87934c90, /*  146 */
128'he28505130000a5174b3060ef953e4611, /*  147 */
128'h978a350a879364f040efde0254e25a52, /*  148 */
128'h439060ef854a55fd4619993ecf840913, /*  149 */
128'h879346f115231350079300f103a3478d, /*  150 */
128'h85a6460594becb740493c2a6978a350a, /*  151 */
128'h06a303200793461060efc0d246c10513, /*  152 */
128'h4a1195becf040593978a350a879346f1, /*  153 */
128'h079343d060ef4741072346f105134611, /*  154 */
128'hcf440593978a350a879346f109a30360, /*  155 */
128'h41b060ef47410a2347510513461195be, /*  156 */
128'h03a346f10ca347b1051385a6460557fd, /*  157 */
128'h061310200793401060ef47310d230001, /*  158 */
128'h079339b060efde3e37a1051345810f00, /*  159 */
128'h3961051385de4799464136f11d231010, /*  160 */
128'h13232637879377e13d3060ef36f10e23, /*  161 */
128'h350a879346f1142335378793679946f1, /*  162 */
128'h0440061304300693943ecec40413978a, /*  163 */
128'h85a2460156fdba1ff0ef3721051385a2, /*  164 */
128'h0e8885de86ca5672bd5ff0ef35e10513, /*  165 */
128'h3a0134033a813083911a6305cebff0ef, /*  166 */
128'h38013a03388139833901390339813483, /*  167 */
128'h36013c0336813b8337013b0337813a83, /*  168 */
128'h851380823b01011335013d0335813c83, /*  169 */
128'ha00d953e978a3507879367854611cd04, /*  170 */
128'h953e866af0048513978a350787936785, /*  171 */
128'h85564611b39df00d0023325060ef9d22, /*  172 */
128'h87936785bfdd855a4611bbb1317060ef, /*  173 */
128'h2fb060ef4611953ece048513978a3507, /*  174 */
128'h00f40123ce14478300f401a3ce044783, /*  175 */
128'h00f40023ce34478300f400a3ce244783, /*  176 */
128'h866ab759cc048513bb29cef42023401c, /*  177 */
128'h2783b311d00d00232c3060ef9d228562, /*  178 */
128'h0000a51700fa2023478512079a63000a, /*  179 */
128'h0e88010905934611451040efc3c50513, /*  180 */
128'hcb840513978a350487936485297060ef, /*  181 */
128'h3531470327f060ef014905934611953e, /*  182 */
128'h0000a517350145833511460335214683, /*  183 */
128'h00a1468335015783411040efc0c50513, /*  184 */
128'h35215783fcf71e230000b71700914603, /*  185 */
128'h0000b717c0c505130000a51700814583, /*  186 */
128'h01b147033dd040ef00b14703fcf71323, /*  187 */
128'h0000a517018145830191460301a14683, /*  188 */
128'h01214683013147033c1040efc0c50513, /*  189 */
128'hc10505130000a5170101458301114603, /*  190 */
128'h05130000a51755c2010157833a5040ef, /*  191 */
128'hb71701215783f6f713230000b717c1e5, /*  192 */
128'hf6bb02f5d63b03c00793f4f71e230000, /*  193 */
128'h02f5d5bbe107879b678502f6763b02f5, /*  194 */
128'h95bee0040593978a35048793365040ef, /*  195 */
128'h3504879334d040efbf8505130000a517, /*  196 */
128'hbf0505130000a51795be978af0040593, /*  197 */
128'h40efbfa505130000a517b501335040ef, /*  198 */
128'h20234785de0796e3000a2783bbcd3270, /*  199 */
128'ha51730b040efbee505130000a51700fa, /*  200 */
128'h3507879367852ff040efbf2505130000, /*  201 */
128'hbf8505130000a51795be978ad0040593, /*  202 */
128'hb35d2db040efbfe505130000a517bf45, /*  203 */
128'hf852fc4ee0cae4a6e8a2ec86711d737d, /*  204 */
128'h6a85c12505130000a517911a89aaf456, /*  205 */
128'h0493978a020a8793747d2b3040efca02, /*  206 */
128'hb79709b060ef852655fd461994beff84, /*  207 */
128'hc83e4a05fef40913439cd02787930000, /*  208 */
128'h993e978a020a879312f11d2313500793, /*  209 */
128'h07930bd060ef014107a31a68460585ca, /*  210 */
128'h020a879312f10f23479112f10ea30370, /*  211 */
128'h60ef13f10513461195beff040593978a, /*  212 */
128'h14f101a314510513460585ca57fd0990, /*  213 */
128'h0fc0079307f060ef000107a315410223, /*  214 */
128'h019060efca3e04a1051345810f000613, /*  215 */
128'h05134641479985ce04f1152310100793, /*  216 */
128'h2637879377e1051060ef04f106230661, /*  217 */
128'h879312f11c2335378793679912f11b23, /*  218 */
128'h06930421051385a2943e1451978a020a, /*  219 */
128'h02e1051385a2821ff0ef044006130430, /*  220 */
128'h85ce86a610084652855ff0ef460156fd, /*  221 */
128'h64a66446450160e6911a630596bff0ef, /*  222 */
128'ha51785aa808261257aa27a4279e26906, /*  223 */
128'h34238101011318f0406fb02505130000, /*  224 */
128'h34237d2138237c913c237e8130237e11, /*  225 */
128'h893689b2e04605a1051384aa71597d31, /*  226 */
128'h101867857ae060efd602e83eec3ae442, /*  227 */
128'h943e7fc404136762747d97ba81078793, /*  228 */
128'hf8aff0efd64e0521051385a2864a86ba, /*  229 */
128'hf0ef03e10513863e86c285a267c26822, /*  230 */
128'h8cfff0ef86c685a6180856326882fbaf, /*  231 */
128'h7d8134837e01340345017e8130836165, /*  232 */
128'h716d80827f0101137c8139837d013903, /*  233 */
128'h003547830045480300554883e222e606, /*  234 */
128'ha597842a000546030015468300254703, /*  235 */
128'h40efa52505130000a517a52585930000, /*  236 */
128'ha597860ac10d842adedff0ef85220c70, /*  237 */
128'h40efa5a505130000a517a32585930000, /*  238 */
128'h0000a51780826151641260b285220a70, /*  239 */
128'h089040efbe07ae230000b797a7450513, /*  240 */
128'hf85afc56e0d2e4ceeca6f0a27159b7cd, /*  241 */
128'h8a2ae46ee8caf486e86aec66f062f45e, /*  242 */
128'h718a8a930000aa974401ff05049389ae, /*  243 */
128'h0000ac1706000b93a48b0b130000ab17, /*  244 */
128'hfff58d1ba44c8c930000ac97a54c0c13, /*  245 */
128'h6a0669a6694664e6740670a603344163, /*  246 */
128'h61656da26d426ce27c027ba27b427ae2, /*  247 */
128'h009040ef855ae7a9c42900f477938082, /*  248 */
128'hfe05879b0007c583012487b34dc14901, /*  249 */
128'h09057ea040ef856602fbe2630ff7f793, /*  250 */
128'h7d8040ef574505130000a517ffb912e3, /*  251 */
128'hb7c57ca040ef8562a0317d2040ef8556, /*  252 */
128'h40ef9d2505130000a5170104c583dbe5, /*  253 */
128'h00f979134d81fffd4913028d1d637b60, /*  254 */
128'h855aff2dcce32d857a0040ef8556a029, /*  255 */
128'h00f45b630009079bff047913794040ef, /*  256 */
128'h0485240577c040ef518505130000a517, /*  257 */
128'hf793fe05879b0007c583012a07b3b781, /*  258 */
128'hb7e9090575c040ef856600fbe7630ff7, /*  259 */
128'he44ee84aec267179bfdd752040ef8562, /*  260 */
128'h86930000a697893289ae84b6f022f406, /*  261 */
128'h0000971794c686930000a697c50919e6, /*  262 */
128'h854a85a6944606130000a617dfc70713, /*  263 */
128'h85bb00955d6300098f63842a6d4040ef, /*  264 */
128'h40ef954a92c606130000a61786ce40a4, /*  265 */
128'hffd4841b00f44463ffe4879b9c296b60, /*  266 */
128'h26e060ef8fc585930000a59700890533, /*  267 */
128'h8082614569a2694264e2854a740270a2, /*  268 */
128'h0613002c7115f73ff06f4581862e86b2, /*  269 */
128'h0000a517002cfebff0efed8645050c80, /*  270 */
128'h8082612d450160ee6a0040ef8e450513, /*  271 */
128'h47b704a76963862e9ff787133b9ad7b7, /*  272 */
128'hf7633e70079304a7676323f78713000f, /*  273 */
128'h8e8707130000b7173e80079346890ca7, /*  274 */
128'he426e822ec0600074903e04a97361101, /*  275 */
128'ha51785aa690264a260e2644202091663, /*  276 */
128'h8793468163c0406f610588a505130000, /*  277 */
128'h02f57433bf7d240787934685b7d9a007, /*  278 */
128'h0287e66347293e800793c02102f555b3, /*  279 */
128'h0287746306300713c70502f4773347a9, /*  280 */
128'h0324341302e4743302f457b306400713, /*  281 */
128'h5433bfc102e45433a039943e00144413, /*  282 */
128'h40ef84b2834505130000a517f86102f4, /*  283 */
128'h40ef82a505130000a51785a2c8015d60, /*  284 */
128'ha517690264a285ca862660e264425c60, /*  285 */
128'h951785aa5ac0406f610581a505130000, /*  286 */
128'h481958d94781862eb78d7ea505130000, /*  287 */
128'h1782cd8500e555b303c6871b02f886bb, /*  288 */
128'he42697c211017f6808130000a8179381, /*  289 */
128'h60e26442e495e04ae822ec060007c483, /*  290 */
128'h61057ca505130000951785aa690264a2, /*  291 */
128'h0000951785aafb079de327855540406f, /*  292 */
128'hfff7c79300e797b357fdb7f57b450513, /*  293 */
128'h03b6869b02f5053347a9c10d44018d7d, /*  294 */
128'hf46300e45433942a47a500d414334405, /*  295 */
128'h89327625051300009517058514590087, /*  296 */
128'h758505130000951785a2c801504040ef, /*  297 */
128'h64a2690285a6864a60e264424f4040ef, /*  298 */
128'h71514da0406f61057605051300009517, /*  299 */
128'he96ae5cee9caf1a202c7073b8cbaed66, /*  300 */
128'he56ef162f55ef95afd56e1d2eda6f586, /*  301 */
128'h00e7f66384368d3289ae892a04000793, /*  302 */
128'hdcbb4cc1000c956302ccdcbb04000c93, /*  303 */
128'h0017849be03e020d1a13001d179b03ac, /*  304 */
128'h708b0b1300009b1703810a93020a5a13, /*  305 */
128'h5d8c0c1300008c17670b8b9300009b97, /*  306 */
128'h6a0e69ae694e64ee740e70ae4501e00d, /*  307 */
128'h616d6daa6d4a6cea7c0a7baa7b4a7aea, /*  308 */
128'h438040ef6c4505130000951785ca8082, /*  309 */
128'h470186ce000c8d9b008cf46300040d9b, /*  310 */
128'h971305b66c630007061b430948a14811, /*  311 */
128'h06bb0d9de66399ba034707339301020d, /*  312 */
128'h415705bb0006861b02e00813875603bd, /*  313 */
128'h05130000951785d6963e011c0ac5ed63, /*  314 */
128'h043b66a23dc040effa060c23e43667e5, /*  315 */
128'h557dd1350b8070ef99369281168241b4, /*  316 */
128'h260195d6002715934290030d1b63b795, /*  317 */
128'hec42f046f41a855a658292011602c190, /*  318 */
128'h96d27322674266a23a0040efe436e83a, /*  319 */
128'h15936290011d1863bf85686278820705, /*  320 */
128'h0006d603006d1c63bfc1e19095d60037, /*  321 */
128'hbf6500c590239241164295d600171593, /*  322 */
128'h00c580230ff6761300ea85b30006c603, /*  323 */
128'h6ae3270567220e4070efe43a855eb75d, /*  324 */
128'h053300074583bfdd4701bf1d3cfdfe97, /*  325 */
128'h0185959bc519097575130005450300bc, /*  326 */
128'hbf390705010700230005d4634185d59b, /*  327 */
128'h8082e21c00b7f4634501918187aa1582, /*  328 */
128'h89aa04000613fd4e7115bfd58f8d2505, /*  329 */
128'hf556f952e1cae5a6e9a2ed8600884581, /*  330 */
128'h577d67869982e16ae566e962ed5ef15a, /*  331 */
128'h55796318474707130000a7178ff98361, /*  332 */
128'h00009b174a8503800a13440106e79d63, /*  333 */
128'h80000c3758cb8b9300009b97554b0b13, /*  334 */
128'h07815783564d0d1300009d1708000cb7, /*  335 */
128'h06137786028a05bba091656600f46463, /*  336 */
128'h77c20957926347a299829dbd00280380, /*  337 */
128'h04090863792226e040ef855a85a2cfbd, /*  338 */
128'h0000951785a60397e863018487b37482, /*  339 */
128'h64ae644e60ee5575250040ef50450513, /*  340 */
128'h6caa6c4a6bea7b0a7aaa7a4a79ea690e, /*  341 */
128'h40ef856a86ca85a666428082612d6d0a, /*  342 */
128'h77a274c2998285260009061b45c22260, /*  343 */
128'h855e85ca993e86268c9d79020097ff63, /*  344 */
128'h24057fb050ef854a45818626204040ef, /*  345 */
128'ha7178082400005378082057e4505bfb1, /*  346 */
128'h869300756513157d631c57a707130000, /*  347 */
128'h057e450597aa20000537e30895360017, /*  348 */
128'h862a0ce507638207871367858082953e, /*  349 */
128'h4b050513000095178087871308a74463, /*  350 */
128'h000095178006079b04c7496306e60b63, /*  351 */
128'h0000951787f787936785c3ad48c50513, /*  352 */
128'h11417c07879b77fd04c7c96350c50513, /*  353 */
128'h05130000a5174fe58593000095979e3d, /*  354 */
128'h05130000a51760a213c040efe4064de5, /*  355 */
128'h05130000951781078713808201414ce5, /*  356 */
128'h0513000095178187879300e60a6345e5, /*  357 */
128'h00009517830787138082faf612e345e5, /*  358 */
128'h8287879300c74963fee609e347c50513, /*  359 */
128'h951783878713bfe94585051300009517, /*  360 */
128'h951784078793fce608e346a505130000, /*  361 */
128'h4205051300009517bf7546a505130000, /*  362 */
128'h84ae892af406e84aec26f02271798082, /*  363 */
128'h942a9041144201045513029044634401, /*  364 */
128'h1542fff54513740270a2952201045513, /*  365 */
128'h0068460985ca808261459141694264e2, /*  366 */
128'h00f107a334f9090900c147836f7050ef, /*  367 */
128'hbf55943e00e1578300f1072300d14783, /*  368 */
128'h8793f44ef84afc26e486e0a26785715d, /*  369 */
128'h0e636dd7879367a13cf50563842e8067, /*  370 */
128'h082884b205e944079a638005079b0af5, /*  371 */
128'ha517461985ca006409136a5050ef4611, /*  372 */
128'h079301744583691050ef3d2505130000, /*  373 */
128'h1cf5826347b108b7e76332f5896302e0, /*  374 */
128'h478502b7e3631af58363479104b7e563, /*  375 */
128'h83633aa5051300009517478910f58463, /*  376 */
128'ha41d7fb030ef546505130000951702f5, /*  377 */
128'h3b0505130000951747a118f582634799, /*  378 */
128'h2cf5826347f5a4317e1030effef591e3, /*  379 */
128'h0000951747d916f58a6347c500b7ed63, /*  380 */
128'h866302100793bf6dfef580e33cc50513, /*  381 */
128'h051300009517faf596e3029007932af5, /*  382 */
128'h04b7e2632cf5826306200793b7c93e65, /*  383 */
128'h02f0079300b7ef632af5826303300793, /*  384 */
128'h3e850513000095170320079328f58763, /*  385 */
128'h079328f5846305c00793b7bdf8f58ae3, /*  386 */
128'hbf91f6f58de33fe505130000951705e0, /*  387 */
128'h0670079300b7ef6328f5866308400793, /*  388 */
128'h410505130000951706c0079326f58b63, /*  389 */
128'h079326f5886308900793b73df4f58ae3, /*  390 */
128'h9517f0f59ce30880079326f589630ff0, /*  391 */
128'h0000a79701e45703b73d41a505130000, /*  392 */
128'h12f714632dc989930000a9972e47d783, /*  393 */
128'h10f71c632ce7d7830000a79702045703, /*  394 */
128'h0000a5974619531050ef852285ca4619, /*  395 */
128'h012301a45783521050ef854a29c58593, /*  396 */
128'h859b01c4578300f41f23020412230204, /*  397 */
128'h1d230009d78302f4102302240513fde4, /*  398 */
128'h0ea3db9ff0ef00f41e230029d78300f4, /*  399 */
128'h1223862601c1578300a10e23812100a1, /*  400 */
128'h00009517a06ddcbfe0ef450185a202f4, /*  401 */
128'hb55922a5051300009517bd4121c50513, /*  402 */
128'h470302444783bdb52385051300009517, /*  403 */
128'h178300f10e230254478300f10ea30264, /*  404 */
128'h00e10e2327810274470300e10ea301c1, /*  405 */
128'h0234470300e10ea301c1190302244703, /*  406 */
128'h04e79b6301c156830450071300e10e23, /*  407 */
128'h0000a597461947e21ad79e230000a797, /*  408 */
128'h0000a71719c505130000a51719458593, /*  409 */
128'ha79766a24762441050efe43618f72e23, /*  410 */
128'h450102a40593ff89061b172787930000, /*  411 */
128'h616179a2794274e2640660a6552060ef, /*  412 */
128'h0000a71747e204e69463043007138082, /*  413 */
128'hc799439c160787930000a79714f72e23, /*  414 */
128'h0000a697f7e9439c150787930000a797, /*  415 */
128'h0000a597140606130000a61714468693, /*  416 */
128'h0713b765d6dfe0ef02a4051314458593, /*  417 */
128'h30ef152505130000951702e798634d20, /*  418 */
128'h051300009517cdcff0ef852285a65670, /*  419 */
128'hcc6ff0ef02a4051385ca553030ef14e5, /*  420 */
128'h67c101e45703f6e787e35fe00713bf95, /*  421 */
128'h4611f4f70de302045703f6f701e317fd, /*  422 */
128'hb79936d050ef0868100585930000a597, /*  423 */
128'h051300009517b3351285051300009517, /*  424 */
128'h9517bb211445051300009517b30d12e5, /*  425 */
128'h1685051300009517b339152505130000, /*  426 */
128'h00009517b9ed16e5051300009517b311, /*  427 */
128'hb1dd19a5051300009517b9c518c50513, /*  428 */
128'h051300009517b9f11b05051300009517, /*  429 */
128'hd703b1e11e45051300009517b9c91d65, /*  430 */
128'h84930000a49707e7d7830000a7970265, /*  431 */
128'hd7830000a7970285d703ecf711e30764, /*  432 */
128'h89930205891320000793eaf719e30687, /*  433 */
128'h2bb050ef854a85ce461900f59a230165, /*  434 */
128'h2ab050ef854e026585930000a5974619, /*  435 */
128'h50ef00640513016585930000a5974619, /*  436 */
128'h01c4578328f050ef852285ca46192990, /*  437 */
128'h02f4142301e4578302f4132302a00613, /*  438 */
128'h00f41f230024d78300f41e230004d783, /*  439 */
128'h0000951785aab36900f4162360800793, /*  440 */
128'h300017b7bba54601401030ef16c50513, /*  441 */
128'h74132601608130239f0101138307b603, /*  442 */
128'h8406871b0387759366850034171b00f6, /*  443 */
128'h3c23630c8387b783972a300005379f2d, /*  444 */
128'h5f200813ffc5849b2581601134235e91, /*  445 */
128'h00c5963b101005938a1d08b8696335b9, /*  446 */
128'h87930000a797cfb527818ff1fff7c793, /*  447 */
128'h869b7007f7930084179bea254390f4e7, /*  448 */
128'h00d100a3872646d496aa068e9ebd8006, /*  449 */
128'h00d100230086d69b0106d69b0106969b, /*  450 */
128'h806686936685c6918005069b00015503, /*  451 */
128'h67139fad377d8005859b658502d51a63, /*  452 */
128'h868a83f502d7473b1782270546a10077, /*  453 */
128'h862602e6446397c285b6300008378f95, /*  454 */
128'h30838287b823300017b70405aa1ff0ef, /*  455 */
128'h610101135f8134838526600134036081, /*  456 */
128'hbc2306a126050008380300d788338082, /*  457 */
128'he42643c0e8220c2007b71101b7e1ff06, /*  458 */
128'h16938304b703300014b747812401ec06, /*  459 */
128'h0485051300009517e7990206c1630337, /*  460 */
128'h64a2644260e2c3c00c2007b72c5030ef, /*  461 */
128'hf0227179bfc14785eb9ff0ef80826105, /*  462 */
128'he78585930000a597461184ae8432ec26, /*  463 */
128'he30787930000a7970e3050eff4060068, /*  464 */
128'h88930000a89785a6862247b20007a803, /*  465 */
128'ha51704500693e1a757030000a717e168, /*  466 */
128'h740270a285228d4ff0efe22505130000, /*  467 */
128'h15428d5d05220085579b8082614564e2, /*  468 */
128'h8fd966c10185579b0185171b80829141, /*  469 */
128'h0085151b8fd98f750085571bf0068693, /*  470 */
128'h07b7715d808225018d5d8d7900ff0737, /*  471 */
128'h04b005134585460100740207879b0700, /*  472 */
128'hc63eec56f052f44efc26e0a2e486f84a, /*  473 */
128'h30eff825051300009517892a06d070ef, /*  474 */
128'hd8f70c230000a71757b90a091d631e70, /*  475 */
128'h0000a7175789d8f707a30000a7175785, /*  476 */
128'h5791d6f70ea30000a717578dd8f70323, /*  477 */
128'h6513893d003070efd6f70a230000a717, /*  478 */
128'h0000a5974611d6a781a30000a797fe05, /*  479 */
128'h0000a59746097e0050ef0048d5658593, /*  480 */
128'hf39ff0ef45127d0050ef0028d4458593, /*  481 */
128'h83210087179bf0060613010006374722, /*  482 */
128'h9101300016b78fd915020ff777138ff1, /*  483 */
128'h8006b78380f6b42393c180a6b02317c2, /*  484 */
128'h74e282f6b42347a1640660a68086b783, /*  485 */
128'h0000a497808261616ae27a0279a27942, /*  486 */
128'hec0a0a1300009a175ae14401ce448493, /*  487 */
128'h061b04852405855285a2028a863b4999, /*  488 */
128'h30effec48fa30ff6761300c956330286, /*  489 */
128'h8007b603300017b7bf91ff3410e30f70, /*  490 */
128'h8f4d91c115c20080073771398087b583, /*  491 */
128'he05ae456e852ec4ef04af426f822fc06, /*  492 */
128'h0b9030efe7c505130000951780e7b423, /*  493 */
128'hc6c7c7830000a797c73747030000a717, /*  494 */
128'hc5a6c6830000a697c65848030000a817, /*  495 */
128'hc485c5830000a597c51646030000a617, /*  496 */
128'h0000a41707d030efe505051300009517, /*  497 */
128'h89930000a997448100044783c3440413, /*  498 */
128'haa1700144783c2f703230000a717c0e9, /*  499 */
128'hc0f708a30000a7176a89c02a0a130000, /*  500 */
128'h0000a7173000193700262b3700244783, /*  501 */
128'hbef709a30000a71700344783bef70f23, /*  502 */
128'h00544783bef704230000a71700444783, /*  503 */
128'hba079a230000a797bcf70ea30000a717, /*  504 */
128'hba07a8230000a797ba07a4230000a797, /*  505 */
128'hb807ac230000a797ba07a2230000a797, /*  506 */
128'h0493ee5fe0ef8522e78d0009a783e4a9, /*  507 */
128'h37830207456303379713830937835a0b, /*  508 */
128'hbfc5bc3ff0effc075de3033797138309, /*  509 */
128'h849377d050ef4501dff154fd000a2783, /*  510 */
128'h4783b7d914fdb7e9ba9ff0efbfc1710a, /*  511 */
128'h4503002547838f5d07a2000547030015, /*  512 */
128'h57fd808225018d5d05628fd907c20035, /*  513 */
128'h058505050005c703808200f61363367d, /*  514 */
128'h808200f61363367d57fdb7f5fee50fa3, /*  515 */
128'hec06e8221101495cbfcd050500b50023, /*  516 */
128'h478101853903cfa500958413e04ae426, /*  517 */
128'h462d02e0031348a5481586ca02000513, /*  518 */
128'h07130107146300a70e6327850006c703, /*  519 */
128'h00e40023040500640023011795630e50, /*  520 */
128'h01c9051300b94783fcc79ee306850405, /*  521 */
128'h01994783c088f59ff0ef00f5842384ae, /*  522 */
128'h478300f492238fd90087979b01894703, /*  523 */
128'h00f493238fd90087979b016947030179, /*  524 */
128'h80826105690264a2644260e200040023, /*  525 */
128'h468303a0061302000593cf99873e611c, /*  526 */
128'h06630017869300c6986302d5fc630007, /*  527 */
128'h46050007c683b7dd0705a00d577d00d7, /*  528 */
128'h078900b666630ff6f593fd06869b577d, /*  529 */
128'h47030000a7178082853ae11c0006871b, /*  530 */
128'hc70d0007c703cb85611cc915bfd5a5e7, /*  531 */
128'he406114102e69063008557030067d683, /*  532 */
128'hc3914501001577933c4060ef0017c503, /*  533 */
128'h01b5c783808245258082014160a24525, /*  534 */
128'h0007079b8f5d0087979b468d01a5c703, /*  535 */
128'h0087979b0145c6830155c78300d51d63, /*  536 */
128'h71798082853e27818fd90107979b8fd5, /*  537 */
128'h0993e052e84af4065904e44eec26f022, /*  538 */
128'h60ef85ce8626468500154503842a0345, /*  539 */
128'h87bb000402234c58505ce13125013520, /*  540 */
128'h694264e2740270a2450100e7eb6340f4, /*  541 */
128'h74e34a0500344903808261456a0269a2, /*  542 */
128'h85ce86269cbd4685001445034c5cff2a, /*  543 */
128'h00454783b7f94505b7e5397d310060ef, /*  544 */
128'he8221101591c80824501f8dff06fc399, /*  545 */
128'h892e84aa02b787634401e04ae426ec06, /*  546 */
128'h46850014c503ec190005041bfddff0ef, /*  547 */
128'h4405c1192501298060ef03448593864a, /*  548 */
128'h690264a2644260e285220324a823597d, /*  549 */
128'h57fde04ae426ec06e822110180826105, /*  550 */
128'he52d2501fa3ff0ef842ad91c00050223, /*  551 */
128'h8fd90087979b45092324470323344783, /*  552 */
128'h1f63a55707134107d79b776d0107979b, /*  553 */
128'h05370005079bd59ff0ef06a4051302f7, /*  554 */
128'hf7b31465049300544537fff509130100, /*  555 */
128'hd33ff0ef0864051300978c6345010127, /*  556 */
128'h644260e200a035338d05012575332501, /*  557 */
128'hf84a715dbfcd450d80826105690264a2, /*  558 */
128'h3023e85aec56f052fc26e0a2e486f44e, /*  559 */
128'h4e6347addd9ff0ef8932852e89aa0005, /*  560 */
128'h97ba862787930000a797003517130205, /*  561 */
128'h000447830089b023c01547b184aa6380, /*  562 */
128'he38d001577931e2060ef00144503cb85, /*  563 */
128'h74e2640660a647a9c111891100090563, /*  564 */
128'h80826161853e6b426ae27a0279a27942, /*  565 */
128'h0f4060ef00a400a3000400230ff4f513, /*  566 */
128'hf569891100090463fb71478d00157713, /*  567 */
128'h848a04f51a634785ee1ff0ef85224581, /*  568 */
128'h4501ffc9478389a623a40a131fa40913, /*  569 */
128'h094100a9a0232501c5bff0ef854ac789, /*  570 */
128'h45090004aa8301048913ff2a14e30991, /*  571 */
128'h0491c10de9dff0ef852285d6000a8763, /*  572 */
128'h470db7bd00e519634785470dfe9915e3, /*  573 */
128'h4783bfb947b5c1194a81f6e504e34785, /*  574 */
128'h0107979b8fd90087979b03f447030404, /*  575 */
128'h04b44983fef711e3200007134107d79b, /*  576 */
128'h1a09866300f9e9b30089999b04a44783, /*  577 */
128'hfff9079b470501342e23044449032981, /*  578 */
128'h04144b03faf769e30ff7f793012401a3, /*  579 */
128'h00fb77b3fffb079bfa0b03e301640123, /*  580 */
128'h6a33008a1a1b0454478304644a03ffc9, /*  581 */
128'h04844503f3c100fa77930144142300fa, /*  582 */
128'h478314050e638d450085151b04744483, /*  583 */
128'hdfb18fd90087979b2501042447030434, /*  584 */
128'h00d7063b9f3d004a571b2781033906bb, /*  585 */
128'h84ae0364d5bb40c504bbf4c564e38732, /*  586 */
128'h0905165500b93933664119556905dd8d, /*  587 */
128'h015787bb248900ea873b490d00b67363, /*  588 */
128'h10e91263470dd05c03542023cc04d458, /*  589 */
128'h949bd408b17ff0ef06040513f00a15e3, /*  590 */
128'hee99e7e324810094d49b1ff4849b0024, /*  591 */
128'h478d00f402a3f8000793c45cc81c57fd, /*  592 */
128'h0087979b064447030654478308f91963, /*  593 */
128'h06f71b6347054107d79b0107979b8fd9, /*  594 */
128'h4783e13d2501ce5ff0ef8522001a859b, /*  595 */
128'h8fd90087979b000402a3232447032334, /*  596 */
128'h1263a55707134107d79b776d0107979b, /*  597 */
128'h2501416157b7a99ff0ef0344051304f7, /*  598 */
128'ha83ff0ef2184051302f5176325278793, /*  599 */
128'h051300f51c63272787932501614177b7, /*  600 */
128'ha63ff0ef22040513c808a6dff0ef21c4, /*  601 */
128'h93c117c227855e87d78300009797c448, /*  602 */
128'h0124002300f413235cf71d2300009717, /*  603 */
128'ha33ff0ef05840513b351478100042a23, /*  604 */
128'hb545a25ff0ef05440513b5b90005099b, /*  605 */
128'h949b00f915634789d41c9fb5e00a05e3, /*  606 */
128'h0017d79b8885029787bb478db7010014, /*  607 */
128'hf0ef842ae426ec06e8221101bdc59cbd, /*  608 */
128'h0cf71063478d00044703ed692501bfff, /*  609 */
128'h0613034404930af71b63478500544703, /*  610 */
128'h092305500793a01ff0ef852645812000, /*  611 */
128'h0a230520079322f409a3faa0079322f4, /*  612 */
128'h0da302f40b230610079302f40aa302f4, /*  613 */
128'h20e40d2302e40ba304100713481c20f4, /*  614 */
128'h20f40e230087571b0107571b0107971b, /*  615 */
128'h20f40fa30187d79b0107d71b20e40ea3, /*  616 */
128'h0107571b0107971b501020e40f23445c, /*  617 */
128'h22f4002307200693001445030087571b, /*  618 */
128'h0c230187d79b0107d71b260522e400a3, /*  619 */
128'hd81022f401a322e4012320d40ca320d4, /*  620 */
128'h00144503000402a363d050ef85a64685, /*  621 */
128'h60e200a035332501631050ef45814601, /*  622 */
128'h37f9ffe5869b4d1c8082610564a26442, /*  623 */
128'h9d2d02d585bb55480025458300f6f963, /*  624 */
128'h71794d180eb7f7634785808245018082, /*  625 */
128'h02e5f963892ae44eec26f022f406e84a, /*  626 */
128'h0e63468d06d70c63842e468900054703, /*  627 */
128'hd59b9cad515c0015d49b00f71e6308d7, /*  628 */
128'h70a257fdc9112501ac7ff0ef9dbd0094, /*  629 */
128'h278380826145853e69a2694264e27402, /*  630 */
128'h94ca1ff4f4930099d59b0014899b0249, /*  631 */
128'hf5792501a93ff0ef0344c483854a9dbd, /*  632 */
128'h0087979b880503494783994e1ff9f993, /*  633 */
128'hbf458fe9157d6505bf658391c0198fc5, /*  634 */
128'hfd592501a63ff0ef9dbd0085d59b515c, /*  635 */
128'h45030359478399221fe474130014141b, /*  636 */
128'h0075d59b515cb7598fc90087979b0349, /*  637 */
128'h75130024151bf9352501a39ff0ef9dbd, /*  638 */
128'h100007b7807ff0ef954a034505131fc5, /*  639 */
128'hf82271398082853e4785b76517fd2501, /*  640 */
128'h1523e456e852ec4ef426fc06f04a4540, /*  641 */
128'h744270e2450900f41c63892a478500b5, /*  642 */
128'h611c808261216aa26a4269e2790274a2, /*  643 */
128'h470d0007c683e02184aefee474e34f98, /*  644 */
128'hfce4f7e30087d703eb15579800e69463, /*  645 */
128'h37839d3d0044d79bd171008928235788, /*  646 */
128'h00a92a2394be03478793049688bd0009, /*  647 */
128'h843a0027c9838722b75d450100993c23, /*  648 */
128'h0134f66385a2000935034a8509925a7d, /*  649 */
128'h0005041be6fff0efbf752501e59ff0ef, /*  650 */
128'h76e34f9c00093783f68afbe301440c63, /*  651 */
128'h00a55583b78d4505bfc1413484bbf6f4, /*  652 */
128'h049bf33ff0ef842aec06e426e8221101, /*  653 */
128'h0005049b933ff0ef6008484ce4950005, /*  654 */
128'h6c1cf3cff0ef4581020006136c08ec99, /*  655 */
128'h60e200e782234705601c00e780235715, /*  656 */
128'hfc06e85271398082610564a285266442, /*  657 */
128'h16ba75634a05e456ec4ef04af426f822, /*  658 */
128'h4709000547830af5f063498984aa4d1c, /*  659 */
128'h94630ee78863470d0ae78f63842e8932, /*  660 */
128'h009a559b00ba0a3b515c0015da1b1547, /*  661 */
128'h8805060996630005099b8b9ff0ef9dbd, /*  662 */
128'h87b3cc191ffa7a130ff97793001a0a9b, /*  663 */
128'h179b00f7f71316c166850347c7830144, /*  664 */
128'h02fa0a239a260ff7f7938fd98ff50049, /*  665 */
128'h9dbd8526009ad59b50dc00f482234785, /*  666 */
128'h1ffafa9300099f630005099b86bff0ef, /*  667 */
128'h032a8a239aa60ff979130049591bc40d, /*  668 */
128'h790274a2854e744270e200f482234785, /*  669 */
128'hc783015487b3808261216aa26a4269e2, /*  670 */
128'h0127e9339bc100f979130089591b0347, /*  671 */
128'h099b811ff0ef9dbd0085d59b515cb7e9, /*  672 */
128'h94261fe474130014141bfc0992e30005, /*  673 */
128'h0089591b0109591b0109191b03240a23, /*  674 */
128'h0075d59b515cbf790144822303240aa3, /*  675 */
128'h141bf80996e30005099bfd8ff0ef9dbd, /*  676 */
128'hf0ef85569aa603440a931fc474130024, /*  677 */
128'h179b012569338d71f00006372501da0f, /*  678 */
128'h0087d79b03240a230107d79b94260109, /*  679 */
128'h00fa81230189591b0109579b00fa80a3, /*  680 */
128'hec4ef4267139bf3d4989b745012a81a3, /*  681 */
128'he19d89ae84aae456e852f04af822fc06, /*  682 */
128'h844a04f977634d1c04090a6300c52903, /*  683 */
128'h052a606304f4636324054c9c5afd4a05, /*  684 */
128'hf86347850005041bc43ff0efa8214401, /*  685 */
128'h744270e28522547d00f41d6357fd0887, /*  686 */
128'h4c9c808261216aa26a4269e2790274a2, /*  687 */
128'h85a24409bf554905b7d5faf47ee3894e, /*  688 */
128'h0863fd5507e3c9012501c05ff0ef8526, /*  689 */
128'h85a2167d10000637b76dfb2411e30545, /*  690 */
128'h489c02099063e9052501de9ff0ef8526, /*  691 */
128'h0054c783c89c37fdfae783e3577dc4c0, /*  692 */
128'h852685ce8622bf4900f482a30017e793, /*  693 */
128'h4405f6f50fe34785dd612501dbbff0ef, /*  694 */
128'h2905f822fc0600a55903f04a7139bfad, /*  695 */
128'heb9993c1e456e852ec4ef42603091793, /*  696 */
128'h6aa26a4269e2790274a2744270e24511, /*  697 */
128'h842a8a2e00f97993d7ed495c80826121, /*  698 */
128'h5783e18dc85c61082785480c00099d63, /*  699 */
128'h15230996601cfcf775e30009071b0085, /*  700 */
128'h4783bf5d4501ec1c97ce034787930124, /*  701 */
128'hfc0a9fe30157fab337fd00495a9b0025, /*  702 */
128'h45090097e46347850005049bb27ff0ef, /*  703 */
128'h4d1c6008b761450500f4946357fdbf49, /*  704 */
128'h049be81ff0ef480cf60a0ee306f4e063, /*  705 */
128'h8de357fdfcf48be34785d4bd451d0005, /*  706 */
128'h06136008f5792501dd8ff0ef6008fcf4, /*  707 */
128'h00043a03beeff0ef0345051345812000, /*  708 */
128'h60084a0502aa2823aa5ff0ef855285a6, /*  709 */
128'hd91c415787bb591c00faed6300254783, /*  710 */
128'h0223b7b9c848a83ff0ef85a6c8046008, /*  711 */
128'h5b1c2a856018f1412501d1cff0ef0145, /*  712 */
128'hf04afc06f426f8227139b7e9db1c2785, /*  713 */
128'h02f007130005c783e05ae456e852ec4e, /*  714 */
128'h0ce7906305c0071300e78663842e84aa, /*  715 */
128'h0ae7fc6347fd000447030004a6230405, /*  716 */
128'h47834b2102e0099305c00a9302f00a13, /*  717 */
128'h462d0204b9030d5780630d4782630004, /*  718 */
128'h926300044783b40ff0ef854a02000593, /*  719 */
128'h07930b37906300144783013900230d37, /*  720 */
128'h470d1b378e630024478300f900a302e0, /*  721 */
128'h458100f905a302000793943a09479763, /*  722 */
128'h608848cc100510632501adbff0ef8526, /*  723 */
128'hc7e5000747836c98e96d2501cdaff0ef, /*  724 */
128'h8d6300b78593709cef918ba100b74783, /*  725 */
128'h08e3fff7c683fff74603078507050cb7, /*  726 */
128'h4bdc611cbf75dfdff0ef85264581fed6, /*  727 */
128'hbc232501a85ff0ef85264581b791c55c, /*  728 */
128'h6aa26a4269e2790274a2744270e20004, /*  729 */
128'h8be3bf954709bf1d0405808261216b02, /*  730 */
128'h02400793943a12f6e06302000693f757, /*  731 */
128'h486502000313478145a147014681b7ad, /*  732 */
128'h9101020695130027e793a8dd0505a0d1, /*  733 */
128'h4503c6ed4711a06d268500e50023954a, /*  734 */
128'h00d90023469500d515630e5006930009, /*  735 */
128'h0037f6930ff7f7930027979b01659663, /*  736 */
128'h946346918bb10107671300b694634585, /*  737 */
128'h00e905a39432920116020087671300d7, /*  738 */
128'hc50500b7c783709c4511bf654701bdfd, /*  739 */
128'hcb890207f7930047f713f4e518e34711, /*  740 */
128'hbf154501e80703e30004bc230004a623, /*  741 */
128'h00b5c7836c8cfbf58b91b73d4515fb0d, /*  742 */
128'hc4c8af2ff0ef0007c503609cdbe58bc1, /*  743 */
128'h46a10ff7f7930027979b05659a63bdb9, /*  744 */
128'h47039722930117020017061b873245ad, /*  745 */
128'h0ae3f95704e3f94706e3f4e374e30007, /*  746 */
128'h4c634185551b0187151b02b6f263fd37, /*  747 */
128'h866300054883ece50513000085170005, /*  748 */
128'h7513fbf7051bbd6d4519f11710e30008, /*  749 */
128'h66e30ff57513f9f7051beea87ae30ff5, /*  750 */
128'h7179bdf90ff777130017e7933701eea8, /*  751 */
128'h451184aef406842ae44ee84aec26f022, /*  752 */
128'h6008a0b1c90de199484c49bd0e500913, /*  753 */
128'hc3210007c7036c1ce1292501afaff0ef, /*  754 */
128'h033780630327026303f7f79300b7c783, /*  755 */
128'h70a2450100979a630017b79317e18bfd, /*  756 */
128'h852245818082614569a2694264e27402, /*  757 */
128'h4511b7cd00042a23d9452501c13ff0ef, /*  758 */
128'hf0ef842ae426ec06e82245811101bfe5, /*  759 */
128'hf0ef6008484c0e500493e50d250188ff, /*  760 */
128'h00978d630007c7836c1ced092501a8cf, /*  761 */
128'h4791dd792501bcdff0ef85224585cb99, /*  762 */
128'h8082610564a2644260e2451d00f51363, /*  763 */
128'h049bfa9ff0ef842aec06e426e8221101, /*  764 */
128'h0005049ba42ff0ef6008484ce49d0005, /*  765 */
128'h700c84cff0ef4581020006136c08e085, /*  766 */
128'h00e782234705601c82aff0ef462d6c08, /*  767 */
128'hed6347858082610564a28526644260e2, /*  768 */
128'h694264e2740270a245098082450900b7, /*  769 */
128'hec26f02271794d1c808261456a0269a2, /*  770 */
128'hfcf5fde384ae842ae052e44ee84af406, /*  771 */
128'hf0ef852285a600f4fa634c1c59fd4a05, /*  772 */
128'h0ce3bf754501000914630005091bec8f, /*  773 */
128'h8afff0ef852285a6460103390763fb49, /*  774 */
128'h4783c81c278501378a63481cf15d2501, /*  775 */
128'hbf5d0009049b00f402a30017e7930054, /*  776 */
128'he432e82efc061028ec2a7139b7594505, /*  777 */
128'h8793000097970405426383eff0eff42e, /*  778 */
128'h0023c3196622631800a78733050eace7, /*  779 */
128'h4501e39897aa00070023c31967620007, /*  780 */
128'hf0ef0828080c460100f618634785cb11, /*  781 */
128'h7175bfe5452d8082612170e22501a0ef, /*  782 */
128'he8daecd6f0d2f4cefca6e122e506f8ca, /*  783 */
128'h84aa89b20005302314050d634925e42e, /*  784 */
128'h10630005091b9d6ff0ef1028002c8a79, /*  785 */
128'h2501b6dff0efe4be1028083c65a21409, /*  786 */
128'h01f9fa1301c9f7934519e011e1196406, /*  787 */
128'he75ff0ef102800f516634791c54dc3e1, /*  788 */
128'hcfcd008a77936406e949008a6a132501, /*  789 */
128'h0ca300f408a302100713046007937aa2, /*  790 */
128'h0b2300e40823000407a30004072300f4, /*  791 */
128'h0e23000405a300e40c2300040ba30004, /*  792 */
128'hc50300040fa300040f2300040ea30004, /*  793 */
128'h0da300040d234785fc9fe0ef85a2000a, /*  794 */
128'h82230005099b00040aa300040a230004, /*  795 */
128'hf0ef030aab03855685ce04098b6300fa, /*  796 */
128'h0135262385da39fd7522e9112501e3ff, /*  797 */
128'h00b44783a895892ac90d250183aff0ef, /*  798 */
128'ha0854921f60981e30049f993e3d98bc5, /*  799 */
128'h0029f993e72d0107f71300b44783f565, /*  800 */
128'h6a13c399008a7793e3ad8b8500098463, /*  801 */
128'h01448523f4800309a78385a279a2020a, /*  802 */
128'hc8c8f33fe0ef0009c503000485a3d09c, /*  803 */
128'ha623c8880069d783dbbfe0ef01c40513, /*  804 */
128'h60aa00f494230134b0230004ae230004, /*  805 */
128'h6b466ae67a0679a6794674e6854a640a, /*  806 */
128'hf8a27119b7d5491db7e5491180826149, /*  807 */
128'hfc5ee0daf0caf4a6fc86e4d6e8d2ecce, /*  808 */
128'h8a2e842a0006a023ec6ef06af466f862, /*  809 */
128'h000998630005099be91fe0ef8ab6e432, /*  810 */
128'h744670e60007899bc39d662200b44783, /*  811 */
128'h7be26b066aa66a4669e6790674a6854e, /*  812 */
128'h00a44783808261096de27d027ca27c42, /*  813 */
128'h40f907bb445c01042903160789638b85, /*  814 */
128'h0b1320000b930006091b00f67463893e, /*  815 */
128'h90631ff777934458fa090ce35c7d0304, /*  816 */
128'hfcb337fd0025478300975c9b60081207, /*  817 */
128'h47854848eb11020c99630ffcfc930197, /*  818 */
128'h4c0cb741498900f405a3478900a7ec63, /*  819 */
128'h05a3478501851763b7e52501bd6ff0ef, /*  820 */
128'h856e4c0c00043d83cc08b7a5498500f4, /*  821 */
128'h0099579b000c861bd5792501b98ff0ef, /*  822 */
128'h002dc683c4b58d3a0007849b00a6073b, /*  823 */
128'h86a6001dc503419684bb00f6f4639fb1, /*  824 */
128'h00a44783f94d250114a050ef85d2863a, /*  825 */
128'h0097fc6341a507bb4c48c3850407f793, /*  826 */
128'h955285da20000613910115020097951b, /*  827 */
128'h9a3e9381020497930094949bc5ffe0ef, /*  828 */
128'h9fa5000aa783c45c9fa54099093b445c, /*  829 */
128'h00a4478304e601634c50b70500faa023, /*  830 */
128'he43a85da4685001dc503c38d0407f793, /*  831 */
128'hf793672200a44783f1392501110050ef, /*  832 */
128'h0017c503863a4685601c00f40523fbf7, /*  833 */
128'h444c01a42e23f11525010bc050ef85da, /*  834 */
128'h0127f46340bb87bb1ff5f5930009049b, /*  835 */
128'he0ef855295a28626030585930007849b, /*  836 */
128'he4cee8caf0a27159b59d499dbf9dbd1f, /*  837 */
128'hec66f062f45ef85aeca6f486fc56e0d2, /*  838 */
128'h8ab689328a2e842a0006a023e46ee86a, /*  839 */
128'h00b44783000997630005099bcb5fe0ef, /*  840 */
128'h694664e6854e740670a60007899bc39d, /*  841 */
128'h6d426ce27c027ba27b427ae26a0669a6, /*  842 */
128'h18078f638b8900a44783808261656da2, /*  843 */
128'h0b1320000b9304f76c630127873b445c, /*  844 */
128'h93631ff777930409046344585c7d0304, /*  845 */
128'hfcb337fd0025478300975c9b60081407, /*  846 */
128'h4581485cef01040c9a630ffcfc930197, /*  847 */
128'h498900f405a3478902e798634705cb91, /*  848 */
128'h445cf3fd0005079bd86ff0ef4c0cb759, /*  849 */
128'h05230207e79300a4478312f76a634818, /*  850 */
128'h498500f405a3478501879763b79500f4, /*  851 */
128'hf79300a44783c85ce311cc1c4858bf99, /*  852 */
128'h85da0017c50346854c50601cc38d0407, /*  853 */
128'hfbf7f79300a44783f96925017b1040ef, /*  854 */
128'h97cff0ef856e4c0c00043d8300f40523, /*  855 */
128'h00a6863b0099579b000c869bd1592501, /*  856 */
128'h74639fb5002dc703c4b58d320007849b, /*  857 */
128'h40ef85d286a6001dc503419704bb00f7, /*  858 */
128'h0297f26341a587bb4c4cf15125017630, /*  859 */
128'h855a95d220000613918115820097959b, /*  860 */
128'h00f40523fbf7f79300a44783a4ffe0ef, /*  861 */
128'h093b445c9a3e9381020497930094949b, /*  862 */
128'h00faa0239fa5000aa783c45c9fa54099, /*  863 */
128'h00e7fa63445c481800c78e634c5cbdd1, /*  864 */
128'hfd0925016c7040ef85da4685001dc503, /*  865 */
128'h87bb1ff575130009049b444801a42e23, /*  866 */
128'h8626030505130007849b0127f46340ab, /*  867 */
128'h0407e79300a447839dbfe0ef952285d2, /*  868 */
128'h1141bd2d499db5f9c81cbf4100f40523, /*  869 */
128'h4783e1752501acffe0ef842ae406e022, /*  870 */
128'h601cc3950407f793cf690207f71300a4, /*  871 */
128'h685040ef030405930017c50346854c50, /*  872 */
128'h00f40523fbf7f79300a44783ed552501, /*  873 */
128'hc703741ce15d2501b77fe0ef6008500c, /*  874 */
128'h0107169b481800e785a30207671300b7, /*  875 */
128'h00d78ea300e78e230086d69b0106d69b, /*  876 */
128'h00e78fa300d78f230187571b0107569b, /*  877 */
128'h169b00e78d2300078ba300078b234858, /*  878 */
128'h0107171b00e78a2327010107571b0107, /*  879 */
128'h0106d69b00e78aa30087571b0107571b, /*  880 */
128'h046007130086d69b00e78c2302100713, /*  881 */
128'h000789a30007892300e78ca300d78da3, /*  882 */
128'h478500f40523fdf7f793600800a44783, /*  883 */
128'h4505ebbfe06f014160a2640200f50223, /*  884 */
128'h842ae406e022114180820141640260a2, /*  885 */
128'h25019cbfe0ef8522e9012501effff0ef, /*  886 */
128'h110180820141640260a200043023e119, /*  887 */
128'h879700054a6395bfe0efec060028e42a, /*  888 */
128'h452d8082610560e245013ea78d230000, /*  889 */
128'hf486f0a21028002c4601e42a7159bfe5, /*  890 */
128'h083c65a2ec190005041bb3bfe0efeca6, /*  891 */
128'h6586e41d0005041bcd2ff0efe4be1028, /*  892 */
128'h64e6740670a68522cbd8575277a2e991, /*  893 */
128'hc50374a2cb998bc100b5c78380826165, /*  894 */
128'hfcf41ee34791b7c5c8c897bfe0ef0004, /*  895 */
128'hf8cae122e506e42afca67175bfd94415, /*  896 */
128'h1828002c460184ae00050023f0d2f4ce, /*  897 */
128'h842677e2ecbe081ce5292501acdfe0ef, /*  898 */
128'h040a12634a16c2be02f009934bdc597d, /*  899 */
128'h071b3427470300008717e50567a24501, /*  900 */
128'h186300e780a303a0071300e780230307, /*  901 */
128'h00078023078d00e7812302f007130e94, /*  902 */
128'h808261497a0679a6794674e6640a60aa, /*  903 */
128'h18284581fd452501f89fe0ef18284585, /*  904 */
128'h0007c50365c677e2f5552501e6eff0ef, /*  905 */
128'h2501f63fe0ef18284581c2aa8cdfe0ef, /*  906 */
128'h77e2e1052501e48ff0ef18284581f949, /*  907 */
128'h01450e6325018a7fe0ef0007c50365c6, /*  908 */
128'h67a24711dd612501a9eff0ef18284581, /*  909 */
128'hf5cfe0ef1828100cb7594509f8e516e3, /*  910 */
128'hfc974703973610949301020797134781, /*  911 */
128'h05bbfff7871b04e462630037871beb05, /*  912 */
128'h96b2920166a20206961300e586bb40f4, /*  913 */
128'hb7319c3d01368023fff7c79301271a63, /*  914 */
128'h4603962a1088920102071613b7c12785, /*  915 */
128'h0789bddd4545b7e900c68023377dfc96, /*  916 */
128'h07850007470397369281020416936722, /*  917 */
128'hf8227139b709fe9465e3fee78fa32405, /*  918 */
128'h84ae842ae456e852ec4efc06f04af426, /*  919 */
128'h00b44783000917630005091bfb4fe0ef, /*  920 */
128'h790274a2854a744270e20007891bcf89, /*  921 */
128'h009777634818808261216aa26a4269e2, /*  922 */
128'h00042623445884bae3918b8900a44783, /*  923 */
128'h00a44783c81cfcf778e34818445ce4bd, /*  924 */
128'hf793445c4481bf7d00f405230207e793, /*  925 */
128'h099300a44783fc960ee34c50d3e51ff7, /*  926 */
128'hc50385ce4685601cc3850407f7930304, /*  927 */
128'hf79300a44783ed51250130f040ef0017, /*  928 */
128'h0017c50386264685601c00f40523fbf7, /*  929 */
128'h6008bf59cc44ed3525012bd040ef85ce, /*  930 */
128'hfff4869b377dc7290097999b00254783, /*  931 */
128'h413007bb02c6ed630337563b0336d6bb, /*  932 */
128'h4a855a7dd1c19c9dc45c27814c0c8ff9, /*  933 */
128'hd7b51ff4f793c45c9fa5445c0499ea63, /*  934 */
128'h9ca90094d49bcd112501c87fe0ef6008, /*  935 */
128'h47850005059b814ff0efe595484cbfb1, /*  936 */
128'h57fdbded490900f405a3478900f59763, /*  937 */
128'hc84cb5ed490500f405a3478500f59763, /*  938 */
128'he0efcb818b89600800a44783b765cc0c, /*  939 */
128'hc4bfe0efbf6984cee5990005059bfddf, /*  940 */
128'h4f9c601cfabafee3fd4588e30005059b, /*  941 */
128'h013787bb413484bbcc0c445cfaf5fae3, /*  942 */
128'h842ac52de42ef822fc067139b7bdc45c, /*  943 */
128'h67e2e1152501fe6fe0ef0828002c4601, /*  944 */
128'h250197cff0eff01c101ce01c852265a2, /*  945 */
128'h4515e7898bc100b5c783cd996c0ce529, /*  946 */
128'he30fe0ef0007c50367e2a02d00043023, /*  947 */
128'h00f414230067d7838522458167e2c448, /*  948 */
128'h70e2f971fcf50be347912501cbdfe0ef, /*  949 */
128'hfcf501e34791bfdd4525808261217442, /*  950 */
128'h2501dbafe0ef842ae406e0221141b7c1, /*  951 */
128'h717980820141640260a200043023e119, /*  952 */
128'hd98fe0ef892e842af406e84aec26f022, /*  953 */
128'he0ef8522458100091f63e8890005049b, /*  954 */
128'h64e269428526740270a20005049bc5ff, /*  955 */
128'hb32ff0ef852245810224302380826145, /*  956 */
128'h852285ca00042a2302f5136347912501, /*  957 */
128'h47912501f8bfe0ef85224581c68fe0ef, /*  958 */
128'hbf6584aad16dbf7d00042a2300f51663, /*  959 */
128'hf0a21028002c460184aee42aeca67159, /*  960 */
128'h083c65a2e00d0005041bedafe0eff486, /*  961 */
128'h6786e8010005041b872ff0efe4be1028, /*  962 */
128'h70a68522c10fe0ef102885a6c489cf81, /*  963 */
128'hf0a27159bfcd44198082616564e67406, /*  964 */
128'he0d28522002c46018b2ee42af85a8432, /*  965 */
128'hec66f062f45efc56e4cee8caeca6f486, /*  966 */
128'h2c836000000a1c6300050a1be7cfe0ef, /*  967 */
128'h00fb202302f76263ffec871b481c0184, /*  968 */
128'h7ae26a0669a6694664e68552740670a6, /*  969 */
128'h00044b83808261656ce27c027ba27b42, /*  970 */
128'h85ca4a8559fd4481490902fb9f634785, /*  971 */
128'h09550863093508632501a55fe0ef8522, /*  972 */
128'h00544783fef963e329054c1c2485e111, /*  973 */
128'hb74d009b202300f402a30017e793c804, /*  974 */
128'h1afd4c0944814981490110000ab7504c, /*  975 */
128'h2501d10fe0ef0015899b852200099e63, /*  976 */
128'h038b9163200009930344091385cee921, /*  977 */
128'he3918fd90087979b0009470300194783, /*  978 */
128'h854ab745fc0c94e33cfd39f909092485, /*  979 */
128'he1116582015575332501abcfe0efe02e, /*  980 */
128'hbfbd4a09b7494a05b7c539f109112485, /*  981 */
128'h842ae04aec06e426e8221101bfad8a2a, /*  982 */
128'hcb9100b44783e4910005049bbc4fe0ef, /*  983 */
128'h610564a269028526644260e20007849b, /*  984 */
128'h48144458cf390027f71300a447838082, /*  985 */
128'h600800f40523c8180207e793fed772e3, /*  986 */
128'hc53900042a232501a58ff0ef484cef01, /*  987 */
128'h091b94dfe0ef4c0cbf7d84aa00a405a3, /*  988 */
128'h06374c0cb7dd450502f9146357fd0005, /*  989 */
128'h85ca6008f9792501b37fe0ef167d1000, /*  990 */
128'h45094785b769449db7e12501a1cff0ef, /*  991 */
128'h00a44783fcf96ae34d1c6008fcf900e3, /*  992 */
128'h0017c50346854c50601cdba50407f793, /*  993 */
128'h00a44783f55d25016ec040ef03040593, /*  994 */
128'h4605e42a7175b7b100f40523fbf7f793, /*  995 */
128'hca0fe0eff8cafca6e122e5061008002c, /*  996 */
128'he3bfe0efe0be1008081c65a2e9052501, /*  997 */
128'h0207f79300b7c78345196786e1052501, /*  998 */
128'hcb810014f79300b5c483c59975e2eb89, /*  999 */
128'h790280826149794674e6640a60aa451d, /* 1000 */
128'h88c1cc0d0005041bad8fe0ef00094503, /* 1001 */
128'h100c02800613fc878de301492783c89d, /* 1002 */
128'h951fe0efcaa200a8458996cfe0ef00a8, /* 1003 */
128'hd94d2501836ff0ef00a84581f1612501, /* 1004 */
128'hf15525019f5fe0ef1008faf518e34791, /* 1005 */
128'h85a27502bf612501f20fe0ef7502e411, /* 1006 */
128'h4605e42a7171b769d575250191cff0ef, /* 1007 */
128'he152e54ee94aed26f506f1221028002c, /* 1008 */
128'hbd0fe0efe8eaece6f0e2f4def8dafcd6, /* 1009 */
128'he4be1028083c65a21c0414630005041b, /* 1010 */
128'h176347911c0409630005041bd67fe0ef, /* 1011 */
128'h9f630207f79300b7c783441967a61af4, /* 1012 */
128'h02630005091bb45fe0ef458175221807, /* 1013 */
128'h0b63440557fd16f90f63440947851809, /* 1014 */
128'h160414630005041ba98fe0ef752216f9, /* 1015 */
128'h0a13f6efe0ef85220109549b85ca7422, /* 1016 */
128'he0ef855200050c1b4581200006130344, /* 1017 */
128'h248188cfe0ef855202000593462d898f, /* 1018 */
128'h0fa30104949b0109199b0ff4fb1347c1, /* 1019 */
128'h0b930104d49b021007930109d99b02f4, /* 1020 */
128'hd99b046007930ff97a9304f4062302e0, /* 1021 */
128'h0a230200061304f406a30084d49b0089, /* 1022 */
128'h07a305540723040405a3040405230374, /* 1023 */
128'h0544051385d2049404a3056404230534, /* 1024 */
128'h00074603468d05740aa3772280efe0ef, /* 1025 */
128'h0723478100f69363571400d6166357d2, /* 1026 */
128'h06f4042327810107d79b0107969b06f4, /* 1027 */
128'h0086d69b0107d79b0106d69b0107979b, /* 1028 */
128'h00274b8306f404a306d407a30087d79b, /* 1029 */
128'h0005041bf59fe0ef1028040b99634c85, /* 1030 */
128'h0210071300e785a3752247416786e835, /* 1031 */
128'h00078ba300078b230460071300e78c23, /* 1032 */
128'h01678a2301378da301578d2300e78ca3, /* 1033 */
128'h041bd5afe0ef00f50223478500978aa3, /* 1034 */
128'h022303852823001c0d1b7522a82d0005, /* 1035 */
128'h20000613ec090005041b8dcfe0ef0195, /* 1036 */
128'h8c6a0ffbfb93f61fd0ef3bfd85524581, /* 1037 */
128'h70aa8522f25fe0ef85ca7522441db749, /* 1038 */
128'h7ba67b467ae66a0a69aa694a64ea740a, /* 1039 */
128'h7159b7c544218082614d6d466ce67c06, /* 1040 */
128'h10284605002c843284aee42aeca6f0a2, /* 1041 */
128'h1028083c65a2e13125019cafe0eff486, /* 1042 */
128'hc783451967a6e9152501b65fe0efe4be, /* 1043 */
128'h00b74783c30d6706e39d0207f79300b7, /* 1044 */
128'h008705a38c3d027474138c658cbd7522, /* 1045 */
128'h740670a62501c9efe0ef00f502234785, /* 1046 */
128'h002c4605e02ee42a71718082616564e6, /* 1047 */
128'h0005079b964fe0efed26f122f5060088, /* 1048 */
128'hf0be083cf4be008865a2678612079663, /* 1049 */
128'hc703778610079a630005079baf7fe0ef, /* 1050 */
128'h479165e61007126302077713479900b7, /* 1051 */
128'h0613e55fd0ef102805ad46550e058e63, /* 1052 */
128'hf05fd0ef850ae49fd0ef10a8008c0280, /* 1053 */
128'h079baadfe0ef10a865820c054d6347ad, /* 1054 */
128'hdc5fe0ef10a80ce793634711cbf90005, /* 1055 */
128'h851302a10593464d648aefc50005079b, /* 1056 */
128'h0207e793640602814783e0dfd0ef00d4, /* 1057 */
128'h8bc100b4c78300f40223478500f485a3, /* 1058 */
128'h85a60004450306f7086357d64736cbbd, /* 1059 */
128'h059bcaefe0ef85220005059bf2dfd0ef, /* 1060 */
128'h0005079bfc3fd0ef8522c5a547890005, /* 1061 */
128'h02f69d630557468302e007936706efb1, /* 1062 */
128'h27810107d79b06f707230107969b57d6, /* 1063 */
128'h0087d79b0107d79b0107979b06f70423, /* 1064 */
128'h07a3478506f704a30086d69b0106d69b, /* 1065 */
128'h0005079be24fe0ef008800f7022306d7, /* 1066 */
128'h740a70aa0005079bb50fe0ef6506e791, /* 1067 */
128'he8a2711dbfcd47a18082614d853e64ea, /* 1068 */
128'h810fe0efec861028002c4605842ee42a, /* 1069 */
128'h9abfe0efe4be1028083c65a2e9292501, /* 1070 */
128'h0207f79300b7c783451967a6e1292501, /* 1071 */
128'h00e78b23752200645703cb856786eb95, /* 1072 */
128'h00e78c230044570300e78ba30087571b, /* 1073 */
128'he0ef00f50223478500e78ca30087571b, /* 1074 */
128'he4a6711d80826125644660e62501ad6f, /* 1075 */
128'he8a208284601002c893284aee42ae0ca, /* 1076 */
128'h4581c4b9e0510005041bf9bfd0efec86, /* 1077 */
128'h08284585e5592501ca8fe0efd2020828, /* 1078 */
128'hd0ef8526462d75c2e93d2501b8ffe0ef, /* 1079 */
128'h000700230200061346ad00b48713ca1f, /* 1080 */
128'h97a6938117820007869bfff6879bce89, /* 1081 */
128'h656202090a63fec783e3177d0007c783, /* 1082 */
128'h470d6562e0150005041be69fd0ef510c, /* 1083 */
128'h0270079300e684630005468304300793, /* 1084 */
128'h852200a92023c29fd0ef953e03478793, /* 1085 */
128'h1563479180826125690664a6644660e6, /* 1086 */
128'he42a711db7d5842abf550004802300f5, /* 1087 */
128'h041bee3fd0efec86e8a21028002c4605, /* 1088 */
128'h02061793460100010c2366a2ec550005, /* 1089 */
128'hea2902000593eba10007c78397b69381, /* 1090 */
128'he8410005041bbd6fe0efda0210284581, /* 1091 */
128'h01814783e1792501abbfe0ef10284585, /* 1092 */
128'h07136786bc7fd0ef082c462dc3dd6506, /* 1093 */
128'h8ba300078b230460071300e78c230210, /* 1094 */
128'hbf45863eb74d2605a06100e78ca30007, /* 1095 */
128'h000747039736930102079713fff6079b, /* 1096 */
128'h07f00e9343658e2e4781082cfeb706e3, /* 1097 */
128'h91411542f9f7051b27850006c70348b1, /* 1098 */
128'h05130000751793411742370100a36c63, /* 1099 */
128'h8522441900eef863a82100070f1b8e65, /* 1100 */
128'h48030505bfcdf36d80826125644660e6, /* 1101 */
128'h00fe06b3b7cdffe81be3060805630005, /* 1102 */
128'h752200f500235795a885078500c68023, /* 1103 */
128'hb7c10005041b8fefe0ef00f502234785, /* 1104 */
128'he0ef1028dbd50181478302f51b634791, /* 1105 */
128'h4581020006136506f4450005041ba55f, /* 1106 */
128'h6786ae5fd0ef082c462d6506b07fd0ef, /* 1107 */
128'hf91780e3b751842abf1900e785a34721, /* 1108 */
128'h93811782f4c7e5e30585068500e58023, /* 1109 */
128'h4703f8d771e30007869b020006134729, /* 1110 */
128'h05052e83bf89eaf71de30e5007930181, /* 1111 */
128'hec22110105c528830585230305452e03, /* 1112 */
128'h87f2869a8646040502938f2ae44ae826, /* 1113 */
128'h8dfd00c6c5b345ef8f9300005f978876, /* 1114 */
128'h008fa403000f2583000fa38300b64733, /* 1115 */
128'h004f2703ff4fa3839db9007585bb0fc1, /* 1116 */
128'h0105e8330198581b0078159b0105883b, /* 1117 */
128'h8e6d00f6c6339f3100f805bb0077073b, /* 1118 */
128'h0146561b00c6171b9e39008f23838e35, /* 1119 */
128'hc6b300d383bb00c5873b008383bb8e59, /* 1120 */
128'hd39b007686bb8ebd00cf24038ef900b7, /* 1121 */
128'hffcfa4039fa100d3e6b30116969b00f6, /* 1122 */
128'h9fa1007777338f2d0007061b00d703bb, /* 1123 */
128'h0f418f5d0167171b00a7579b9f3d8f2d, /* 1124 */
128'hf45f17e300e387bb0003869b0005881b, /* 1125 */
128'h3d8f8f9300005f974a05859300005597, /* 1126 */
128'h00cf7f3300d7cf334a02829300005297, /* 1127 */
128'h0025c4030015c383000faf0301e6c733, /* 1128 */
128'h972a070a93aa038a0005c70300ef0f3b, /* 1129 */
128'h083b004fa70300ef0f3b942a040a4318, /* 1130 */
128'h0003a70301b8581b9e3900581f1b010f, /* 1131 */
128'h8e7501e7c6339f3100f80f3b010f6833, /* 1132 */
128'h0176561b0096139b008fa7039e398e3d, /* 1133 */
128'h05919f3500cf03bb00c3e63340189eb9, /* 1134 */
128'h0fc101e6c6b3fff5c4838efd007f46b3, /* 1135 */
128'h9fb900e6941b94aa048affcfa7039eb9, /* 1136 */
128'hc7339fb900d3843b8ec140980126d69b, /* 1137 */
128'h00c7579b9f3d0077473301e777330083, /* 1138 */
128'h069b0003861b000f081b8f5d0147171b, /* 1139 */
128'h0f1300005f17f25599e300e407bb0004, /* 1140 */
128'h010fc40332c38393000053978ffa3b6f, /* 1141 */
128'h00c2c4b3942a040a00d7c2b30003a703, /* 1142 */
128'h048a0043a4039f21011fc4839f254000, /* 1143 */
128'h171b012fc4830107083b40809e2194aa, /* 1144 */
128'h0083a4039e210107683301c8581b0048, /* 1145 */
128'h863b9ea194aa00e2c2b3048a00f8073b, /* 1146 */
128'h0156561b013fc90300b6129b408000c2, /* 1147 */
128'hffc3a4839c3500c702bb03c100c2e633, /* 1148 */
128'h941b992a9ea1090a0056c6b300e7c6b3, /* 1149 */
128'h843b8ec1000924830106d69b9fa50106, /* 1150 */
128'h9f3d8f219fa5005747330007081b00d2, /* 1151 */
128'h0002861b0f918f5d0177171b0097579b, /* 1152 */
128'h00005297f5f592e300e407bb0004069b, /* 1153 */
128'ha70300d745b38f5dfff647132a428293, /* 1154 */
128'h020f45839f2d022f4403021f43830002, /* 1155 */
128'h9f2d942a040a418c95aa058a93aa038a, /* 1156 */
128'ha5839e2d0068171b0107083b0042a583, /* 1157 */
128'h9db100f8073b0107683301a8581b0003, /* 1158 */
128'h139b0082a5839e2d8e3d8e59fff6c613, /* 1159 */
128'h03bb00c3e633400c9ead0166561b00a6, /* 1160 */
128'h0075e5b3fff7c593023f44839ead00c7, /* 1161 */
128'h00f5969b048a9db5ffc2a4038db902c1, /* 1162 */
128'h00b385bb40809fa18dd50115d59b94aa, /* 1163 */
128'h007747339fa18f4dfff747130007081b, /* 1164 */
128'h861b0f118f5d0157171b00b7579b9f3d, /* 1165 */
128'h6462f3ef9de300e587bb0005869b0003, /* 1166 */
128'h00c8863b00d306bb00fe07bb010e883b, /* 1167 */
128'h6105692264c2cd70cd34c97c05052823, /* 1168 */
128'he85af44ef84afc26e0a2715d653c8082, /* 1169 */
128'h84aa97b203f7f413ec56f052e486e45e, /* 1170 */
128'h07bb04000b9304000b13e53c893289ae, /* 1171 */
128'h0a1b00f974639381178200078a1b408b, /* 1172 */
128'h0084853385ce020ada93020a1a930009, /* 1173 */
128'h99d641590933481020ef0144043b8656, /* 1174 */
128'h60a6b7c997824401852660bc01741763, /* 1175 */
128'h6ba26b426ae27a0279a2794274e26406, /* 1176 */
128'h842a03f7f793f0227179653c80826161, /* 1177 */
128'hf800071300178513e84af406e44eec26, /* 1178 */
128'h40a9863b449d0400099300e7802397a2, /* 1179 */
128'h3c9020ef95224581920116020006091b, /* 1180 */
128'h97828522603cfc1c078e643c0124f563, /* 1181 */
128'h69a2694264e2740270a2fd24fde34501, /* 1182 */
128'h3423639cf4c787930000779780826145, /* 1183 */
128'hed3c639cf447879300007797e93c0405, /* 1184 */
128'h059311018082e13cb6c7879300000797, /* 1185 */
128'h769747013bf020efec06850a46410505, /* 1186 */
128'h454137a5859300006597162686930000, /* 1187 */
128'h0047d613070506890007c78300e107b3, /* 1188 */
128'h8f230007c78397ae000646038bbd962e, /* 1189 */
128'h0000751760e2fca71de3fef68fa3fec6, /* 1190 */
128'h0808842ae12271758082610512450513, /* 1191 */
128'hf0ef080885a26622f71ff0efe42ee506, /* 1192 */
128'h60aaf83ff0ef0808f01ff0ef0808e85f, /* 1193 */
128'h00d70d63711c46a1595880826149640a, /* 1194 */
128'h80824501cf980200071300d717634691, /* 1195 */
128'he426e82211018082556dbfe50007ac23, /* 1196 */
128'h569702f5026384ae842a200007b7ec06, /* 1197 */
128'h85930000659708800613052686930000, /* 1198 */
128'hfc2419b030ef2ee50513000065172de5, /* 1199 */
128'h6100e82211018082610564a2644260e2, /* 1200 */
128'h569702f4026384ae200007b7ec06e426, /* 1201 */
128'h85930000659702f0061302a686930000, /* 1202 */
128'he00415b030ef2ae505130000651729e5, /* 1203 */
128'h6100e82211018082610564a2644260e2, /* 1204 */
128'h569702f4026384ae200007b7ec06e426, /* 1205 */
128'h85930000659703600613ffa686930000, /* 1206 */
128'he40411b030ef26e505130000651725e5, /* 1207 */
128'h6104e42611018082610564a2644260e2, /* 1208 */
128'h769702f48263842e200007b7ec06e822, /* 1209 */
128'h85930000659703e00613ea2686930000, /* 1210 */
128'h14020db030ef22e505130000651721e5, /* 1211 */
128'h11018082610564a2644260e2e8809001, /* 1212 */
128'h8263842e200007b7ec06e8226104e426, /* 1213 */
128'h659704500613e56686930000769702f4, /* 1214 */
128'h30ef1ea50513000065171da585930000, /* 1215 */
128'h610564a2644260e2ec80900114020970, /* 1216 */
128'h200007b7ec06e4266100e82211018082, /* 1217 */
128'h0613f42686930000569702f4026384ae, /* 1218 */
128'h051300006517196585930000659704c0, /* 1219 */
128'h610564a2644260e2f004053030ef1a65, /* 1220 */
128'h200007b7ec06e4266100e82211018082, /* 1221 */
128'h0613f12686930000569702f4026384ae, /* 1222 */
128'h05130000651715658593000065970530, /* 1223 */
128'h610564a2644260e2f404013030ef1665, /* 1224 */
128'hf04af426f82200053983ec4e71398082, /* 1225 */
128'h02f984638436893284ae200007b7fc06, /* 1226 */
128'h0000659705a00613ed86869300005697, /* 1227 */
128'h30efe43a11c505130000651710c58593, /* 1228 */
128'h0029191b8b0589890014159b67227c60, /* 1229 */
128'h88a10125e5b30034949b8dd900497913, /* 1230 */
128'h69e2790274a202b9b8238dc5744270e2, /* 1231 */
128'h4605468147057100e022114180826121, /* 1232 */
128'hf0ef45818522f7dff0efe40645818522, /* 1233 */
128'hf67ff0ef45814605468547058522f35f, /* 1234 */
128'h01414501640260a2d97ff0ef45816008, /* 1235 */
128'h3c23460546814705e022e40611418082, /* 1236 */
128'h8522f39ff0ef842a4581040530230205, /* 1237 */
128'h46054685470545818522ef1ff0ef4581, /* 1238 */
128'hf06f0141458160a264026008f23ff0ef, /* 1239 */
128'h200007b7ec06e8226104e4261101d4df, /* 1240 */
128'h0613e02686930000569702f48263842e, /* 1241 */
128'h05130000651702658593000065970610, /* 1242 */
128'h644260e2fc80904114426e2030ef0365, /* 1243 */
128'hec06e8226104e42611018082610564a2, /* 1244 */
128'h86930000569702f48263842e200007b7, /* 1245 */
128'h6517fe2585930000659706800613dce6, /* 1246 */
128'h8c7d17fd678569e030efff2505130000, /* 1247 */
128'he82211018082610564a2644260e2e0a0, /* 1248 */
128'h02f4026384ae200007b7ec06e4266100, /* 1249 */
128'h0000659706f00613d986869300005697, /* 1250 */
128'h658030effac5051300006517f9c58593, /* 1251 */
128'he04a11018082610564a2644260e2e424, /* 1252 */
128'h842a200007b7ec06e426e82200053903, /* 1253 */
128'h0613d62686930000569702f9026384ae, /* 1254 */
128'h051300006517f5658593000065970760, /* 1255 */
128'h644260e2c84404993c23612030eff665, /* 1256 */
128'heca67100f0a2715980826105690264a2, /* 1257 */
128'hf062f45ef85afc56e0d2e4cef486e8ca, /* 1258 */
128'he03084b2892e0005d783020408a3ec66, /* 1259 */
128'h9c636ca020ef00c9051345814611d01c, /* 1260 */
128'h07b700043983bf5ff0ef458560080e04, /* 1261 */
128'h44810049278316f99a6304043a032000, /* 1262 */
128'h4c1c4485e391448d8b89c7090017f713, /* 1263 */
128'h8b85008a2783000a09638cdd03243c23, /* 1264 */
128'h45814605468147050144e49316078663, /* 1265 */
128'h2583be1ff0ef85224581d71ff0ef8522, /* 1266 */
128'hc4fff0efcdcc0c1300005c1785220089, /* 1267 */
128'hf0efe82a0a1300006a17852200095583, /* 1268 */
128'hf0ef85224581cbdff0ef852285a6c81f, /* 1269 */
128'hd27ff0ef85224581460546854705cf5f, /* 1270 */
128'h4585e93ff0ef852224058593000f45b7, /* 1271 */
128'h009899b785220d89b583cd1ff0ef8522, /* 1272 */
128'h6a9768198993eb7ff0ef25810015e593, /* 1273 */
128'h64e6740670a6efe9485ce42a8a930000, /* 1274 */
128'h6ce27c027ba27b427ae26a0669a66946, /* 1275 */
128'hdb7ff0efe024852244cc808261654501, /* 1276 */
128'hee079be38b85449cdf3ff0ef8522488c, /* 1277 */
128'h458163900107e683654100043883603c, /* 1278 */
128'h6e89f005051300ff0e37431147014781, /* 1279 */
128'h183b070500371f1b00064803ec0689e3, /* 1280 */
128'h0067036316fd060527810107e7b301e8, /* 1281 */
128'h981b010767330187971b0187d81bf2e5, /* 1282 */
128'h8fe9010767330087d79b01c878330087, /* 1283 */
128'h9746938183751782170200be873b8fd9, /* 1284 */
128'h869300005697b765470147812585e31c, /* 1285 */
128'h6517d62585930000659714900613b7e6, /* 1286 */
128'h00c4e493bd8541e030efd72505130000, /* 1287 */
128'h5597000b1d633b7d20000bb78b4ebd61, /* 1288 */
128'h00efd625051300006517b62585930000, /* 1289 */
128'h061386e20179096300043903b7116f60, /* 1290 */
128'h485c070934833de030ef855685d20f20, /* 1291 */
128'h37830209370312048e6324818cfd4c81, /* 1292 */
128'hcc5cf9200793c7817c1c00f76f630c89, /* 1293 */
128'hb27ff0ef85224581b6fff0ef85224581, /* 1294 */
128'hff397913852201442903c3950044f793, /* 1295 */
128'h0000651785cad47ff0ef85ca00896913, /* 1296 */
128'h2903c3950084f793680000efd0450513, /* 1297 */
128'hf0ef85ca00496913ff39791385220144, /* 1298 */
128'h658000efd04505130000651785cad1ff, /* 1299 */
128'h8c630384390300043c83cfb50014f793, /* 1300 */
128'h85d209c00613ace6869300005697017c, /* 1301 */
128'h3c2300492783cba97c1c332030ef8556, /* 1302 */
128'h018c871308e69f630037f693470d0204, /* 1303 */
128'hff87051363104591480d468100c90793, /* 1304 */
128'h8361ff87370301068763c3900086161b, /* 1305 */
128'h603cfeb690e30791872a2685c3988f51, /* 1306 */
128'hc85c9bf9485cc85c0027e793485ccbb5, /* 1307 */
128'h01748c63040439036004cc9d4c858889, /* 1308 */
128'h855685d20ca00613a686869300005697, /* 1309 */
128'h0089278300090963040430232b4030ef, /* 1310 */
128'h9bf54c85485cb4dff0ef8522ef8d8b85, /* 1311 */
128'h4505d80c8ee3c47ff0ef8522484cc85c, /* 1312 */
128'h2623000cb783dbd98b85bd95641020ef, /* 1313 */
128'h97a667a1bf41b1dff0ef8522b77100f9, /* 1314 */
128'h8913fa978de394be00093c8301096483, /* 1315 */
128'h39a020efe43e002c46218566639c0087, /* 1316 */
128'h0513717908b041635535b7dd87ca0ca1, /* 1317 */
128'h892e84b2e44ef406e84aec26f0220480, /* 1318 */
128'h0000551785a2cc1d5551842a1a4030ef, /* 1319 */
128'h6517862285aa89aa785010ef9d450513, /* 1320 */
128'h07b702098b634fe000efbd2505130000, /* 1321 */
128'hcb990024f793f40401242423e01c2000, /* 1322 */
128'h69a2694264e2740270a24501c45c4789, /* 1323 */
128'hb7e5c45c4785d4fd4501888580826145, /* 1324 */
128'h458146098082bff9557d18c030ef8522, /* 1325 */
128'h953e050e200007b7f73ff06f20000537, /* 1326 */
128'he4066380e0221141711c808225016108, /* 1327 */
128'h970686930000569702f40263200007b7, /* 1328 */
128'h00006517ab4585930000659734c00613, /* 1329 */
128'h557de3914505703c170030efac450513, /* 1330 */
128'h4501842ae822110180820141640260a2, /* 1331 */
128'h60e26622644285a24d3010efe42eec06, /* 1332 */
128'hf4062000051371797940006f61054685, /* 1333 */
128'h84aa0aa030efe052e44ee84aec26f022, /* 1334 */
128'h0001b5031b2030efb285051300006517, /* 1335 */
128'h206010ef842a491010ef450144b010ef, /* 1336 */
128'h3f8000ef638cb0e5051300006517681c, /* 1337 */
128'h3e8000efb0c505130000651706f44583, /* 1338 */
128'h15c20085d59bb165051300006517546c, /* 1339 */
128'h0000651706c44583583c3d2000ef91c1, /* 1340 */
128'h0187d61b0107d69b0087d71bb0c50513, /* 1341 */
128'h00ef26010ff6f6930ff7f7930ff77713, /* 1342 */
128'h398000efafc50513000065175c0c3a60, /* 1343 */
128'h00006597c789a865859300006597545c, /* 1344 */
128'h378000efaec5051300006517a7458593, /* 1345 */
128'h65977448102030efaf85051300006517, /* 1346 */
128'h584c19c42783dc3fb0ef0fa585930000, /* 1347 */
128'h061300006617e789a506061300006617, /* 1348 */
128'h852633a000efad65051300006517dae6, /* 1349 */
128'h0a1300006a174481ed5ff0ef84264581, /* 1350 */
128'hf79320000913ad69899300006997ad6a, /* 1351 */
128'h0004458330c000ef855285a6e78901f4, /* 1352 */
128'h04052fa000ef819100f5f6132485854e, /* 1353 */
128'h2e8000ef0845051300006517fd249fe3, /* 1354 */
128'h614545016a0269a2694264e2740270a2, /* 1355 */
128'h07b30003b6830083b7830103b7038082, /* 1356 */
128'h0017079300d7fe6393811782278540f7, /* 1357 */
128'h802345050103b78300a7002300f3b823, /* 1358 */
128'h0103b7830083b7038082450180820007, /* 1359 */
128'hfff706930003b7038f99920102059613, /* 1360 */
128'h86bb87aa9d9dfff7059b00c6f5638e9d, /* 1361 */
128'h852e0007002300b6e6630103b70340a7, /* 1362 */
128'h07850007c68300d3b823001706938082, /* 1363 */
128'h053be681000556634881bfe900d70023, /* 1364 */
128'hf81304100693c21906100693488540a0, /* 1365 */
128'h02b6733b0005061b385986ba4e250ff6, /* 1366 */
128'h02b6563b0305051b046e67630ff37513, /* 1367 */
128'h85bbfe718532fea68fa306850ff57513, /* 1368 */
128'h07930008876302f5e9630300051340e6, /* 1369 */
128'h0015559b40e6853b068500f6802302d0, /* 1370 */
128'h00b61b63fff5081b86ba258100068023, /* 1371 */
128'h2585fea68fa30685bf5d00a8053b8082, /* 1372 */
128'h0007c30397ba9381178240c807bbb7d9, /* 1373 */
128'h0685011780230066802326050006c883, /* 1374 */
128'heccef4a6f8a2597d011cf0ca7119b7f1, /* 1375 */
128'hf42afc3e843684b2e0dafc86e4d6e8d2, /* 1376 */
128'h03000a9306c00a1302500993f82af02e, /* 1377 */
128'hc52d8f1d0004c50377a2774202095913, /* 1378 */
128'h086304d7ff639381178276820017079b, /* 1379 */
128'hc503bfe1e7bff0ef0201039304850135, /* 1380 */
128'hc783035510634781048905450f630014, /* 1381 */
128'hf36346a50ff7f793fd07879bcb9d0004, /* 1382 */
128'h0f630640069304890014c503478100f6, /* 1383 */
128'h079304d50f630580069302a6eb6306d5, /* 1384 */
128'h790674a6744670e6f55d08f509630630, /* 1385 */
128'h808261090007051b6b066aa66a4669e6, /* 1386 */
128'h06e50e6307300713b74d048d0024c503, /* 1387 */
128'h00840b13f6e51ee30700071300a76c63, /* 1388 */
128'h02e5006307500713a00d460146850038, /* 1389 */
128'h00840b13fa850613f6e510e307800713, /* 1390 */
128'hf8b50693a81145c10016361346850038, /* 1391 */
128'h400845a946010016b693003800840b13, /* 1392 */
128'hf0ef0028020103930005059be37ff0ef, /* 1393 */
128'h00840b130201039300044503a809ddbf, /* 1394 */
128'h7433600000840b13b5fd845ad93ff0ef, /* 1395 */
128'h020103930005059b4db010ef85220124, /* 1396 */
128'hfc3ef83aec061034f436715db7f18522, /* 1397 */
128'h8082616160e2e8dff0efe436e4c6e0c2, /* 1398 */
128'hec06100005931014862ef436f032715d, /* 1399 */
128'h60e2e69ff0efe436e4c6e0c2fc3ef83a, /* 1400 */
128'h1234862afe36fa32f62e710d80826161, /* 1401 */
128'heac2e6bee2baea22ee06080810000593, /* 1402 */
128'h129020ef0808842ae3fff0efe436eec6, /* 1403 */
128'hb303679c691c80826135645260f28522, /* 1404 */
128'hee63479d808245018302000303630087, /* 1405 */
128'h83f94ca70713000047170205979304b7, /* 1406 */
128'h878297bae426e822ec061101439c97ba, /* 1407 */
128'h97930c5010ef7540f55c08c52483795c, /* 1408 */
128'he91c64a2644260e202f457b393810204, /* 1409 */
128'h35f1bfd9617cbfe97d5c808261054501, /* 1410 */
128'h557d8082557db7e9659c95aa058e05e1, /* 1411 */
128'h5e63ff5ff0ef842ae406e02211418082, /* 1412 */
128'h8522000307630207b303679c681c0005, /* 1413 */
128'h0141640260a245018302014160a26402, /* 1414 */
128'h4797150200a7eb6347ad8082557d8082, /* 1415 */
128'h551780826108953e8175452787930000, /* 1416 */
128'h0007b303679c691c80826d2505130000, /* 1417 */
128'h4785d23e47d502f1102347a1715d8302, /* 1418 */
128'h100c200007930030e83ee42e07851782, /* 1419 */
128'h8082616160a6fd3ff0efcc3ed402e486, /* 1420 */
128'h45018082450100e6fe63400407374d14, /* 1421 */
128'h24010113228134832301340323813083, /* 1422 */
128'h980101f1041322813823dc0101138082, /* 1423 */
128'hf0ef1a05348322113c232291342385a2, /* 1424 */
128'h02f71c630a0447830a04c703f579f95f, /* 1425 */
128'h0c04c70302f716630dd447830dd4c703, /* 1426 */
128'h0e0447830e04c70302f710630c044783, /* 1427 */
128'h10ef0d4485130d440593461100f71a63, /* 1428 */
128'h842af0227179b761fb600513d55156f0, /* 1429 */
128'h858a460185226ea020eff4063e800513, /* 1430 */
128'he509842af21ff0efc202c40200011023, /* 1431 */
128'h6145740270a285226cc020ef7d000513, /* 1432 */
128'hf406f022478500f11023478571798082, /* 1433 */
128'h008007b745386914c195842ac402c23e, /* 1434 */
128'h8f75600006b78ff58ff9f80787934ad4, /* 1435 */
128'h8522858a4601c43e8fd98f55400006b7, /* 1436 */
128'h6145740270a2c43c47b2e119ec9ff0ef, /* 1437 */
128'h5783c23e47d500f1102347b5711d8082, /* 1438 */
128'hfdf949370107979bf852fc4ee0ca07c5, /* 1439 */
128'h842e8aaaec86f456e4a6e8a26a056989, /* 1440 */
128'he00a0a13e0098993080909134495c43e, /* 1441 */
128'hf79345b2ed0de73ff0ef8556858a4601, /* 1442 */
128'h0125f7b3054793630135f7b3c7891005, /* 1443 */
128'h0513d4bff0ef52e5051300005517c78d, /* 1444 */
128'h7aa27a4279e2690664a6644660e6fba0, /* 1445 */
128'h0014079b347dfe04c6e334fd80826125, /* 1446 */
128'h4501b7555d8020ef3e80051300f05763, /* 1447 */
128'hd09ff0ef5045051300005517fc8049e3, /* 1448 */
128'h47c17139e7a919c52783bf7df9200513, /* 1449 */
128'hfc06f822858a460147d5c42e00f11023, /* 1450 */
128'h1b842783c11dde3ff0efc23e842af426, /* 1451 */
128'hdcdff0ef8522858a46014495cb918b89, /* 1452 */
128'h8082612174a2744270e2f8ed34fdc901, /* 1453 */
128'hec86e0cae4a6711d80824501bfd54501, /* 1454 */
128'h270347c906d7f66384b6892a4785e8a2, /* 1455 */
128'hd432cf3108c92783260102f1102302c9, /* 1456 */
128'hd23a854a100c47850030cc3ee42e4755, /* 1457 */
128'hf0634785e529842ad75ff0efc83eca26, /* 1458 */
128'h854a100c47f5460102f1102347b10497, /* 1459 */
128'h051300005517c11dd55ff0efd23ed402, /* 1460 */
128'h690664a6644660e68522c43ff0ef45e5, /* 1461 */
128'h841bb74d02f6063bbf6147c580826125, /* 1462 */
128'hf426f822fc067139b7c54401b7d50004, /* 1463 */
128'h8a2e4148842ace05e456e852ec4ef04a, /* 1464 */
128'h00b44583c11d892a482010ef8ab684b2, /* 1465 */
128'h014485b3681000054d638d3fa0ef8522, /* 1466 */
128'hbd9ff0ef414505130000551700b67a63, /* 1467 */
128'hf96decdff0ef854a08c92583a0894481, /* 1468 */
128'h844e0089f3630207e4030109378389a6, /* 1469 */
128'hfc851ae3f01ff0ef854a85d6865286a2, /* 1470 */
128'h9aa2028784339a22408989b308c96783, /* 1471 */
128'h69e274a279028526744270e2fc0999e3, /* 1472 */
128'h00f1102347997139808261216aa26a42, /* 1473 */
128'h161b8edd030007b70086969bc23e47f5, /* 1474 */
128'h440dc43684aafc06f426f8228ed10106, /* 1475 */
128'h3e800593e919c53ff0ef8526858a4601, /* 1476 */
128'h8082612174a2744270e2d91ff0ef8526, /* 1477 */
128'hbffc07b7db0101134d18bfcdfc79347d, /* 1478 */
128'h3c2324813023241134239fb923213823, /* 1479 */
128'h1ce7f56349013ffc0737233134232291, /* 1480 */
128'h892ac09ff0ef84aa85a2980101f10413, /* 1481 */
128'h20ef20000513e7991a04b7831e051863, /* 1482 */
128'h06131e0503631a04b5031aa4b0237660, /* 1483 */
128'h6b6347210c044783123010ef85a22000, /* 1484 */
128'h53b897ba078affe70713000047171cf7, /* 1485 */
128'h278300e7fd63cc981ff78793400407b7, /* 1486 */
128'h73630147d69307a68007071367050d44, /* 1487 */
128'h06f48f2309b449830a044783f8dc00d7, /* 1488 */
128'h4783c7890e244783e7810019f9938b85, /* 1489 */
128'h8b890a04478300098a6308f480a30b34, /* 1490 */
128'h07130e24478306f48fa309c44783c789, /* 1491 */
128'h05130a844783fcdc07c60c8486130914, /* 1492 */
128'h00074583fff74783e0fc07c6468109d4, /* 1493 */
128'h97aeffe745839fad0105959b0087979b, /* 1494 */
128'h02f585b30e04458300098c634685c391, /* 1495 */
128'h0621070de21c07ce02b787b30dd44783, /* 1496 */
128'h08d4470308e4478304098f63fca714e3, /* 1497 */
128'h08c447039fb90087171b0107979b4685, /* 1498 */
128'h87b30dd4478302f707330e04470397ba, /* 1499 */
128'h979b08a4470308b44783f8fc07ce02e7, /* 1500 */
128'h0087171b089447039fb90107171b0187, /* 1501 */
128'h07a6c319f4fc54d89fb9088447039fb9, /* 1502 */
128'h8bfd09c44783c7898b850a044783f4fc, /* 1503 */
128'hf0ef852645850af006134685ce81e391, /* 1504 */
128'h46830af447830af407a34785ed35e0bf, /* 1505 */
128'h54dc08f4aa2300a6979bc7b98b850e04, /* 1506 */
128'h4783f8dc07a60d44278300098663c799, /* 1507 */
128'h478308d4ac2302f686bb00a6969b0dd4, /* 1508 */
128'h854a240134032481308308f480230a74, /* 1509 */
128'h25010113228139832301390323813483, /* 1510 */
128'h8bfd8b7d0057d79b00a7d71b50fc8082, /* 1511 */
128'h892abf4d08f4aa2302f707bb27852705, /* 1512 */
128'hbf651a04b0235c8020efd1691a04b503, /* 1513 */
128'h22113c23dc010113bf455929bf555951, /* 1514 */
128'h88634789232130232291342322813823, /* 1515 */
128'h2381308354a9c585468102b7e16302f5, /* 1516 */
128'h01132281348322013903852623013403, /* 1517 */
128'h4685fef760e34705ffc5879b80822401, /* 1518 */
128'h84aad1fff0ef892a45850b900613842e, /* 1519 */
128'h01f10413f1e9258199f5ffe4059bf571, /* 1520 */
128'h0b944783e51998dff0ef854a85a29801, /* 1521 */
128'hec267179b74d84aab75ddf400493f7d5, /* 1522 */
128'h0ff5f99308154783f022f406e44ee84a, /* 1523 */
128'h45850b3006138edd892e9be10079f693, /* 1524 */
128'h00f51e63842a57b5c519cc7ff0ef84aa, /* 1525 */
128'h8526842a875ff0ef852685ca00091c63, /* 1526 */
128'h64e2740270a28522013505a315e010ef, /* 1527 */
128'h28113c23d60101138082614569a26942, /* 1528 */
128'h27313c23292130232891342328813823, /* 1529 */
128'h25713c23276130232751342327413823, /* 1530 */
128'h23b13c2325a130232591342325813823, /* 1531 */
128'hbff7879bbffc07b74d180ac7e9634789, /* 1532 */
128'h84ae8b32892abfe787933ffc07b79f3d, /* 1533 */
128'h07e9460300e7eb630185051300005517, /* 1534 */
128'hf0ef03a5051300005517e7b900167793, /* 1535 */
128'h29013403298130838522f8400413f96f, /* 1536 */
128'h27013a03278139832801390328813483, /* 1537 */
128'h25013c0325813b8326013b0326813a83, /* 1538 */
128'h2a01011323813d8324013d0324813c83, /* 1539 */
128'hdb450125051300005517098927038082, /* 1540 */
128'hac83e79102eaf7bb060a81630045aa83, /* 1541 */
128'h0185051300005517cb8902ecf7bb0005, /* 1542 */
128'h02eadabb02c92783bf415429f24ff0ef, /* 1543 */
128'h856200c488138c0a009c9c9be3994b85, /* 1544 */
128'h0017859b000828834e114e85478189d6, /* 1545 */
128'h010505130000551700030d6302e8f33b, /* 1546 */
128'hd33bb7f14b814a814c81b7c1ee4ff0ef, /* 1547 */
128'hc78397a6078e020880630065202302e8, /* 1548 */
128'hfb9300dbebb300be96bbcb898b850107, /* 1549 */
128'hfbc596e387ae05110821013309bb0ffb, /* 1550 */
128'h00e3ff250513000055178a09000b8963, /* 1551 */
128'hf0ef854a85d2fe0a7a1302f10a13f006, /* 1552 */
128'h09ea478309fa4603ee0519e3842af94f, /* 1553 */
128'h963e09da47839e3d0087979b0106161b, /* 1554 */
128'hf0effe2505130000551785ce01367a63, /* 1555 */
128'h0017f7130a7a46830084c783b5c1e56f, /* 1556 */
128'h0016e993c3990fe6f9938b89c71989b6, /* 1557 */
128'h4b189726070e0017059b461145054701, /* 1558 */
128'h00b517bb02080463001878130017581b, /* 1559 */
128'hd79b8b050189999b0187979b0027571b, /* 1560 */
128'h0ff9f99300f9e9b3c70d4189d99b4187, /* 1561 */
128'h8b850a6a478302d98263fcc592e3872e, /* 1562 */
128'hb591370020eff965051300005517ef89, /* 1563 */
128'h8b8509ba4783bfd100f9f9b3fff7c793, /* 1564 */
128'h547ddbaff0effc65051300005517cb89, /* 1565 */
128'h4685e3958b850afa4783e20b02e3b51d, /* 1566 */
128'h4785e569a21ff0ef854a45850af00613, /* 1567 */
128'h08f92a2300a7979b0e0a47830afa07a3, /* 1568 */
128'hf69301acd6bb08c00d934d0108800493, /* 1569 */
128'h2485ed499f1ff0ef854a458586260ff6, /* 1570 */
128'h08f00d134c81ffb492e32d210ff4f493, /* 1571 */
128'hf0ef854a458586260ff6f693019ad6bb, /* 1572 */
128'hffa492e32ca10ff4f4932485e9359cbf, /* 1573 */
128'h8656000c26834c818aa609b00d934d61, /* 1574 */
128'h99dff0ef854a0ff6f6930196d6bb4585, /* 1575 */
128'h248dffac90e30ffafa932ca12a85e139, /* 1576 */
128'h09c0061386defdb498e30c110ff4f493, /* 1577 */
128'hd4fb0de34785ed19975ff0ef854a4585, /* 1578 */
128'h458509b00613468501379b630a7a4783, /* 1579 */
128'h0a70061386cebb3d842a957ff0ef854a, /* 1580 */
128'h1141b32ddd79842a945ff0ef854a4585, /* 1581 */
128'h681c00055e63810ff0ef842ae406e022, /* 1582 */
128'h60a264028522000307630187b303679c, /* 1583 */
128'h713980820141640260a2450583020141, /* 1584 */
128'h00f5866384aa4791f04af822fc06f426, /* 1585 */
128'h00f110230370079304f5926355294785, /* 1586 */
128'h858a46010107979b4955842e07c4d783, /* 1587 */
128'h10234799ed19d52ff0efc43ec24a8526, /* 1588 */
128'h4601c43e478900f41f634791c24a00f1, /* 1589 */
128'h790274a2744270e2d34ff0ef8526858a, /* 1590 */
128'hee09b7cdc402fef414e3478580826121, /* 1591 */
128'h85be27814f1887ae00f5f3634f5c6918, /* 1592 */
128'hf06f02c50823dd0c0007059b00e7f463, /* 1593 */
128'h4b9c711910000737691c80828082c2cf, /* 1594 */
128'he4d6e8d2eccef0caf4a6fc86f8a2070d, /* 1595 */
128'hf0ef842ac17c8fd9f466f862fc5ee0da, /* 1596 */
128'h02042423eb8d6b9c679c681cc509f11f, /* 1597 */
128'hf8500493bacff0efdd85051300005517, /* 1598 */
128'h6aa66a4669e674a679068526744670e6, /* 1599 */
128'h4481541c808261097ca27c427be26b06, /* 1600 */
128'h082347851af42c23478df93ff0eff3e5, /* 1601 */
128'h7d000513ba2ff0ef852202042c2302f4, /* 1602 */
128'h84aa97826b9c679c8522681c421010ef, /* 1603 */
128'h22231a04282318042e2308842783f945, /* 1604 */
128'h45814601b72ff0ef8522d85c478508f4, /* 1605 */
128'hf14984aacf2ff0ef8522f1dff0ef8522, /* 1606 */
128'h00f1102347a1000505a345d000ef8522, /* 1607 */
128'he3991aa007138ff94bdc00ff8737681c, /* 1608 */
128'hc23ec43a8522858a460147d50aa00713, /* 1609 */
128'h15630aa0079300c14703e911bf8ff0ef, /* 1610 */
128'h037009933e900913cc1c800207b700f7, /* 1611 */
128'h80020c3700ff8bb74b0502900a934a55, /* 1612 */
128'hc252013110238522858a460140000cb7, /* 1613 */
128'h015110234c18681ce13dbb6ff0efc402, /* 1614 */
128'he7b301871563c43e0177f7b3c25a4bdc, /* 1615 */
128'hed1db8eff0ef8522858a4601c43e0197, /* 1616 */
128'h3e80051306090863397d0007ca6347b2, /* 1617 */
128'h00e68563800207374c14bf45331010ef, /* 1618 */
128'hd45c8b8541e7d79bc43ccc1880010737, /* 1619 */
128'hf9200793b55d18f40ca3478506041e23, /* 1620 */
128'hf0ef85224581c04ff0ef852202f51f63, /* 1621 */
128'h18f40c2347850007d663443ced09c34f, /* 1622 */
128'h00005517d965c1cff0ef85224585bfd1, /* 1623 */
128'h84aab595fa100493a10ff0efc5450513, /* 1624 */
128'he74eeb4aef26f706f3227161551cb585, /* 1625 */
128'he6eeeaeaeee6f2e2f6defadafed6e352, /* 1626 */
128'h199bc7831ff010ef45018baae3b54401, /* 1627 */
128'h10234789e7b5180b8ca3198bc783c7b1, /* 1628 */
128'hf0efc482c2be855e008c479d460104f1, /* 1629 */
128'hcf818b851b8ba783120500e3842aabaf, /* 1630 */
128'h03e3842aaa0ff0ef855e008c46014495, /* 1631 */
128'hf0ef855ea031020ba423f4fd34fd1005, /* 1632 */
128'h695a64fa741a70ba8522d55d842ad99f, /* 1633 */
128'h6d566cf67c167bb67b567af66a1a69ba, /* 1634 */
128'hc163180b8c23048ba7838082615d6db6, /* 1635 */
128'h149316d010ef4501b16ff0ef855e0407, /* 1636 */
128'hb36ff0ef855e45853e80091390810205, /* 1637 */
128'h10ef85260007cc63048ba783f155842a, /* 1638 */
128'hbfe91d7010ef0640051312a96ee31490, /* 1639 */
128'h41e7d79b048ba78300fbac23400007b7, /* 1640 */
128'h450dbf0506fb9e23478502fba6238b85, /* 1641 */
128'ha029400406370ea61ee345111aa60f63, /* 1642 */
128'h0036d61b00cbac234006061b40010637, /* 1643 */
128'h964e068a8a3d60e98993000039978a9d, /* 1644 */
128'h018ba88345051086a6830f86460396ce, /* 1645 */
128'hae231a0ba8238a0500c7d61b02d606bb, /* 1646 */
128'hd69b08dba22308dba42304cba823180b, /* 1647 */
128'h1408dc63090ba62300d5183b8abd0107, /* 1648 */
128'h0107979b14068e6302cba683090ba823, /* 1649 */
128'h938117828fd98ff50107571b003f06b7, /* 1650 */
128'hbc23030787b300e797b3070907854721, /* 1651 */
128'hbc230c0bb8230c0bb4230c0bb0230a0b, /* 1652 */
128'hd463200007930afbb8230e0bb0230c0b, /* 1653 */
128'hf46320000793090ba70308fba6230107, /* 1654 */
128'h8e63577d04cba783c21508fba82300e7, /* 1655 */
128'h1023855e008c46010107979b471100e7, /* 1656 */
128'h04f11023479d902ff0efc282c4be04e1, /* 1657 */
128'h855e008c0107979b4601495507cbd783, /* 1658 */
128'h4785e40516e3842a8e4ff0efc4bec2ca, /* 1659 */
128'hc9aff0ef855e08fb80a357fd08fbaa23, /* 1660 */
128'h00b545830f7000ef855ee2051ae3842a, /* 1661 */
128'h018ba703e0051fe3842affbfe0ef855e, /* 1662 */
128'h079304fba0232789100007b754075a63, /* 1663 */
128'h979b108c460107cbd78306f110230370, /* 1664 */
128'hd2caed05880ff0efd4bed2ca855e0107, /* 1665 */
128'h988102091a93033007930bf104934905, /* 1666 */
128'h108c08104b210a854a11d48206f11023, /* 1667 */
128'h3a7dc131850ff0efd05aec56e826855e, /* 1668 */
128'h0637a7a940020637bb45842afe0a16e3, /* 1669 */
128'ha82300b515bb89bd0165d59bbd994003, /* 1670 */
128'h569b8ff50027979b16f16685b54d08bb, /* 1671 */
128'hb5558b1d938100f7571b17828fd501e7, /* 1672 */
128'h161b0187179b0187569b00ff05374098, /* 1673 */
128'h06138fd167410087569b8e698fd50087, /* 1674 */
128'h559b40d804fbaa2327818fd58ef1f007, /* 1675 */
128'h571b8de90087159b8ecd0187169b0187, /* 1676 */
128'h0187d71b04ebac238f558f718ecd0087, /* 1677 */
128'h8001073720d702634689212700638b3d, /* 1678 */
128'h040ba7830007596302d7971300ebac23, /* 1679 */
128'h07b7018ba70304fba0238fd920000737, /* 1680 */
128'h639c03a78793000057971ef718638001, /* 1681 */
128'h020d1a13044ba783f0be4d05040ba903, /* 1682 */
128'h0ff1079300f979334284849300003497, /* 1683 */
128'h97bb478540980a05fe07fc1383f97913, /* 1684 */
128'h017d8b3716078563278100f977b300e7, /* 1685 */
128'h40dc0007ac8397d6109c840b0b1b4a81, /* 1686 */
128'h400007b7140781630197f7b300f977b3, /* 1687 */
128'h00fc88634591200007b700fc8d6345a1, /* 1688 */
128'hf0ef855e0015b59340bc85b3100005b7, /* 1689 */
128'h8d6347a1400007370e051c638daa971f, /* 1690 */
128'h100007b700ec886347912000073700ec, /* 1691 */
128'he0ef855e02fbaa23001cb79340fc8cb3, /* 1692 */
128'h4d850ce79163470d01a78663409cdfdf, /* 1693 */
128'h2d81810007b7d33e47d50af110234799, /* 1694 */
128'h110c040007930110d53e00fde7b317c1, /* 1695 */
128'h4783e941e91fe0efc93ee552e162855e, /* 1696 */
128'h9a631afba823409c09b794638bbd010c, /* 1697 */
128'h08bba2230017b79317ed088ba5831407, /* 1698 */
128'h0ff10793947ff0ef855e460118fbae23, /* 1699 */
128'h07cbd7830af1102303700793fe07fd93, /* 1700 */
128'hd33a8cee855e110c0107979b46014755, /* 1701 */
128'h102347b56702e915e35fe0efd53ee03a, /* 1702 */
128'h110c0110040007134791d502d33a0af1, /* 1703 */
128'he0dfe0efe03ac93ae552e16ee43e855e, /* 1704 */
128'h85b74785f3ed37fd670267a20e050c63, /* 1705 */
128'h4601180bae23096ba2231afba823017d, /* 1706 */
128'h94e347a10a918c9ff0ef855e84058593, /* 1707 */
128'he6f49fe32a4787930000379704a1eafa, /* 1708 */
128'hdf400413cbdfe0ef7305051300004517, /* 1709 */
128'h80020737b519a007071b80011737b61d, /* 1710 */
128'h80030737de075ee30307971300ebac23, /* 1711 */
128'h9881190201000ab70ff104934905bbc5, /* 1712 */
128'h10234799020a08633a7d09053ac54a15, /* 1713 */
128'h855e010c040007931030c33e47d508f1, /* 1714 */
128'hd0051ce3d61fe0efdc3ef84af426c556, /* 1715 */
128'hf006869366c144dcfbe18b8583a54cdc, /* 1716 */
128'h02e796938fd18ff50087d79b0087961b, /* 1717 */
128'h04fba02300876793da06d9e3040ba703, /* 1718 */
128'h837902079713eaf768e34581472db35d, /* 1719 */
128'h0537040d859366c1b54511872583974e, /* 1720 */
128'h0187d61b0d91000da783f006869300ff, /* 1721 */
128'h0087d79b8e690087961b8f510187971b, /* 1722 */
128'ha703fdb59ee3fefdae238fd98ff58f51, /* 1723 */
128'ha60300f6f8638bbd00c7579b46a5008c, /* 1724 */
128'h86930000369704d61c63800306b7018b, /* 1725 */
128'hae230087171b1487a78397b6078a0f66, /* 1726 */
128'h0186d61b8ff917fd67c100cca68308fb, /* 1727 */
128'hc305c38d03f7771327810126d71b8fd1, /* 1728 */
128'h57bb8a8d0106d69b02e6073b3e800613, /* 1729 */
128'ha7830adba2230afba02302d606bb02f7, /* 1730 */
128'h20000793c79919cba7831afbaa231b0b, /* 1731 */
128'h1523484000ef855e08fba82308fba623, /* 1732 */
128'hd6b7aaaab7b708cba703000506230005, /* 1733 */
128'h27818ef98ff9ccc68693aaa78793cccc, /* 1734 */
128'hf0f0f6b79fb500f037b3068600d036b3, /* 1735 */
128'h06b79fb5068a00d036b38ef90f068693, /* 1736 */
128'h9fb5068e00d036b38ef9f0068693ff01, /* 1737 */
128'h9fb9071200e037338f750207161376c1, /* 1738 */
128'hd70302c7d7b3ed1092010a8bb783d11c, /* 1739 */
128'h0000459784aa06fbc603074bd68307ab, /* 1740 */
128'ha95fe0effef536230245051356c58593, /* 1741 */
128'h0088579b06cbc603077bc883070ba803, /* 1742 */
128'h0ff878130ff7f7930188569b0108571b, /* 1743 */
128'h851354a585930000459726810ff77713, /* 1744 */
128'h859300004597074ba603a5ffe0ef04d4, /* 1745 */
128'h8abd0146561b0106569b062485135465, /* 1746 */
128'ha42347857e4010ef8526a3ffe0ef8a3d, /* 1747 */
128'h07b704fba0232785100007b7b8d102fb, /* 1748 */
128'h00004517e691ecf76ce31a0bb6834004, /* 1749 */
128'ha0230017079b70000737bb954c450513, /* 1750 */
128'hf6931adba42303f7f6930c46c78304fb, /* 1751 */
128'ha0230217071bc68900c7f693ce910027, /* 1752 */
128'h8b8504eba02301076713040ba70304eb, /* 1753 */
128'haa0304fba02300c7e793040ba783c799, /* 1754 */
128'h7a33855e4601088ba583044ba783040b, /* 1755 */
128'h4a85db4ff0effa6484930000349700fa, /* 1756 */
128'h8c9300003c974c2dfb8b0b1300003b17, /* 1757 */
128'hcbb5278100fa77b300fa97bb409cfeac, /* 1758 */
128'h10000db720000d37f989091300003917, /* 1759 */
128'h04f718630017b79317ed00494703409c, /* 1760 */
128'h4683c3a18ff900fa77b30009270340dc, /* 1761 */
128'he0ef855e0fb6f69345850b7006130089, /* 1762 */
128'he0ef855e45850b7006134681c131debf, /* 1763 */
128'ha223180bae231a0ba823088ba783ddbf, /* 1764 */
128'h11e30931973fe0ef855e035baa2308fb, /* 1765 */
128'h3985051300004517f7649fe304a1fb99, /* 1766 */
128'h4721400006b700092783bb6d925fe0ef, /* 1767 */
128'hb71341b787b301a78663471100d78963, /* 1768 */
128'h855e408c933fe0ef855e02ebaa230017, /* 1769 */
128'he79d0046f79300892683f941808ff0ef, /* 1770 */
128'hb79317ed088ba583ef8d1afba823409c, /* 1771 */
128'hf0ef855e460118fbae2308bba2230017, /* 1772 */
128'h0ff6f693bb91fd319fdfe0ef855ecb0f, /* 1773 */
128'hb7c9f521d31fe0ef855e45850b700613, /* 1774 */
128'h2583974e837902079713fcfc65e34581, /* 1775 */
128'h6da000ef06cb851300ec4641bf6d1187, /* 1776 */
128'h979b008c460107cbd78304f11023478d, /* 1777 */
128'h842a96ffe0efc2be47d5855ec4be0107, /* 1778 */
128'h04e157830007d663018ba783ec051b63, /* 1779 */
128'hd783c2be479d04f1102347a506fb9e23, /* 1780 */
128'he0efc4be855e0107979b008c460107cb, /* 1781 */
128'h45e6475647c646b6ea051163842a93bf, /* 1782 */
128'h06eba22306fba02304dbae23018ba503, /* 1783 */
128'h01a6d61bf2c51a634000063706bba423, /* 1784 */
128'h09634505f0c543638ca602e345098a3d, /* 1785 */
128'h0413f0eff06f2006061b40010637f0a6, /* 1786 */
128'h8082557d80824501c56ce54ff06ffa10, /* 1787 */
128'h879300005797808218b50d238082557d, /* 1788 */
128'h842ae406e02247851141ef9d439cbea7, /* 1789 */
128'he0ef852212a000efbcf72a2300005717, /* 1790 */
128'h02c00513fc5ff0ef852200055563aeef, /* 1791 */
128'h01414501640260a20dc000ef13e000ef, /* 1792 */
128'h631cba27071300005717808245018082, /* 1793 */
128'h05130000451785aa114102e790636394, /* 1794 */
128'h0141853e478160a2f60fe0efe4063465, /* 1795 */
128'h853ebfd187b600a604630fc7a6038082, /* 1796 */
128'hc105fbdff0efe42eec06110141488082, /* 1797 */
128'h07930815470302b7006365a210354703, /* 1798 */
128'h5535eb3fe06f610560e200f70c630ff0, /* 1799 */
128'hbfcdf8400513bfe545018082610560e2, /* 1800 */
128'hcd09f7dff0ef84aee822ec06e4261101, /* 1801 */
128'h60e2e0800f840413e501cf0ff0ef842a, /* 1802 */
128'h00005797bfd555358082610564a26442, /* 1803 */
128'h05138082c3980015071b438898c78793, /* 1804 */
128'h80824388974787930000579780820f85, /* 1805 */
128'he4266380e822ad678793000057971101, /* 1806 */
128'h610564a2644260e20094176384beec06, /* 1807 */
128'h6000a9cff0ef8522c78119a447838082, /* 1808 */
128'h5797e79ce39caa67879300005797b7d5, /* 1809 */
128'h879300005797e50880829207a5230000, /* 1810 */
128'h711d8082e308e518e11ce7886798a8e7, /* 1811 */
128'hfc4e6080e8a2a764849300005497e4a6, /* 1812 */
128'hec86e06ae466e862ec5ef05af456f852, /* 1813 */
128'h00004a97234a0a1300004a1789aae0ca, /* 1814 */
128'h00004b9722cb0b1300004b17224a8a93, /* 1815 */
128'h810c8c9300004c9700050c1b22cb8b93, /* 1816 */
128'h79e2690664a660e66446029415634d29, /* 1817 */
128'h45176d026ca26c426be27b027aa27a42, /* 1818 */
128'h4901541cddcfe06f612537a505130000, /* 1819 */
128'h2603681c89560007c36389524c1cc791, /* 1820 */
128'h85ca00090663dbefe0ef638c855a0fc4, /* 1821 */
128'h856685e200978e63601cdb2fe0ef855e, /* 1822 */
128'h798505130000351701a98863da4fe0ef, /* 1823 */
128'he426ec06e8221101b771600032a010ef, /* 1824 */
128'hcbbd4d5ccfad44014d1cc1414401e04a, /* 1825 */
128'h84aa892ec7ad639cc7bd651ccbad511c, /* 1826 */
128'h57fdcd21842a200010ef45051c000593, /* 1827 */
128'he90410f502a347850ef52c234799c57c, /* 1828 */
128'hfffff797e65ff0ef0405282303253023, /* 1829 */
128'h2be787930000179716f43c2391c78793, /* 1830 */
128'h18f434232ae787930000179718f43023, /* 1831 */
128'h10f400230247c78385220ea42e23681c, /* 1832 */
128'h6105690264a2644260e28522e99ff0ef, /* 1833 */
128'h611c6b268693000046971bc0106f8082, /* 1834 */
128'he11897360017671302d786b365186294, /* 1835 */
128'h07b300f7553b93ed836d8f3d0127d713, /* 1836 */
128'h00005517808225018d5d00f717bb40f0, /* 1837 */
128'hf0efe022e4061141fc3ff06f8ec50513, /* 1838 */
128'h60a28d410105151bfe9ff0ef842afeff, /* 1839 */
128'hf0efe022e40611418082014125016402, /* 1840 */
128'h15029001fd1ff0ef14020005041bfdbf, /* 1841 */
128'hc703058587aa80820141640260a28d41, /* 1842 */
128'h87aa962a8082fb75fee78fa30785fff5, /* 1843 */
128'hfee78fa30785fff5c703058500c78963, /* 1844 */
128'heb09001786930007c70387aa8082fb65, /* 1845 */
128'h8082fb75fee78fa30785fff5c7030585, /* 1846 */
128'h0007c70387b68082e21987aab7d587b6, /* 1847 */
128'h8713fff5c6830585963efb7d00178693, /* 1848 */
128'h80a300c715638082e291fed70fa30017, /* 1849 */
128'hc783000547030585b7cd87ba80820007, /* 1850 */
128'he3994187d79b0187979b40f707bbfff5, /* 1851 */
128'h478100c59463962e8082853ef37d0505, /* 1852 */
128'h40f707bbfff5c783000547030585a839, /* 1853 */
128'h853eff790505e3994187d79b0187979b, /* 1854 */
128'h808200b79363000547830ff5f5938082, /* 1855 */
128'h47830ff5f59380824501bfcd0505c399, /* 1856 */
128'h87aabfcd0505dffd808200b793630005, /* 1857 */
128'hbfcd0785808240a78533e7010007c703, /* 1858 */
128'h65a2fe5ff0efec06842ae42ee8221101, /* 1859 */
128'h157d00b78663000547830ff5f5939522, /* 1860 */
128'h95aa80826105644260e24501fe857be3, /* 1861 */
128'h40a78533e7010007c70300b7856387aa, /* 1862 */
128'h85330007c68387aa862ab7fd07858082, /* 1863 */
128'h000748030705fed80fe38082ea9940c7, /* 1864 */
128'h87aa86aabfcd872eb7d50785fe081be3, /* 1865 */
128'h00c80a638082ea1140d785330007c603, /* 1866 */
128'hbfd5872e8082fe081be3000748030705, /* 1867 */
128'h8fe380824501eb1900054703bff90785, /* 1868 */
128'h87aeb7e50505fafd0007c6830785fee6, /* 1869 */
128'he519842a84aeec06e426e8221101bfd5, /* 1870 */
128'h85a68522cc1163806e87879300004797, /* 1871 */
128'h00004797ef8100044783942af9dff0ef, /* 1872 */
128'h610564a2644260e2852244016c07b623, /* 1873 */
128'h00054783c519f9fff0ef852285a68082, /* 1874 */
128'h6aa7b02300004797050500050023c781, /* 1875 */
128'h842ac891e822ec066104e4261101bfd9, /* 1876 */
128'he008050500050023c501f73ff0ef8526, /* 1877 */
128'h4783c11d8082610564a28526644260e2, /* 1878 */
128'h0017c703ce810007c68387aacf990005, /* 1879 */
128'hb7e5078900d780a300e780238082e311, /* 1880 */
128'h9063963e87aacb9d0075779380824501, /* 1881 */
128'h08b3872aff6d377d8fd507a2808204c7, /* 1882 */
128'h003657930106ef6340e88833469d00c5, /* 1883 */
128'h4725bfc1963a97aa078e02e787335761, /* 1884 */
128'h0785bfe1fef73c230721bfd10ff5f693, /* 1885 */
128'h8b9d00a5e7b300b50a63bf6dfeb78fa3, /* 1886 */
128'h38030721808202c79e63963e87aacb9d, /* 1887 */
128'hff06e8e340f88833ff07bc2307a1ff87, /* 1888 */
128'h963e95ba070e02f707b357e100365713, /* 1889 */
128'h469d00c508b387aa872ebfc100e507b3, /* 1890 */
128'hbf65fee78fa30785fff5c7030585bfe1, /* 1891 */
128'he84af406e432ec26852e842af0227179, /* 1892 */
128'h6582892ace1184aa6622dcdff0efe02e, /* 1893 */
128'hf0ef944a864a8522fff6091300c56463, /* 1894 */
128'h64e269428526740270a200040023f79f, /* 1895 */
128'h00a5e963842ae406e022114180826145, /* 1896 */
128'h95b280820141640260a28522f57ff0ef, /* 1897 */
128'h15fdd7e500e587b340b6073300c506b3, /* 1898 */
128'h1563962ab7fd00f6802316fd0005c783, /* 1899 */
128'h0005c703000547838082853e478100c5, /* 1900 */
128'h00c51363962ab7dd05850505fbed9f99, /* 1901 */
128'h7179bfc50505feb78de3000547838082, /* 1902 */
128'h89aee84af406e44eec26852e842af022, /* 1903 */
128'hd13ff0ef8522c8890005049bd1fff0ef, /* 1904 */
128'h740270a28522440100995b630005091b, /* 1905 */
128'h852285ce86268082614569a2694264e2, /* 1906 */
128'hf593962abfe90405d175f8bff0ef397d, /* 1907 */
128'h0793000547038082450100c514630ff5, /* 1908 */
128'h0ff5f59347c1b7ed853efeb70be30015, /* 1909 */
128'h8082853e4781e60187aa260100c7ef63, /* 1910 */
128'h7713b7f5367d0785feb71ce30007c703, /* 1911 */
128'h87aa0007069b40e7873b47a1c31d0075, /* 1912 */
128'h1793faf5078536fdfcb81ce30007c803, /* 1913 */
128'h00b7e733008597938e1d953e93810207, /* 1914 */
128'h8edd00365713020796938fd901071793, /* 1915 */
128'h1fe30007c703d24d8a1deb1187aa2701, /* 1916 */
128'h008785130007b803bfcd367d0785f8b7, /* 1917 */
128'h1be30785f8b712e30007c70300d80a63, /* 1918 */
128'h4703e7a9419cb7f1377d87aabfa5fef5, /* 1919 */
128'h27970015470308f71163030007930005, /* 1920 */
128'h8a850006c68300e786b30f2787930000, /* 1921 */
128'h1b63078006930ff777130207071bc689, /* 1922 */
128'h0447f7930007c78397ba0025470304d7, /* 1923 */
128'h470302f71c6347c14198c19c47c1c3b1, /* 1924 */
128'h27170015478302f71663030007930005, /* 1925 */
128'hc7098b0500074703973e0a2707130000, /* 1926 */
128'h00e79363078007130ff7f7930207879b, /* 1927 */
128'he8221101bf6d47a9bf7d47a180820509, /* 1928 */
128'h00c16583f63ff0efc632ec06006c842e, /* 1929 */
128'h079b0005470305e80813000028174681, /* 1930 */
128'h9863044678930006460300f806330007, /* 1931 */
128'h7893808261058536644260e2ec050008, /* 1932 */
128'h86b3feb7f4e3fd07879b00088b630046, /* 1933 */
128'hfe07079bc6098a09b7d196be050502d5, /* 1934 */
128'h7139b7e1e008b7cdfc97879b0ff7f793, /* 1935 */
128'h842ae42e00063023f04afc06f426f822, /* 1936 */
128'h744270e25529e90165a2b0dff0ef84b2, /* 1937 */
128'h8522082c892a862e80826121790274a2, /* 1938 */
128'hcb010007c703fe8782e367e2f5dff0ef, /* 1939 */
128'he088fcf718e347a9fd279be307858f81, /* 1940 */
128'h00e6846302d0071300054683b7e94501, /* 1941 */
128'h60a2f23ff0efe40605051141f2dff06f, /* 1942 */
128'h842ee406e02211418082014140a00533, /* 1943 */
128'h04630007c70304b00693601cf0dff0ef, /* 1944 */
128'h60a202d70e630470069300e6ea6302d7, /* 1945 */
128'h069302d7076304d00693808201416402, /* 1946 */
128'h052a069007130017c683fed716e306b0, /* 1947 */
128'h00e69863042007130027c683fce69fe3, /* 1948 */
128'hbfd50789bff1052a052ab7e9e01c078d, /* 1949 */
128'he0fff0efc632ec06006c842ee8221101, /* 1950 */
128'h4703f0a8081300002817468100c16583, /* 1951 */
128'h78930006460300f806330007079b0005, /* 1952 */
128'h61058536644260e2ec05000898630446, /* 1953 */
128'hf4e3fd07879b00088b63004678938082, /* 1954 */
128'hc6098a09b7d196be050502d586b3feb7, /* 1955 */
128'he008b7cdfc97879b0ff7f793fe07079b, /* 1956 */
128'h601cf87ff0ef842ee406e0221141b7e1, /* 1957 */
128'h00e6ea6302d704630007c70304b00693, /* 1958 */
128'h80820141640260a202d70e6304700693, /* 1959 */
128'hfed716e306b0069302d7076304d00693, /* 1960 */
128'hc683fce69fe3052a069007130017c683, /* 1961 */
128'hb7e9e01c078d00e69863042007130027, /* 1962 */
128'he406e0221141bfd50789bff1052a052a, /* 1963 */
128'hfff5c70300a405b395bff0efe589842a, /* 1964 */
128'h4703973efff58513e307879300002797, /* 1965 */
128'h80820141557d640260a2e7198b110007, /* 1966 */
128'h00074703973e00054703fea47ae3157d, /* 1967 */
128'h014105054581462960a26402f77d8b11, /* 1968 */
128'h00a107a31141fa5ff06f4581d7dff06f, /* 1969 */
128'h47978082014100e1550300a107238121, /* 1970 */
128'h9201160291811582639c2c2787930000, /* 1971 */
128'h0005470345a946254781aa5ff06f95be, /* 1972 */
128'h67630ff6f693fd07069b8082853ee319, /* 1973 */
128'hbff90505fd07879b9fb902f587bb00d6, /* 1974 */
128'hf86347a500a04563842ee406e0221141, /* 1975 */
128'h4529fe7ff0ef357d02b455bb45a900b7, /* 1976 */
128'h006f03050513014160a2640202a4753b, /* 1977 */
128'h24f734230000471707e2081007935000, /* 1978 */
128'h4417e8221101808224f7342300004717, /* 1979 */
128'h600885aa84ae862ee42623a404130000, /* 1980 */
128'h6442e00c95a660e2600ca15ff0efec06, /* 1981 */
128'h210787930000479711018082610564a2, /* 1982 */
128'h6380e82260901fe4849300004497e426, /* 1983 */
128'hd0ef85a29c11ec067b85051300003517, /* 1984 */
128'h862286aa608ce63fc0ef85a26088b87f, /* 1985 */
128'h00003517b6dfd0ef7b05051300003517, /* 1986 */
128'hef65051300000517b61fd0ef7bc50513, /* 1987 */
128'h05b364a260e2644200055e63857f90ef, /* 1988 */
128'hb39fd06f61057ae505130000351740a0, /* 1989 */
128'he02211416680006f610564a260e26442, /* 1990 */
128'h60a2557d00850363878fa0ef8432e406, /* 1991 */
128'h8413f222716980824501808201416402, /* 1992 */
128'h892eea4aee26f606852289aae64e0125, /* 1993 */
128'hf72ff0ef852600a404b30505f7eff0ef, /* 1994 */
128'h1ff00793fff5071be93ff0ef95260505, /* 1995 */
128'hf0ef852212a7a2230000479704e7ee63, /* 1996 */
128'hf42ff0ef524505130000351784aaf50f, /* 1997 */
128'hf32ff0ef852204a7f2630ff007939526, /* 1998 */
128'h05b3f24ff0ef5065051300003517842a, /* 1999 */
128'h70b2a8bfd0ef71e505130000351700a4, /* 2000 */
128'h200007938082615569b2695264f27412, /* 2001 */
128'h458110000613b7550cf7242300004717, /* 2002 */
128'h850a4c25859300003597863ff0ef850a, /* 2003 */
128'h00f7096302f0079301294703deaff0ef, /* 2004 */
128'h85a2dfaff0ef850a6f05859300003597, /* 2005 */
128'h43900827879300004797df2ff0ef850a, /* 2006 */
128'h0793a1bfd0ef6d65051300003517858a, /* 2007 */
128'h471706f7352300004717451107e20810, /* 2008 */
128'h932300004797d85ff0ef06f735230000, /* 2009 */
128'he2a79d2300004797d77ff0ef4501e4a7, /* 2010 */
128'heb1ff0ef854ee2e58593000045974611, /* 2011 */
128'he8221101b79102f71523000047174785, /* 2012 */
128'h892a08c7df638432478de04ae426ec06, /* 2013 */
128'h956325010004d783d37ff0ef84ae450d, /* 2014 */
128'hd783d21ff0efffa555030000451708a7, /* 2015 */
128'h00448513ffc4059b06a79a6325010024, /* 2016 */
128'h932300004797d05ff0ef4511dabff0ef, /* 2017 */
128'h4611cf1ff0effca5550300004517dca7, /* 2018 */
128'hda85859300004597daa7992300004797, /* 2019 */
128'h00004597256000ef4535e2bff0ef854a, /* 2020 */
128'h00ef02000513d1bff0ef4515fa05d583, /* 2021 */
128'h27850007d783f8a78793000047972400, /* 2022 */
128'hf707879300004797f6f71e2300004717, /* 2023 */
128'h5e050513000035170087cf63278d439c, /* 2024 */
128'hf06f6105690264a260e26442905fd0ef, /* 2025 */
128'h717980826105690264a2644260e2d49f, /* 2026 */
128'hc78300f10fa347090105c783f022f406, /* 2027 */
128'h470d00e78e6301e1578300f10f230115, /* 2028 */
128'h5c0505130000351770a2740202e78a63, /* 2029 */
128'h5985051300003517842a8b3fd06f6145, /* 2030 */
128'h614570a265a2740285228a3fd0efe42e, /* 2031 */
128'hf06f614505c170a241907402d8bff06f, /* 2032 */
128'h30232291342322813823dc010113ebff, /* 2033 */
128'h0028218006134581893284ae842a2321, /* 2034 */
128'h08282040061385a6e60ff0ef22113c23, /* 2035 */
128'hf63ff0ef8522002cea2ff0efe802c44a, /* 2036 */
128'h22013903228134832301340323813083, /* 2037 */
128'hcb81e867d78300004797808224010113, /* 2038 */
128'h8082cf3ff06fc6e58593000045974611, /* 2039 */
128'h7763878e1041e703504000efe4061141, /* 2040 */
128'h10a7a22310e1a02327051001a70300e5, /* 2041 */
128'h01418d5d91011782150260a21007e783, /* 2042 */
128'h84aae426e822ec061101808245018082, /* 2043 */
128'h07b33e800793440000ef842afc1ff0ef, /* 2044 */
128'h8d0502a7d533644260e29101150202f4, /* 2045 */
128'hf95ff0efe022e40611418082610564a2, /* 2046 */
128'h07b324078793000f47b7414000ef842a, /* 2047 */
128'h02a7d533014191011502640260a202f4, /* 2048 */
128'hf0ef84aae04ae426e822ec0611018082, /* 2049 */
128'h000f443702a485333e2000ef892af63f, /* 2050 */
128'hf45ff0ef0405944a0285543324040413, /* 2051 */
128'h80826105690264a2644260e2fe856ee3, /* 2052 */
128'h842ae04aec06e822009894b7e4261101, /* 2053 */
128'h0433854a89260084f363892268048493, /* 2054 */
128'h690264a2644260e2f47dfa1ff0ef4124, /* 2055 */
128'h808200054503808200b5002380826105, /* 2056 */
128'h07378082020575130147c503100007b7, /* 2057 */
128'h00a70023dfe50207f793014747831000, /* 2058 */
128'h8623f800071300078223100007b78082, /* 2059 */
128'h8623470d0007822300e78023476d00e7, /* 2060 */
128'h88230200071300e78423fc70071300e7, /* 2061 */
128'h00044503842ae406e0221141808200e7, /* 2062 */
128'h0405fa5ff0ef80820141640260a2e509, /* 2063 */
128'h811100f57713d567879300002797b7f5, /* 2064 */
128'h00e580a30007c7830007470397aa973e, /* 2065 */
128'h8121842a002ce8221101808200f58023, /* 2066 */
128'h4503f65ff0ef00814503fd1ff0efec06, /* 2067 */
128'hfb7ff0ef0ff47513002cf5dff0ef0091, /* 2068 */
128'hf43ff0ef00914503f4bff0ef00814503, /* 2069 */
128'he84aec26f022717980826105644260e2, /* 2070 */
128'h7513002c0089553b54e14461892af406, /* 2071 */
128'hf13ff0ef346100814503f81ff0ef0ff5, /* 2072 */
128'h740270a2fe9410e3f0bff0ef00914503, /* 2073 */
128'he84aec26f022717980826145694264e2, /* 2074 */
128'h002c0089553354e103800413892af406, /* 2075 */
128'hf0ef346100814503f3fff0ef0ff57513, /* 2076 */
128'h70a2fe9410e3ec9ff0ef00914503ed1f, /* 2077 */
128'hec06002c110180826145694264e27402, /* 2078 */
128'h00914503ea7ff0ef00814503f13ff0ef, /* 2079 */
128'h8793000047978082610560e2e9fff0ef, /* 2080 */
128'hec4efc06f04af426f8227139439ce2e7, /* 2081 */
128'h05130000451702b7856384b2842e892a, /* 2082 */
128'ha12300004797c10d2501f3afb0efbd65, /* 2083 */
128'h8082612169e2790274a2744270e2e0a7, /* 2084 */
128'h85ca86260074def723230000471757fd, /* 2085 */
128'hc50d2501814fb0efba05051300004517, /* 2086 */
128'h85a6049675634632dca7a62300004797, /* 2087 */
128'h47174785d0cfd0ef2385051300003517, /* 2088 */
128'h591be05ff0ef4521b775daf727230000, /* 2089 */
128'h791323278793000037970009099b00c4, /* 2090 */
128'h10ef854ede7ff0ef00094503993e0039, /* 2091 */
128'hbf95d687a923000047979c25bf5d3200, /* 2092 */
128'h2085051300003517842a85aae0221141, /* 2093 */
128'h25730ff0000f0000100fcb2fd0efe406, /* 2094 */
128'hbb8585930000259760a264028322f140, /* 2095 */
128'hef058593000035974605114183020141, /* 2096 */
128'hd79fa0efe022e406d305051300004517, /* 2097 */
128'h60a264021ec5051300003517c9112501, /* 2098 */
128'hd0ef1fa5051300003517c62fd06f0141, /* 2099 */
128'h0000451720c58593000035974605c56f, /* 2100 */
128'h00003517c5112501d9bfa0efab450513, /* 2101 */
128'hd0ef0825051300003517b7e120450513, /* 2102 */
128'ha12300004797e985051300000517c26f, /* 2103 */
128'h842a90cf90efca07ab2300004797cc07, /* 2104 */
128'hcf81439cca8787930000479700054863, /* 2105 */
128'h058505130000351760a26402408005b3, /* 2106 */
128'hb0efa4a5051300004517be2fd06f0141, /* 2107 */
128'hbfb91b25051300003517c5112501b9af, /* 2108 */
128'hcb9fa0ef4501e2658593000035974605, /* 2109 */
128'h8522b7811ac5051300003517c5112501, /* 2110 */
128'he40625011141900200000023ee1ff0ef, /* 2111 */
128'h808224050513000f4537a001d69ff0ef, /* 2112 */
128'h157d631cc1c707130000471780824501, /* 2113 */
128'h10d00513e30895360017869300756513, /* 2114 */
128'hec06e822110102b506338082953e055e, /* 2115 */
128'h45816622c509842afd1ff0efe4328532, /* 2116 */
128'h808280826105644260e28522944ff0ef, /* 2117 */
128'hb28fd0efe40614650513000035171141, /* 2118 */
128'h80820141450160a2ee5fc0ef20000537, /* 2119 */
128'h553347a9b00025738082450180824501, /* 2120 */
128'h351785aa862e86b287361141808202f5, /* 2121 */
128'hf0ef4505aecfd0efe406132505130000, /* 2122 */
128'hf0efe406952e842ae0221141a001cbbf, /* 2123 */
128'h01418d7d640260a29522408007b3f57f, /* 2124 */
128'h71798082450580824505808245058082, /* 2125 */
128'h0096186300c684bb842ef406ec26f022, /* 2126 */
128'h852285b280826145450164e2740270a2, /* 2127 */
128'hbff92605200404136622e37fc0efe432, /* 2128 */
128'h80828082808245098082450980824509, /* 2129 */
128'h1101bbbff06f80824501808245018082, /* 2130 */
128'h00d584b3003796934781e426e822ec06, /* 2131 */
128'h450164a2644260e200c7986300d50433, /* 2132 */
128'h600c02e8036360980004380380826105, /* 2133 */
128'h8626a2afd0ef0a650513000035176090, /* 2134 */
128'ha001a1afd0ef0be505130000351785a2, /* 2135 */
128'h051300003517892ae0ca711dbf5d0785, /* 2136 */
128'he862ec5ef05af456f852fc4ee8a20be5, /* 2137 */
128'h3a179eafd0ef44018b2ee466e4a6ec86, /* 2138 */
128'h49930b2b8b9300003b970aaa0a130000, /* 2139 */
128'hd0ef85524ac10b6c0c1300003c17fff9, /* 2140 */
128'h87ca9bafd0ef855e85e600040c9b9c6f, /* 2141 */
128'h856285e69acfd0ef8552036498634481, /* 2142 */
128'h17e3040502b49b63458187ca9a4fd0ef, /* 2143 */
128'h450198afd0ef0de5051300003517fd54, /* 2144 */
128'h00349713c689873e8a85008486b3a889, /* 2145 */
128'h86b3bf5d07a104856398e39840e98733, /* 2146 */
128'h873300359713c689873e8a8563900085, /* 2147 */
128'h0405051300003517058e02e60d6340e9, /* 2148 */
128'h938fd0ef06c5051300003517944fd0ef, /* 2149 */
128'h7aa27a4279e2690664a6644660e6557d, /* 2150 */
128'h07a10585808261256ca26c426be27b02, /* 2151 */
128'h020005138aaa6a05fc56e0d27159bfa5, /* 2152 */
128'he8caf0a2f486f062f45ef85ae4ceeca6, /* 2153 */
128'hb3fff0ef44818bb28b2ee46ee86aec66, /* 2154 */
128'h97933a2c0c1300003c179c4a0a134981, /* 2155 */
128'h351703749b6300fb0cb300fa8db30034, /* 2156 */
128'h694670a674068befd0ef03a505130000, /* 2157 */
128'h86266da26d426ce27c027ba26a0669a6, /* 2158 */
128'he33ff06f61657ae285567b4264e685da, /* 2159 */
128'hbd1fe0ef8d2abd7fe0ef842abddfe0ef, /* 2160 */
128'h1d1b0105151b0344f7b3bcbfe0ef892a, /* 2161 */
128'h91011402150201a4643300a96533010d, /* 2162 */
128'hf0ef4521ef8100adb02300acb0238d41, /* 2163 */
128'hf0ef0007c50397e20039f7930985aadf, /* 2164 */
128'hf822fc06e032e42e7139b7ad0485a9df, /* 2165 */
128'he0ef842ab75fe0ef89aaec4ef04af426, /* 2166 */
128'h151bb63fe0ef84aab69fe0ef892ab6ff, /* 2167 */
128'h65a2660215028fc18d450109179b0105, /* 2168 */
128'h00e588330037971347818d5d91011782, /* 2169 */
128'h854e790274a270e2744200c79c63974e, /* 2170 */
128'h8ea907856314d79ff06f6121863e69e2, /* 2171 */
128'h7139b7f100e830238f2900083703e314, /* 2172 */
128'h89aaec4ef04af426f822fc06e032e42e, /* 2173 */
128'haf1fe0ef892aaf7fe0ef842aafdfe0ef, /* 2174 */
128'h8d450109179b0105151baebfe0ef84aa, /* 2175 */
128'h47818d5d9101178265a2660215028fc1, /* 2176 */
128'h744200c79c63974e00e5883300379713, /* 2177 */
128'hf06f6121863e69e2854e790274a270e2, /* 2178 */
128'h8f0900083703e3148e8907856314d01f, /* 2179 */
128'hf822fc06e032e42e7139b7f100e83023, /* 2180 */
128'he0ef842aa85fe0ef89aaec4ef04af426, /* 2181 */
128'h151ba73fe0ef84aaa79fe0ef892aa7ff, /* 2182 */
128'h65a2660215028fc18d450109179b0105, /* 2183 */
128'h00e588330037971347818d5d91011782, /* 2184 */
128'h854e790274a270e2744200c79c63974e, /* 2185 */
128'h86b307856314c89ff06f6121863e69e2, /* 2186 */
128'h00e8302302a7073300083703e31402a6, /* 2187 */
128'hf04af426f822fc06e032e42e7139b7e1, /* 2188 */
128'h892aa03fe0ef842aa09fe0ef89aaec4e, /* 2189 */
128'h179b0105151b9f7fe0ef84aa9fdfe0ef, /* 2190 */
128'h9101178265a2660215028fc18d450109, /* 2191 */
128'h9c63974e00e588330037971347818d5d, /* 2192 */
128'h863e69e2854e790274a270e2744200c7, /* 2193 */
128'hd6b3078563144505e111c0dff06f6121, /* 2194 */
128'h00e8302302a7573300083703e31402a6, /* 2195 */
128'hf04af426f822fc06e032e42e7139b7d1, /* 2196 */
128'h892a983fe0ef842a989fe0ef89aaec4e, /* 2197 */
128'h179b0105151b977fe0ef84aa97dfe0ef, /* 2198 */
128'h9101178265a2660215028fc18d450109, /* 2199 */
128'h9c63974e00e588330037971347818d5d, /* 2200 */
128'h863e69e2854e790274a270e2744200c7, /* 2201 */
128'h3703e3148ec907856314b8dff06f6121, /* 2202 */
128'he032e42e7139b7f100e830238f490008, /* 2203 */
128'h911fe0ef89aaec4ef04af426f822fc06, /* 2204 */
128'he0ef84aa905fe0ef892a90bfe0ef842a, /* 2205 */
128'h15028fc18d450109179b0105151b8fff, /* 2206 */
128'h0037971347818d5d9101178265a26602, /* 2207 */
128'h74a270e2744200c79c63974e00e58833, /* 2208 */
128'h6314b15ff06f6121863e69e2854e7902, /* 2209 */
128'h00e830238f6900083703e3148ee90785, /* 2210 */
128'hf04af426f822fc06e032e42e7139b7f1, /* 2211 */
128'h892a893fe0ef842a899fe0ef89aaec4e, /* 2212 */
128'h179b0105151b887fe0ef84aa88dfe0ef, /* 2213 */
128'h9081178265a2660214828fc18cc90109, /* 2214 */
128'h1c6396ae00d988330037169347018fc5, /* 2215 */
128'h863a69e2854e790274a270e2744200c7, /* 2216 */
128'h00a83023e28800f70533a9dff06f6121, /* 2217 */
128'h051300003517892ae8ca7159bfc90705, /* 2218 */
128'hf062f45ef85afc56e0d2e4cef0a2b9e5, /* 2219 */
128'hcc9fc0ef44018b3289aeec66eca6f486, /* 2220 */
128'hb90b8b9300003b97b88a0a1300003a17, /* 2221 */
128'hc0ef855204000a93b98c0c1300003c17, /* 2222 */
128'hc99fc0ef8885855e85a2fff44493ca7f, /* 2223 */
128'h00f905b30036179314fd460140900cb3, /* 2224 */
128'h85a2c7bfc0efe43285520566186397ce, /* 2225 */
128'ha03ff0ef854a85ce6622c73fc0ef8562, /* 2226 */
128'h051300003517fb541be32405e12984aa, /* 2227 */
128'h64e669468526740670a6c53fc0efba65, /* 2228 */
128'h61656ce27c027ba27b427ae26a0669a6, /* 2229 */
128'he198e3988726c2918766001676938082, /* 2230 */
128'h351784aaeca67159bfc154fdbf590605, /* 2231 */
128'hfc56e0d2e4cee8caf0a2aca505130000, /* 2232 */
128'h8ab2892ee86af486ec66f062f45ef85a, /* 2233 */
128'h3b17ab29899300003997bf3fc0ef4401, /* 2234 */
128'h3c17db2b8b9300003b97db2b0b130000, /* 2235 */
128'h0a13ab2c8c9300003c97aaac0c130000, /* 2236 */
128'hbd03cba500147793bc1fc0ef854e0400, /* 2237 */
128'hfffd45134601baffc0ef856285a2000b, /* 2238 */
128'h854e05561c6397ca00f485b300361793, /* 2239 */
128'h6622b8bfc0ef856685a2b93fc0efe432, /* 2240 */
128'h1ae32405e5298d2a91bff0ef852685ca, /* 2241 */
128'h70a6b6bfc0efabe5051300003517fb44, /* 2242 */
128'h7b427ae26a0669a6694664e6856a7406, /* 2243 */
128'h000b3d03808261656d426ce27c027ba2, /* 2244 */
128'he198e398872ac291876a00167693bf49, /* 2245 */
128'h3517842ae8a2711db7e15d7db7790605, /* 2246 */
128'hf05af456f852e0cae4a69da505130000, /* 2247 */
128'hc0ef4c018ab284aefc4eec86e862ec5e, /* 2248 */
128'h0b1300003b179c69091300003917b07f, /* 2249 */
128'h854a10000a139d6b8b9300003b979ceb, /* 2250 */
128'had9fc0ef855a85ce000c099bae5fc0ef, /* 2251 */
128'h17130187e7b38fd9010c1793008c1713, /* 2252 */
128'h8fd9028c17138fd9020c17138fd9018c, /* 2253 */
128'h171346018fd9038c17138fd9030c1713, /* 2254 */
128'he432854a05561763972600e406b30036, /* 2255 */
128'h85a66622a8dfc0ef855e85cea95fc0ef, /* 2256 */
128'hf94c19e30c05e91d89aa81dff0ef8522, /* 2257 */
128'h644660e6a6dfc0ef9c05051300003517, /* 2258 */
128'h6be27b027aa27a4279e2690664a6854e, /* 2259 */
128'h59fdb74d0605e29ce31c808261256c42, /* 2260 */
128'h8f0505130000351784aaf4a67119bff1, /* 2261 */
128'hf862fc5ee0dae4d6e8d2eccef0caf8a2, /* 2262 */
128'hc0ef44018b32892eec6efc86f06af466, /* 2263 */
128'h8c9300003c978d6a0a1300003a17a17f, /* 2264 */
128'h00003d1703f00c13498507f00b938dec, /* 2265 */
128'h85a29ebfc0ef855208000a938dcd0d13, /* 2266 */
128'h95b300e99733408b873b9e3fc0ef8566, /* 2267 */
128'h1a6397ca00f486b30036179346010089, /* 2268 */
128'hc0ef856a85a29bffc0efe43285520566, /* 2269 */
128'he1398daaf46ff0ef852685ca66229b7f, /* 2270 */
128'hc0ef8ea5051300003517fb541be32405, /* 2271 */
128'h6a4669e6790674a6856e744670e6997f, /* 2272 */
128'h61096de27d027ca27c427be26b066aa6, /* 2273 */
128'he398bf610605e28ce38c008c66638082, /* 2274 */
128'h351784aaf4a67119b7f15dfdbfe5e298, /* 2275 */
128'he4d6e8d2eccef0caf8a280a505130000, /* 2276 */
128'h892eec6efc86f06af466f862fc5ee0da, /* 2277 */
128'h7f0a0a1300002a17931fc0ef44018b32, /* 2278 */
128'h0c13498507f00b937f8c8c9300002c97, /* 2279 */
128'h855208000a937f6d0d1300002d1703f0, /* 2280 */
128'h408b87bb8fdfc0ef856685a2905fc0ef, /* 2281 */
128'hfff6c693fff7c793008996b300f997b3, /* 2282 */
128'h05661a63974a00e485b3003617134601, /* 2283 */
128'h8c9fc0ef856a85a28d1fc0efe4328552, /* 2284 */
128'h2405e1398daae58ff0ef852685ca6622, /* 2285 */
128'h8a9fc0ef7fc5051300002517fb5417e3, /* 2286 */
128'h6aa66a4669e6790674a6856e744670e6, /* 2287 */
128'h808261096de27d027ca27c427be26b06, /* 2288 */
128'he19ce31cbf610605e194e314008c6663, /* 2289 */
128'h0000251784aaf4a67119b7f15dfdbfe5, /* 2290 */
128'he0dae4d6e8d2eccef0caf8a271c50513, /* 2291 */
128'h8a32892eec6efc86f06af466f862fc5e, /* 2292 */
128'h2c177029899300002997843fc0ef4401, /* 2293 */
128'h08100b134d0507f00a9370ac0c130000, /* 2294 */
128'hc0ef854e704c8c9300002c9703f00b93, /* 2295 */
128'h07bb408a873b80ffc0ef856285a2817f, /* 2296 */
128'h0024079b8f5d00ed173300fd17b3408b, /* 2297 */
128'hc313fff748938fd5008d16b300fd17b3, /* 2298 */
128'h1c6396ca00d48533003616934601fff7, /* 2299 */
128'hc0ef856685a2fcefc0efe432854e0546, /* 2300 */
128'hed298daad56ff0ef852685ca6622fc6f, /* 2301 */
128'h051300002517f8f41be3080007932405, /* 2302 */
128'h790674a6856e744670e6fa2fc0ef6f65, /* 2303 */
128'h7d027ca27c427be26b066aa66a4669e6, /* 2304 */
128'h859a008bea6300167813808261096de2, /* 2305 */
128'h85c6b7610605e10ce28c85be00081363, /* 2306 */
128'hf0ca7119bf755dfdbfc585bafe081be3, /* 2307 */
128'hfc5ee8d2ecce6065051300002517892a, /* 2308 */
128'he0dae4d6f4a6f8a2fc86ec6ef06af466, /* 2309 */
128'h00002a17f2cfc0ef4b81e03289aef862, /* 2310 */
128'h00002d175f4c8c9300002c975eca0a13, /* 2311 */
128'h003b949b01779c3347854da15fcd0d13, /* 2312 */
128'h856685da00848b3bf00fc0ef85524401, /* 2313 */
128'h0036171367824601fffc4a93ef4fc0ef, /* 2314 */
128'hc0efe432855206f61063974e00e90833, /* 2315 */
128'h854a85ce6622ecefc0ef856a85daed6f, /* 2316 */
128'hfbb41be38c562405e9318b2ac5eff0ef, /* 2317 */
128'h051300002517fafb90e3040007932b85, /* 2318 */
128'h790674a6855a744670e6ea2fc0ef5f65, /* 2319 */
128'h7d027ca27c427be26b066aa66a4669e6, /* 2320 */
128'h85d6e11185e200167513808261096de2, /* 2321 */
128'h7175b7e95b7db749060500b83023e30c, /* 2322 */
128'h698502000513892e84aaf4cef8cafca6, /* 2323 */
128'he122e506fc66e0e2e4dee8daecd6f0d2, /* 2324 */
128'h3c174a01892ff0ef4a81e032f46ef86a, /* 2325 */
128'h8c9300003c979c498993132c0c130000, /* 2326 */
128'h003d969367824d214d818bca8b268eec, /* 2327 */
128'hba2ff0ef852685ca866e04fd956396da, /* 2328 */
128'h5705051300002517020a0863ed45842a, /* 2329 */
128'h79a6794674e6640a60aa8522df4fc0ef, /* 2330 */
128'h7da27d427ce26c066ba66b466ae67a06, /* 2331 */
128'he0efec36b7758ba68b4a4a0580826149, /* 2332 */
128'he42a902fe0efe82a908fe0ef842a90ef, /* 2333 */
128'h161b8d5d0105151b664267a28fcfe0ef, /* 2334 */
128'h37978d4166e29101140215028c510106, /* 2335 */
128'hc683018786b34781e28808a7b9230000, /* 2336 */
128'h00d600230ff6f693078500fb86330006, /* 2337 */
128'he0ef4521ef910ba1033df7b3ffa795e3, /* 2338 */
128'hc50397e68b8d00078a9b001a879bfbdf, /* 2339 */
128'h7175bfa1547dbf0d0d85fa9fe0ef0007, /* 2340 */
128'h6a050200051389ae892af0d2f4cef8ca, /* 2341 */
128'he506f86afc66e0e2e4dee8daecd6fca6, /* 2342 */
128'h34974a81f73fe0ef4b018cb2f46ee122, /* 2343 */
128'h0d1300002d179c4a0a1301a484930000, /* 2344 */
128'h00fc06b3003d97934d818c4e8bca7ced, /* 2345 */
128'ha82ff0ef854a85ce866e059d956397de, /* 2346 */
128'h4505051300002517020a8863e579842a, /* 2347 */
128'h79a6794674e6640a60aa8522cd4fc0ef, /* 2348 */
128'h7da27d427ce26c066ba66b466ae67a06, /* 2349 */
128'he836ec3eb7758c4a8bce4a8580826149, /* 2350 */
128'hfe1fd0efe42afe7fd0ef842afedfd0ef, /* 2351 */
128'h161b0105151b67026622fdbfd0efe02a, /* 2352 */
128'h37978d419101140215028c518d590106, /* 2353 */
128'h0004d783e38866c267e2f6a7bd230000, /* 2354 */
128'h93c117c20024d78300f6902393c117c2, /* 2355 */
128'h00f6922393c117c20044d78300f69123, /* 2356 */
128'h034df7b300f6932393c117c20064d783, /* 2357 */
128'h00078b1b001b079be87fe0ef4521ef91, /* 2358 */
128'hbf290d85e73fe0ef0007c50397ea8b8d, /* 2359 */
128'h86138932f8ca717580826505b789547d, /* 2360 */
128'h251785aa962a84ae842afca6e122fff5, /* 2361 */
128'he4dee8daecd6f0d2f4ce372505130000, /* 2362 */
128'hbd8fc0efec36e506f46ef86afc66e0e2, /* 2363 */
128'h99a20034d793e83e0014d9930044d793, /* 2364 */
128'h2b9735ab0b1300002b1744854a81e43e, /* 2365 */
128'h2c9735ac0c1300002c1735ab8b930000, /* 2366 */
128'h2d97362d0d1300002d1735ac8c930000, /* 2367 */
128'h7863e72a0a1300003a17362d8d930000, /* 2368 */
128'h60aab7afc0ef35650513000025170299, /* 2369 */
128'h6b466ae67a0679a6794674e68556640a, /* 2370 */
128'h85a6808261497da27d427ce26c066ba6, /* 2371 */
128'hc0ef855e85ca00090663b52fc0ef855a, /* 2372 */
128'hb38fc0ef856a85e6b40fc0ef8562b46f, /* 2373 */
128'hb28fc0ef856eed15920ff0ef852265a2, /* 2374 */
128'hc58d000a358302f749636762010a2783, /* 2375 */
128'h008a3783b0cfc0ef2d85051300002517, /* 2376 */
128'h2c850513000025179782852285ce6642, /* 2377 */
128'h0805051300002517b7e94a89af4fc0ef, /* 2378 */
128'h0513000025177179bfa10485ae4fc0ef, /* 2379 */
128'hc19fe0efe44ee84aec26f022f4062b65, /* 2380 */
128'hab8fc0ef2b4505130000251704000593, /* 2381 */
128'h00002517aacfc0ef2d05051300002517, /* 2382 */
128'h0305051300002517aa0fc0ef2f450513, /* 2383 */
128'h95b3497901f499934441a92fc0ef4485, /* 2384 */
128'he6dff0ef240501358533460546850084, /* 2385 */
128'h614569a2694264e2740270a2ff2417e3, /* 2386 */
128'h46814881470100c5131b460580828082, /* 2387 */
128'h000780234000081387f245a901f61e13, /* 2388 */
128'h802397aa0007802397aa0007802397aa, /* 2389 */
128'h02b71d632705fe0813e397aa387d0007, /* 2390 */
128'h86b33e800513c00026f38e15c0202673, /* 2391 */
128'h45bb02c747334000059302a687334116, /* 2392 */
128'h05130000251702a7473302a767b302b3, /* 2393 */
128'h28f3c02026f3fac710e39f2fc06f28e5, /* 2394 */
128'h4505f7bff0ef4501e4061141bf51c000, /* 2395 */
128'hf69ff0ef4511f6fff0ef4509f75ff0ef, /* 2396 */
128'h1502bff1f5dff0ef4541f63ff0ef4521, /* 2397 */
128'h6388400007b78082e388400007b79101, /* 2398 */
128'h25016b880007b823400007b780822501, /* 2399 */
128'h0085979b808225017b88400007b78082, /* 2400 */
128'h2581f7888d51400007b70106161b8d5d, /* 2401 */
128'h06b73e80079300b7ef63400007374781, /* 2402 */
128'h400007b7ffe537fdc3198b097a984000, /* 2403 */
128'hbfe1f710069127850006e60380827388, /* 2404 */
128'h551b00b7d863842a4785e406e0221141, /* 2405 */
128'h00002797883dfebff0ef250135fd0045, /* 2406 */
128'h014160a2640200044503943e20478793, /* 2407 */
128'h67050185579b9d3d00b007b7a1ffe06f, /* 2408 */
128'h8fd9058565133007071311010085151b, /* 2409 */
128'hc43e454d458946010034842ec62ae822, /* 2410 */
128'hf0ef454d460100344589f5bff0efec06, /* 2411 */
128'h802300f556b357610380079385a2f4ff, /* 2412 */
128'h6105644260e2fee79ae3058537e100d5, /* 2413 */
128'hec56f052f44ef84afc26e0a2715d8082, /* 2414 */
128'h0ab7ff86099b440189328a2e84aae486, /* 2415 */
128'hf79ff0ef002c033466630144053b4000, /* 2416 */
128'hecbfd0ef92018526002c16024089063b, /* 2417 */
128'h61616ae27a0279a2794274e2640660a6, /* 2418 */
128'h178200c4579b2421f51ff0ef85a68082, /* 2419 */
128'h000025171141bf6d00fab02304a19381, /* 2420 */
128'h05130000051783efc0efe406c9c50513, /* 2421 */
128'h40a005b360a200055c63d35f70eff885, /* 2422 */
128'h60a281afc06f0141c905051300002517, /* 2423 */
128'he06f1a25051300002517b4ffe06f0141, /* 2424 */
128'he852ec4ef04af426f822fc067139957f, /* 2425 */
128'h0e0505130000251790ffe0efe05ae456, /* 2426 */
128'h091300002917080009b74401935fe0ef, /* 2427 */
128'h0004059b6390078e013407b344950de9, /* 2428 */
128'hda0f80effe9416e3fc1fb0ef0405854a, /* 2429 */
128'h2a97400004b727eb0b1300002b174901, /* 2430 */
128'h49910caa0a1300002a170baa8a930000, /* 2431 */
128'h608ce09c090585560007c783016907b3, /* 2432 */
128'h0004b823f7dfb0ef8622240125816080, /* 2433 */
128'h7413fd391be3f6ffb0ef25818552688c, /* 2434 */
128'h0000071702f7646347190054579b0ff4, /* 2435 */
128'h2517878297ba439c97ba078a65470713, /* 2436 */
128'haa9fe0ef8522f3ffb0ef08a505130000, /* 2437 */
128'h8522f2bfb0ef0865051300002517a001, /* 2438 */
128'hb0ef0825051300002517b7f5edbff0ef, /* 2439 */
128'h0805051300002517bfe9c37ff0eff17f, /* 2440 */
128'h051300002517b7e1e14f80eff05fb0ef, /* 2441 */
128'h00000000bf5dd0fff0efef3fb0ef07e5, /* 2442 */
128'h00000000000000000000000000000000, /* 2443 */
128'h00000000000000000000000000000000, /* 2444 */
128'h00000000000000000000000000000000, /* 2445 */
128'h00000000000000000000000000000000, /* 2446 */
128'h00000000000000000000000000000000, /* 2447 */
128'h08082828282828080808080808080808, /* 2448 */
128'h08080808080808080808080808080808, /* 2449 */
128'h101010101010101010101010101010a0, /* 2450 */
128'h10101010101004040404040404040404, /* 2451 */
128'h01010101010101010141414141414110, /* 2452 */
128'h10101010100101010101010101010101, /* 2453 */
128'h02020202020202020242424242424210, /* 2454 */
128'h08101010100202020202020202020202, /* 2455 */
128'h00000000000000000000000000000000, /* 2456 */
128'h00000000000000000000000000000000, /* 2457 */
128'h101010101010101010101010101010a0, /* 2458 */
128'h10101010101010101010101010101010, /* 2459 */
128'h01010101010101010101010101010101, /* 2460 */
128'h02010101010101011001010101010101, /* 2461 */
128'h02020202020202020202020202020202, /* 2462 */
128'h02020202020202021002020202020202, /* 2463 */
128'hc1bdceee242070dbe8c7b756d76aa478, /* 2464 */
128'hfd469501a83046134787c62af57c0faf, /* 2465 */
128'h895cd7beffff5bb18b44f7af698098d8, /* 2466 */
128'h49b40821a679438efd9871936b901122, /* 2467 */
128'he9b6c7aa265e5a51c040b340f61e2562, /* 2468 */
128'he7d3fbc8d8a1e68102441453d62f105d, /* 2469 */
128'h455a14edf4d50d87c33707d621e1cde6, /* 2470 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /* 2471 */
128'hfde5380c6d9d61228771f681fffa3942, /* 2472 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /* 2473 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /* 2474 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /* 2475 */
128'hfc93a039ab9423a7432aff97f4292244, /* 2476 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /* 2477 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /* 2478 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /* 2479 */
128'h0c07020d08030e09040f0a05000b0601, /* 2480 */
128'h020f0c090603000d0a0704010e0b0805, /* 2481 */
128'h09020b040d060f08010a030c050e0700, /* 2482 */
128'h6c5f7465735f64735f63736972776f6c, /* 2483 */
128'h6e67696c615f64730000000000006465, /* 2484 */
128'h645f6b6c635f64730000000000000000, /* 2485 */
128'h69747465735f64730000000000007669, /* 2486 */
128'h735f646d635f6473000000000000676e, /* 2487 */
128'h74657365725f64730000000074726174, /* 2488 */
128'h6e636b6c625f64730000000000000000, /* 2489 */
128'h69736b6c625f64730000000000000074, /* 2490 */
128'h6f656d69745f6473000000000000657a, /* 2491 */
128'h655f7172695f64730000000000007475, /* 2492 */
128'h5f63736972776f6c000000000000006e, /* 2493 */
128'h00000000646d635f74726174735f6473, /* 2494 */
128'h746e695f746961775f63736972776f6c, /* 2495 */
128'h000000000067616c665f747075727265, /* 2496 */
128'h00007172695f64735f63736972776f6c, /* 2497 */
128'h695f646d635f64735f63736972776f6c, /* 2498 */
128'h5f63736972776f6c0000000000007172, /* 2499 */
128'h007172695f646e655f617461645f6473, /* 2500 */
128'h0000000087fe9c880000000087feaf50, /* 2501 */
128'h004c4b40004c4b400030000020000000, /* 2502 */
128'h6d6d5f6472616f62000000020000ffff, /* 2503 */
128'h0000000087fe4e980064637465675f63, /* 2504 */
128'h0000000087fe4d040000000087fe4aa6, /* 2505 */
128'h00000000000000000000000000000000, /* 2506 */
128'hffffbb7affffbb76ffffbb76ffffbb50, /* 2507 */
128'hffffbb7effffbb7effffbb7effffbb7e, /* 2508 */
128'h0000000087feb2780000000087feb268, /* 2509 */
128'h0000000087feb2a00000000087feb288, /* 2510 */
128'h0000000087feb2d00000000087feb2b8, /* 2511 */
128'h0000000087feb3000000000087feb2e8, /* 2512 */
128'h0000000087feb3300000000087feb318, /* 2513 */
128'h0000000087feb3600000000087feb348, /* 2514 */
128'h40040300400402004004010040040000, /* 2515 */
128'h40050000400405004004040140040400, /* 2516 */
128'h30000000000000030000000040050100, /* 2517 */
128'h60000000000000053000000000000001, /* 2518 */
128'h70000000000000027000000000000004, /* 2519 */
128'h00000001400000007000000000000000, /* 2520 */
128'h00000005000000012000000000000006, /* 2521 */
128'h20000000000000020000000040000000, /* 2522 */
128'h00000000100000000000000100000000, /* 2523 */
128'h1e19140f0d0c0a000000000000000000, /* 2524 */
128'h000186a00000271050463c37322d2823, /* 2525 */
128'h017d7840017d784000989680000f4240, /* 2526 */
128'h031975000319750002faf080018cba80, /* 2527 */
128'h02faf08005f5e10002faf080017d7840, /* 2528 */
128'h00000020000000000bebc2000c65d400, /* 2529 */
128'h00000200000001000000008000000040, /* 2530 */
128'h00002000000010000000080000000400, /* 2531 */
128'h0000c000000080000000600000004000, /* 2532 */
128'h37363534333231300002000000010000, /* 2533 */
128'h2043534952776f4c4645444342413938, /* 2534 */
128'h746f6f622d7520646573696d696e696d, /* 2535 */
128'h00000000647261432d445320726f6620, /* 2536 */
128'hfffff9d0fffff9e6fffff9d2fffff9be, /* 2537 */
128'h00000000fffffa0afffff9d0fffff9f8, /* 2538 */
128'he00600003800000039080000edfe0dd0, /* 2539 */
128'h00000000100000001100000028000000, /* 2540 */
128'h0000000000000000a806000059010000, /* 2541 */
128'h00000000010000000000000000000000, /* 2542 */
128'h02000000000000000400000003000000, /* 2543 */
128'h020000000f0000000400000003000000, /* 2544 */
128'h2c6874651b0000001400000003000000, /* 2545 */
128'h007665642d657261622d656e61697261, /* 2546 */
128'h2c687465260000001000000003000000, /* 2547 */
128'h0100000000657261622d656e61697261, /* 2548 */
128'h1a0000000300000000006e65736f6863, /* 2549 */
128'h303140747261752f636f732f2c000000, /* 2550 */
128'h0000003030323531313a303030303030, /* 2551 */
128'h00000000737570630100000002000000, /* 2552 */
128'h01000000000000000400000003000000, /* 2553 */
128'h000000000f0000000400000003000000, /* 2554 */
128'h40787d01380000000400000003000000, /* 2555 */
128'h03000000000000304075706301000000, /* 2556 */
128'h0300000080f0fa024b00000004000000, /* 2557 */
128'h03000000007570635b00000004000000, /* 2558 */
128'h03000000000000006700000004000000, /* 2559 */
128'h0000000079616b6f6b00000005000000, /* 2560 */
128'h7a6874651b0000001300000003000000, /* 2561 */
128'h0000766373697200656e61697261202c, /* 2562 */
128'h34367672720000000b00000003000000, /* 2563 */
128'h0b000000030000000000636466616d69, /* 2564 */
128'h0000393376732c76637369727c000000, /* 2565 */
128'h01000000850000000000000003000000, /* 2566 */
128'h6f72746e6f632d747075727265746e69, /* 2567 */
128'h04000000030000000000000072656c6c, /* 2568 */
128'h0000000003000000010000008f000000, /* 2569 */
128'h1b0000000f00000003000000a0000000, /* 2570 */
128'h000063746e692d7570632c7663736972, /* 2571 */
128'h01000000b50000000400000003000000, /* 2572 */
128'h01000000bb0000000400000003000000, /* 2573 */
128'h01000000020000000200000002000000, /* 2574 */
128'h0030303030303030384079726f6d656d, /* 2575 */
128'h6f6d656d5b0000000700000003000000, /* 2576 */
128'h67000000100000000300000000007972, /* 2577 */
128'h00000008000000000000008000000000, /* 2578 */
128'h0300000000636f730100000002000000, /* 2579 */
128'h03000000020000000000000004000000, /* 2580 */
128'h03000000020000000f00000004000000, /* 2581 */
128'h616972612c6874651b0000001f000000, /* 2582 */
128'h706d697300636f732d657261622d656e, /* 2583 */
128'h000000000300000000007375622d656c, /* 2584 */
128'h303240746e696c6301000000c3000000, /* 2585 */
128'h0d000000030000000000003030303030, /* 2586 */
128'h30746e696c632c76637369721b000000, /* 2587 */
128'hca000000100000000300000000000000, /* 2588 */
128'h07000000010000000300000001000000, /* 2589 */
128'h00000000670000001000000003000000, /* 2590 */
128'h0300000000000c000000000000000002, /* 2591 */
128'h006c6f72746e6f63de00000008000000, /* 2592 */
128'h7075727265746e690100000002000000, /* 2593 */
128'h3030634072656c6c6f72746e6f632d74, /* 2594 */
128'h04000000030000000000000030303030, /* 2595 */
128'h04000000030000000000000000000000, /* 2596 */
128'h0c00000003000000010000008f000000, /* 2597 */
128'h003063696c702c76637369721b000000, /* 2598 */
128'h03000000a00000000000000003000000, /* 2599 */
128'h0b00000001000000ca00000010000000, /* 2600 */
128'h10000000030000000900000001000000, /* 2601 */
128'h000000000000000c0000000067000000, /* 2602 */
128'he8000000040000000300000000000004, /* 2603 */
128'hfb000000040000000300000007000000, /* 2604 */
128'hb5000000040000000300000003000000, /* 2605 */
128'hbb000000040000000300000002000000, /* 2606 */
128'h75626564010000000200000002000000, /* 2607 */
128'h0000304072656c6c6f72746e6f632d67, /* 2608 */
128'h637369721b0000001000000003000000, /* 2609 */
128'h03000000003331302d67756265642c76, /* 2610 */
128'hffff000001000000ca00000008000000, /* 2611 */
128'h00000000670000001000000003000000, /* 2612 */
128'h03000000001000000000000000000000, /* 2613 */
128'h006c6f72746e6f63de00000008000000, /* 2614 */
128'h30303140747261750100000002000000, /* 2615 */
128'h08000000030000000000003030303030, /* 2616 */
128'h03000000003035373631736e1b000000, /* 2617 */
128'h00000010000000006700000010000000, /* 2618 */
128'h04000000030000000010000000000000, /* 2619 */
128'h040000000300000080f0fa024b000000, /* 2620 */
128'h040000000300000000c2010006010000, /* 2621 */
128'h04000000030000000200000014010000, /* 2622 */
128'h04000000030000000100000025010000, /* 2623 */
128'h04000000030000000200000030010000, /* 2624 */
128'h0100000002000000040000003a010000, /* 2625 */
128'h3030303240636d6d2d63736972776f6c, /* 2626 */
128'h10000000030000000000000030303030, /* 2627 */
128'h00000000000000200000000067000000, /* 2628 */
128'h14010000040000000300000000000100, /* 2629 */
128'h25010000040000000300000002000000, /* 2630 */
128'h1b0000000c0000000300000002000000, /* 2631 */
128'h0200000000636d6d2d63736972776f6c, /* 2632 */
128'h406874652d63736972776f6c01000000, /* 2633 */
128'h03000000000000003030303030303033, /* 2634 */
128'h2d63736972776f6c1b0000000c000000, /* 2635 */
128'h5b000000080000000300000000687465, /* 2636 */
128'h0400000003000000006b726f7774656e, /* 2637 */
128'h04000000030000000200000014010000, /* 2638 */
128'h06000000030000000300000025010000, /* 2639 */
128'h0300000000007fe3023e180047010000, /* 2640 */
128'h00000030000000006700000010000000, /* 2641 */
128'h01000000020000000080000000000000, /* 2642 */
128'h303440646e7277682d63736972776f6c, /* 2643 */
128'h0e000000030000000000303030303030, /* 2644 */
128'h6e7277682d63736972776f6c1b000000, /* 2645 */
128'h67000000100000000300000000000064, /* 2646 */
128'h00100000000000000000004000000000, /* 2647 */
128'h09000000020000000200000002000000, /* 2648 */
128'h2300736c6c65632d7373657264646123, /* 2649 */
128'h61706d6f6300736c6c65632d657a6973, /* 2650 */
128'h6f647473006c65646f6d00656c626974, /* 2651 */
128'h65736162656d697400687461702d7475, /* 2652 */
128'h6b636f6c630079636e6575716572662d, /* 2653 */
128'h63697665640079636e6575716572662d, /* 2654 */
128'h75746174730067657200657079745f65, /* 2655 */
128'h2d756d6d006173692c76637369720073, /* 2656 */
128'h230074696c70732d626c740065707974, /* 2657 */
128'h00736c6c65632d747075727265746e69, /* 2658 */
128'h6f72746e6f632d747075727265746e69, /* 2659 */
128'h646e6168702c78756e696c0072656c6c, /* 2660 */
128'h727265746e69007365676e617200656c, /* 2661 */
128'h6572006465646e657478652d73747075, /* 2662 */
128'h616d2c76637369720073656d616e2d67, /* 2663 */
128'h766373697200797469726f6972702d78, /* 2664 */
128'h70732d746e6572727563007665646e2c, /* 2665 */
128'h61702d747075727265746e6900646565, /* 2666 */
128'h0073747075727265746e6900746e6572, /* 2667 */
128'h6f692d6765720074666968732d676572, /* 2668 */
128'h63616d2d6c61636f6c0068746469772d, /* 2669 */
128'h0000000000000000737365726464612d, /* 2670 */
128'h0000000000203a642520656369766544, /* 2671 */
128'h00203a6425206563697665642073250a, /* 2672 */
128'h00000000203a6425206563697665440a, /* 2673 */
128'h000a656369766564206e776f6e6b6e75, /* 2674 */
128'h00000a2973252c73252870756b6f6f6c, /* 2675 */
128'h7265206c616e7265746e692070636864, /* 2676 */
128'h00000000000000000a7025202c726f72, /* 2677 */
128'h5145525f5043484420676e69646e6553, /* 2678 */
128'h4b434120504348440000000a54534555, /* 2679 */
128'h696c432050434844000000000000000a, /* 2680 */
128'h203a7373657264644120504920746e65, /* 2681 */
128'h0000000a64252e64252e64252e642520, /* 2682 */
128'h73657264644120504920726576726553, /* 2683 */
128'h0a64252e64252e64252e642520203a73, /* 2684 */
128'h6120726574756f520000000000000000, /* 2685 */
128'h252e64252e642520203a737365726464, /* 2686 */
128'h6b73616d2074654e0000000a64252e64, /* 2687 */
128'h64252e642520203a7373657264646120, /* 2688 */
128'h697420657361654c000a64252e64252e, /* 2689 */
128'h7364253a6d64253a686425203d20656d, /* 2690 */
128'h3d206e69616d6f44000000000000000a, /* 2691 */
128'h4820746e65696c4300000a2273252220, /* 2692 */
128'h000a22732522203d20656d616e74736f, /* 2693 */
128'h000000000a44455050494b53204b4341, /* 2694 */
128'h000000000000000a4b414e2050434844, /* 2695 */
128'h73657264646120646574736575716552, /* 2696 */
128'h0000000000000a646573756665722073, /* 2697 */
128'h000000000000000a732520726f727245, /* 2698 */
128'h6e6f6974706f2064656c646e61686e75, /* 2699 */
128'h656c646e61686e55000000000a642520, /* 2700 */
128'h64252065646f63706f20504348442064, /* 2701 */
128'h20676e69646e6553000000000000000a, /* 2702 */
128'h000a595245564f435349445f50434844, /* 2703 */
128'h00000000000a29732528726f72726570, /* 2704 */
128'h3a2043414d2073250000000030687465, /* 2705 */
128'h3a583230253a583230253a5832302520, /* 2706 */
128'h000a583230253a583230253a58323025, /* 2707 */
128'h484420646e65732074276e646c756f43, /* 2708 */
128'h206e6f20595245564f43534944205043, /* 2709 */
128'h00000a7325203a732520656369766564, /* 2710 */
128'h5043484420726f6620676e6974696157, /* 2711 */
128'h2020202020202020000a524546464f5f, /* 2712 */
128'h00000000000063250000000000000020, /* 2713 */
128'h0000005832302520000000000000002e, /* 2714 */
128'h00000000732573250000000000000a0a, /* 2715 */
128'h00000000007325203a646c697542202c, /* 2716 */
128'h73257a4820756c250000000000007325, /* 2717 */
128'h0000000000756c250000000000000000, /* 2718 */
128'h0073257a4863252000000000646c252e, /* 2719 */
128'h00000000007325736574794220756c25, /* 2720 */
128'h00003a786c3830250073254269632520, /* 2721 */
128'h000a73252020202000786c6c2a302520, /* 2722 */
128'h000000203a5d64255b6e6f6974636553, /* 2723 */
128'h727265207974696e6173207264646170, /* 2724 */
128'h2c7825286e666c6500000a702520726f, /* 2725 */
128'h000000000a3b29782578302c78257830, /* 2726 */
128'h782578302c302c7825287465736d656d, /* 2727 */
128'h464f5f4f4c43414d00000000000a3b29, /* 2728 */
128'h464f5f494843414d0000000054455346, /* 2729 */
128'h46464f5f524c50540000000054455346, /* 2730 */
128'h46464f5f534346540000000000544553, /* 2731 */
128'h4c5254434f49444d0000000000544553, /* 2732 */
128'h46464f5f534346520054455346464f5f, /* 2733 */
128'h5346464f5f5253520000000000544553, /* 2734 */
128'h46464f5f444142520000000000005445, /* 2735 */
128'h46464f5f524c50520000000000544553, /* 2736 */
128'h000000003f3f3f3f0000000000544553, /* 2737 */
128'h000064252b54455346464f5f524c5052, /* 2738 */
128'h6f746f72502050490000000000000047, /* 2739 */
128'h00000000000000000a50495049203d20, /* 2740 */
128'h6f746f72502050490000000000000054, /* 2741 */
128'h6f746f7250205049000a504745203d20, /* 2742 */
128'h6165682074736574000a505550203d20, /* 2743 */
128'h6e6f6320747365740000000a3a726564, /* 2744 */
128'h6f746f7250205049000a3a73746e6574, /* 2745 */
128'h6f746f7250205049000a504449203d20, /* 2746 */
128'h6f746f725020504900000a5054203d20, /* 2747 */
128'h00000000000000000a50434344203d20, /* 2748 */
128'h6f746f72502050490000000000000036, /* 2749 */
128'h00000000000000000a50565352203d20, /* 2750 */
128'h000a455247203d206f746f7250205049, /* 2751 */
128'h000a505345203d206f746f7250205049, /* 2752 */
128'h00000a4841203d206f746f7250205049, /* 2753 */
128'h000a50544d203d206f746f7250205049, /* 2754 */
128'h5054454542203d206f746f7250205049, /* 2755 */
128'h6f746f72502050490000000000000a48, /* 2756 */
128'h000000000000000a5041434e45203d20, /* 2757 */
128'h6f746f7250205049000000000000004d, /* 2758 */
128'h00000000000000000a504d4f43203d20, /* 2759 */
128'h0a50544353203d206f746f7250205049, /* 2760 */
128'h6f746f72502050490000000000000000, /* 2761 */
128'h00000000000a4554494c504455203d20, /* 2762 */
128'h0a534c504d203d206f746f7250205049, /* 2763 */
128'h6f746f72502050490000000000000000, /* 2764 */
128'h6f746f7270205049000a574152203d20, /* 2765 */
128'h2820646574726f707075736e75203d20, /* 2766 */
128'h79745f6f746f7270000000000a297825, /* 2767 */
128'h0000000000000a78257830203d206570, /* 2768 */
128'h727265746e692064656c646e61686e75, /* 2769 */
128'h414d2070757465530000000a21747075, /* 2770 */
128'h4d454f2049505351000a726464612043, /* 2771 */
128'h0000000000000a7825203d205d64255b, /* 2772 */
128'h00000a786c253a786c25203d2043414d, /* 2773 */
128'h3025203d20737365726464612043414d, /* 2774 */
128'h3230253a783230253a783230253a7832, /* 2775 */
128'h0000000a2e783230253a783230253a78, /* 2776 */
128'h00007f7c5d5b3f3e3d3c3b3a2c2b2a22, /* 2777 */
128'h007f7c5d5b3f3e3d3c3b3a2e2c2b2a22, /* 2778 */
128'h66656463626139383736353433323130, /* 2779 */
128'h72776f6c2f6372730000000000000000, /* 2780 */
128'h00000000000000632e636d6d5f637369, /* 2781 */
128'h61625f6473203d3d20657361625f6473, /* 2782 */
128'h5f63736972776f6c00726464615f6573, /* 2783 */
128'h000a74756f656d6974207325203a6473, /* 2784 */
128'h616d202c6465766f6d65722064726143, /* 2785 */
128'h6425206f74206465676e616863206b73, /* 2786 */
128'h736e692064726143000000000000000a, /* 2787 */
128'h6e616863206b73616d202c6465747265, /* 2788 */
128'h0000000000000a6425206f7420646567, /* 2789 */
128'h25207461206465746165726320636d6d, /* 2790 */
128'h0000000a7825203d2074736f68202c78, /* 2791 */
128'h0000000000006f4e0000000000736559, /* 2792 */
128'h002020203a434d4d0000000052444420, /* 2793 */
128'h00000000000a7325203a656369766544, /* 2794 */
128'h3a4449207265727574636166756e614d, /* 2795 */
128'h0a7825203a4d454f000000000a782520, /* 2796 */
128'h6325203a656d614e0000000000000000, /* 2797 */
128'h0000000000000a206325632563256325, /* 2798 */
128'h00000a6425203a646565705320737542, /* 2799 */
128'h25203a79746963617061432068676948, /* 2800 */
128'h79746963617061430000000000000a73, /* 2801 */
128'h7464695720737542000000000000203a, /* 2802 */
128'h000000000a73257469622d6425203a68, /* 2803 */
128'h0000007825782520000000203a78250a, /* 2804 */
128'h00000000000064735f63736972776f6c, /* 2805 */
128'h0000000065646f6d206e776f6e6b6e55, /* 2806 */
128'h7830203a726f72724520737574617453, /* 2807 */
128'h2074756f656d69540000000a58383025, /* 2808 */
128'h616572206472616320676e6974696177, /* 2809 */
128'h6c69616620636d6d00000000000a7964, /* 2810 */
128'h6d6320706f747320646e6573206f7420, /* 2811 */
128'h6f6c62203a434d4d0000000000000a64, /* 2812 */
128'h20786c257830207265626d756e206b63, /* 2813 */
128'h6c2578302878616d2073646565637865, /* 2814 */
128'h203d3e20434d4d6500000000000a2978, /* 2815 */
128'h726f6620646572697571657220342e34, /* 2816 */
128'h642072657375206465636e61686e6520, /* 2817 */
128'h000000000000000a6165726120617461, /* 2818 */
128'h757320746f6e2073656f642064726143, /* 2819 */
128'h696e6f697469747261702074726f7070, /* 2820 */
128'h656f64206472614300000000000a676e, /* 2821 */
128'h20434820656e6966656420746f6e2073, /* 2822 */
128'h00000a657a69732070756f7267205057, /* 2823 */
128'h636e61686e6520617461642072657355, /* 2824 */
128'h5720434820746f6e2061657261206465, /* 2825 */
128'h696c6120657a69732070756f72672050, /* 2826 */
128'h72617020692550470000000a64656e67, /* 2827 */
128'h505720434820746f6e206e6f69746974, /* 2828 */
128'h67696c6120657a69732070756f726720, /* 2829 */
128'h656f642064726143000000000a64656e, /* 2830 */
128'h6e652074726f7070757320746f6e2073, /* 2831 */
128'h657475626972747461206465636e6168, /* 2832 */
128'h6e65206c61746f54000000000000000a, /* 2833 */
128'h6563786520657a6973206465636e6168, /* 2834 */
128'h20752528206d756d6978616d20736465, /* 2835 */
128'h656f64206472614300000a297525203e, /* 2836 */
128'h6f682074726f7070757320746f6e2073, /* 2837 */
128'h61702064656c6c6f72746e6f63207473, /* 2838 */
128'h6572206574697277206e6f6974697472, /* 2839 */
128'h6e6974746573207974696c696261696c, /* 2840 */
128'h726c61206472614300000000000a7367, /* 2841 */
128'h64656e6f697469747261702079646165, /* 2842 */
128'h206f6e203a434d4d000000000000000a, /* 2843 */
128'h0000000a746e65736572702064726163, /* 2844 */
128'h73657220746f6e206469642064726143, /* 2845 */
128'h20656761746c6f76206f7420646e6f70, /* 2846 */
128'h00000000000000000a217463656c6573, /* 2847 */
128'h7463656c6573206f7420656c62616e75, /* 2848 */
128'h00000000000000000a65646f6d206120, /* 2849 */
128'h646e756f66206473635f747865206f4e, /* 2850 */
128'h78363025206e614d0000000000000a21, /* 2851 */
128'h000000783430257834302520726e5320, /* 2852 */
128'h00000000632563256325632563256325, /* 2853 */
128'h6167656c20434d4d00000064252e6425, /* 2854 */
128'h636167654c2044530000000000007963, /* 2855 */
128'h6867694820434d4d0000000000000079, /* 2856 */
128'h0000297a484d36322820646565705320, /* 2857 */
128'h35282064656570532068676948204453, /* 2858 */
128'h6867694820434d4d000000297a484d30, /* 2859 */
128'h0000297a484d32352820646565705320, /* 2860 */
128'h7a484d32352820323552444420434d4d, /* 2861 */
128'h31524453205348550000000000000029, /* 2862 */
128'h00000000000000297a484d3532282032, /* 2863 */
128'h7a484d30352820353252445320534855, /* 2864 */
128'h35524453205348550000000000000029, /* 2865 */
128'h000000000000297a484d303031282030, /* 2866 */
128'h7a484d30352820303552444420534855, /* 2867 */
128'h31524453205348550000000000000029, /* 2868 */
128'h0000000000297a484d38303228203430, /* 2869 */
128'h0000297a484d30303228203030325348, /* 2870 */
128'h6f6e2064252065636976654420434d4d, /* 2871 */
128'h00000000000000000a646e756f662074, /* 2872 */
128'h000000000000445300000000434d4d65, /* 2873 */
128'h000000297325282000006425203a7325, /* 2874 */
128'h6e656c20656c69460000000000636d6d, /* 2875 */
128'h000000000000000a6425203d20687467, /* 2876 */
128'h0a7325203d202964252c70252835646d, /* 2877 */
128'h666c652064616f6c0000000000000000, /* 2878 */
128'h000a79726f6d656d20524444206f7420, /* 2879 */
128'h2064656c696166206461657220666c65, /* 2880 */
128'h000000646c252065646f632068746977, /* 2881 */
128'h6f6f7420687461702074736575716552, /* 2882 */
128'h00000000000a646c25202e676e6f6c20, /* 2883 */
128'h732522203a717277000000000000002f, /* 2884 */
128'h0a64253d657a69736b636f6c62202c22, /* 2885 */
128'h20657669656365520000000000000000, /* 2886 */
128'h0000000000000a2e646e6520656c6966, /* 2887 */
128'h656c6c6163207172775f656c646e6168, /* 2888 */
128'h206c6167656c6c4900000000000a2e64, /* 2889 */
128'h0a2e6e6f6974617265706f2050544654, /* 2890 */
128'h75716572206e656c0000000000000000, /* 2891 */
128'h6175746361202c5825203d2064657269, /* 2892 */
128'h000000005c2d2f7c000a7825203d206c, /* 2893 */
128'h20646564616f6c2065687420746f6f42, /* 2894 */
128'h6572646461207461206d6172676f7270, /* 2895 */
128'h000000000000000a2e2e2e7025207373, /* 2896 */
128'h445320746e756f6d206f74206c696146, /* 2897 */
128'h000000000000000a2172657669726420, /* 2898 */
128'h6e69206e69622e746f6f622064616f4c, /* 2899 */
128'h0000000000000a79726f6d656d206f74, /* 2900 */
128'h00000000000000006e69622e746f6f62, /* 2901 */
128'h62206e65706f206f742064656c696146, /* 2902 */
128'h206f74206c6961660000000a21746f6f, /* 2903 */
128'h000000000021656c69662065736f6c63, /* 2904 */
128'h6420746e756f6d75206f74206c696166, /* 2905 */
128'h20746f6f622d750a00000000216b7369, /* 2906 */
128'h67617473207473726966206465736162, /* 2907 */
128'h00000a726564616f6c20746f6f622065, /* 2908 */
128'h696166207325206e6f69747265737361, /* 2909 */
128'h696c202c732520656c6966202c64656c, /* 2910 */
128'h206e6f6974636e7566202c642520656e, /* 2911 */
128'h3a4552554c49414600000000000a7325, /* 2912 */
128'h74612078257830203d21207825783020, /* 2913 */
128'h00000a2e782578302074657366666f20, /* 2914 */
128'h7025203d203270202c7025203d203170, /* 2915 */
128'h2020202020202020000000000000000a, /* 2916 */
128'h08080808080808080000000000202020, /* 2917 */
128'h20676e69747465730000000000080808, /* 2918 */
128'h20676e69747365740000000000007525, /* 2919 */
128'h3a4552554c4941460000000000007525, /* 2920 */
128'h64612064616220656c626973736f7020, /* 2921 */
128'h666f20746120656e696c207373657264, /* 2922 */
128'h00000000000a2e782578302074657366, /* 2923 */
128'h7478656e206f7420676e697070696b53, /* 2924 */
128'h000000000000000a2e2e2e7473657420, /* 2925 */
128'h20202020200808080808080808080808, /* 2926 */
128'h08080808080808080808202020202020, /* 2927 */
128'h00000000000820080000000000000008, /* 2928 */
128'h78302073692065676e61722074736574, /* 2929 */
128'h00000000000a70257830206f74207025, /* 2930 */
128'h000000000075252f00752520706f6f4c, /* 2931 */
128'h6441206b637574530000000000000a3a, /* 2932 */
128'h0000203a732520200000007373657264, /* 2933 */
128'h00000a2e656e6f4400000000000a6b6f, /* 2934 */
128'h4d415244206c6174656d20657261420a, /* 2935 */
128'h65747365746d656d00000a7473657420, /* 2936 */
128'h20302e332e34206e6f69737265762072, /* 2937 */
128'h000000000000000a297469622d642528, /* 2938 */
128'h30322029432820746867697279706f43, /* 2939 */
128'h2073656c7261684320323130322d3130, /* 2940 */
128'h000000000000000a2e6e6f62617a6143, /* 2941 */
128'h74207265646e75206465736e6563694c, /* 2942 */
128'h50206c6172656e654720554e47206568, /* 2943 */
128'h65762065736e6563694c2063696c6275, /* 2944 */
128'h0a2e29796c6e6f282032206e6f697372, /* 2945 */
128'h5f676e696b726f770000000000000000, /* 2946 */
128'h20646c25202c424b6425203d20746573, /* 2947 */
128'h6c25202c736e6f697463757274736e69, /* 2948 */
128'h203d20495043202c73656c6379632064, /* 2949 */
128'h00000000000000000a646c252e646c25, /* 2950 */
128'h46454443424139383736353433323130, /* 2951 */
128'h6f57206f6c6c65480000000000000000, /* 2952 */
128'h205d64255b70777300000a0d21646c72, /* 2953 */
128'h73206863746977530000000a5825203d, /* 2954 */
128'h000a58252c5825203d20676e69747465, /* 2955 */
128'h5825203d2064656573206d6f646e6152, /* 2956 */
128'h0a746f6f62204453000000000000000a, /* 2957 */
128'h6f6f6220495053510000000000000000, /* 2958 */
128'h736574204d4152440000000000000a74, /* 2959 */
128'h6f6f6220505446540000000000000a74, /* 2960 */
128'h65742065686361430000000000000a74, /* 2961 */
128'h00000a0d7061727400000000000a7473, /* 2962 */
128'h00000002464c457fcccccccccccccccd, /* 2963 */
128'h1032547698badcfeefcdab8967452301, /* 2964 */
128'h5851f42d4c957f2d1000000020000000, /* 2965 */
128'haaaaaaaaaaaaaaaa5555555555555555, /* 2966 */
128'h00000000000000000000000000000000, /* 2967 */
128'h00000000000000000000000000000000, /* 2968 */
128'h00000000000000000000000000000000, /* 2969 */
128'h00000000000000000000000000000000, /* 2970 */
128'h00000000000000000000000000000000, /* 2971 */
128'h00000000000000000000000000000000, /* 2972 */
128'h00000000000000000000000000000000, /* 2973 */
128'h00000000000000000000000000000000, /* 2974 */
128'h00000000000000000000000000000000, /* 2975 */
128'h00004b4d47545045000000030f060301, /* 2976 */
128'h000000003000000000000000004b4d47, /* 2977 */
128'h00000000ffffffff0000000000000000, /* 2978 */
128'h0000646d635f6473000000000c000000, /* 2979 */
128'h00000000ffffffff00006772615f6473, /* 2980 */
128'h000000002f7c5c2d0000000087feb1f8, /* 2981 */
128'h000000060000000087feb3b0cc33aa55, /* 2982 */
128'h87fe70900000000000000000ffffffff, /* 2983 */
128'h00000000000000000000000000000000, /* 2984 */
128'h00000000000000000000000000000000, /* 2985 */
128'h00000000000000000000000000000000, /* 2986 */
128'h00000000000000000000000000000000, /* 2987 */
128'h00000000000000000000000000000000, /* 2988 */
128'h00000000000000000000000000000000, /* 2989 */
128'h00000000000000000000000000000000, /* 2990 */
128'h00000000000000000000000000000000, /* 2991 */
128'h00000000000000000000000000000000, /* 2992 */
128'h00000000000000000000000000000000, /* 2993 */
128'h00000000000000000000000000000000, /* 2994 */
128'h00000000000000000000000000000000, /* 2995 */
128'h00000000000000000000000000000000, /* 2996 */
128'h00000000000000000000000000000000, /* 2997 */
128'h00000000000000000000000000000000, /* 2998 */
128'h00000000000000000000000000000000, /* 2999 */
128'h00000000000000000000000000000000, /* 3000 */
128'h00000000000000000000000000000000, /* 3001 */
128'h00000000000000000000000000000000, /* 3002 */
128'h00000000000000000000000000000000, /* 3003 */
128'h00000000000000000000000000000000, /* 3004 */
128'h00000000000000000000000000000000, /* 3005 */
128'h00000000000000000000000000000000, /* 3006 */
128'h00000000000000000000000000000000, /* 3007 */
128'h00000000000000000000000000000000, /* 3008 */
128'h00000000000000000000000000000000, /* 3009 */
128'h00000000000000000000000000000000, /* 3010 */
128'h00000000000000000000000000000000, /* 3011 */
128'h00000000000000000000000000000000, /* 3012 */
128'h00000000000000000000000000000000, /* 3013 */
128'h00000000000000000000000000000000, /* 3014 */
128'h00000000000000000000000000000000, /* 3015 */
128'h00000000000000000000000000000000, /* 3016 */
128'h00000000000000000000000000000000, /* 3017 */
128'h00000000000000000000000000000000, /* 3018 */
128'h00000000000000000000000000000000, /* 3019 */
128'h00000000000000000000000000000000, /* 3020 */
128'h00000000000000000000000000000000, /* 3021 */
128'h00000000000000000000000000000000, /* 3022 */
128'h00000000000000000000000000000000, /* 3023 */
128'h00000000000000000000000000000000, /* 3024 */
128'h00000000000000000000000000000000, /* 3025 */
128'h00000000000000000000000000000000, /* 3026 */
128'h00000000000000000000000000000000, /* 3027 */
128'h00000000000000000000000000000000, /* 3028 */
128'h00000000000000000000000000000000, /* 3029 */
128'h00000000000000000000000000000000, /* 3030 */
128'h00000000000000000000000000000000, /* 3031 */
128'h00000000000000000000000000000000, /* 3032 */
128'h00000000000000000000000000000000, /* 3033 */
128'h00000000000000000000000000000000, /* 3034 */
128'h00000000000000000000000000000000, /* 3035 */
128'h00000000000000000000000000000000, /* 3036 */
128'h00000000000000000000000000000000, /* 3037 */
128'h00000000000000000000000000000000, /* 3038 */
128'h00000000000000000000000000000000, /* 3039 */
128'h00000000000000000000000000000000, /* 3040 */
128'h00000000000000000000000000000000, /* 3041 */
128'h00000000000000000000000000000000, /* 3042 */
128'h00000000000000000000000000000000, /* 3043 */
128'h00000000000000000000000000000000, /* 3044 */
128'h00000000000000000000000000000000, /* 3045 */
128'h00000000000000000000000000000000, /* 3046 */
128'h00000000000000000000000000000000, /* 3047 */
128'h00000000000000000000000000000000, /* 3048 */
128'h00000000000000000000000000000000, /* 3049 */
128'h00000000000000000000000000000000, /* 3050 */
128'h00000000000000000000000000000000, /* 3051 */
128'h00000000000000000000000000000000, /* 3052 */
128'h00000000000000000000000000000000, /* 3053 */
128'h00000000000000000000000000000000, /* 3054 */
128'h00000000000000000000000000000000, /* 3055 */
128'h00000000000000000000000000000000, /* 3056 */
128'h00000000000000000000000000000000, /* 3057 */
128'h00000000000000000000000000000000, /* 3058 */
128'h00000000000000000000000000000000, /* 3059 */
128'h00000000000000000000000000000000, /* 3060 */
128'h00000000000000000000000000000000, /* 3061 */
128'h00000000000000000000000000000000, /* 3062 */
128'h00000000000000000000000000000000, /* 3063 */
128'h00000000000000000000000000000000, /* 3064 */
128'h00000000000000000000000000000000, /* 3065 */
128'h00000000000000000000000000000000, /* 3066 */
128'h00000000000000000000000000000000, /* 3067 */
128'h00000000000000000000000000000000, /* 3068 */
128'h00000000000000000000000000000000, /* 3069 */
128'h00000000000000000000000000000000, /* 3070 */
128'h00000000000000000000000000000000, /* 3071 */
128'h00000000000000000000000000000000, /* 3072 */
128'h00000000000000000000000000000000, /* 3073 */
128'h00000000000000000000000000000000, /* 3074 */
128'h00000000000000000000000000000000, /* 3075 */
128'h00000000000000000000000000000000, /* 3076 */
128'h00000000000000000000000000000000, /* 3077 */
128'h00000000000000000000000000000000, /* 3078 */
128'h00000000000000000000000000000000, /* 3079 */
128'h00000000000000000000000000000000, /* 3080 */
128'h00000000000000000000000000000000, /* 3081 */
128'h00000000000000000000000000000000, /* 3082 */
128'h00000000000000000000000000000000, /* 3083 */
128'h00000000000000000000000000000000, /* 3084 */
128'h00000000000000000000000000000000, /* 3085 */
128'h00000000000000000000000000000000, /* 3086 */
128'h00000000000000000000000000000000, /* 3087 */
128'h00000000000000000000000000000000, /* 3088 */
128'h00000000000000000000000000000000, /* 3089 */
128'h00000000000000000000000000000000, /* 3090 */
128'h00000000000000000000000000000000, /* 3091 */
128'h00000000000000000000000000000000, /* 3092 */
128'h00000000000000000000000000000000, /* 3093 */
128'h00000000000000000000000000000000, /* 3094 */
128'h00000000000000000000000000000000, /* 3095 */
128'h00000000000000000000000000000000, /* 3096 */
128'h00000000000000000000000000000000, /* 3097 */
128'h00000000000000000000000000000000, /* 3098 */
128'h00000000000000000000000000000000, /* 3099 */
128'h00000000000000000000000000000000, /* 3100 */
128'h00000000000000000000000000000000, /* 3101 */
128'h00000000000000000000000000000000, /* 3102 */
128'h00000000000000000000000000000000, /* 3103 */
128'h00000000000000000000000000000000, /* 3104 */
128'h00000000000000000000000000000000, /* 3105 */
128'h00000000000000000000000000000000, /* 3106 */
128'h00000000000000000000000000000000, /* 3107 */
128'h00000000000000000000000000000000, /* 3108 */
128'h00000000000000000000000000000000, /* 3109 */
128'h00000000000000000000000000000000, /* 3110 */
128'h00000000000000000000000000000000, /* 3111 */
128'h00000000000000000000000000000000, /* 3112 */
128'h00000000000000000000000000000000, /* 3113 */
128'h00000000000000000000000000000000, /* 3114 */
128'h00000000000000000000000000000000, /* 3115 */
128'h00000000000000000000000000000000, /* 3116 */
128'h00000000000000000000000000000000, /* 3117 */
128'h00000000000000000000000000000000, /* 3118 */
128'h00000000000000000000000000000000, /* 3119 */
128'h00000000000000000000000000000000, /* 3120 */
128'h00000000000000000000000000000000, /* 3121 */
128'h00000000000000000000000000000000, /* 3122 */
128'h00000000000000000000000000000000, /* 3123 */
128'h00000000000000000000000000000000, /* 3124 */
128'h00000000000000000000000000000000, /* 3125 */
128'h00000000000000000000000000000000, /* 3126 */
128'h00000000000000000000000000000000, /* 3127 */
128'h00000000000000000000000000000000, /* 3128 */
128'h00000000000000000000000000000000, /* 3129 */
128'h00000000000000000000000000000000, /* 3130 */
128'h00000000000000000000000000000000, /* 3131 */
128'h00000000000000000000000000000000, /* 3132 */
128'h00000000000000000000000000000000, /* 3133 */
128'h00000000000000000000000000000000, /* 3134 */
128'h00000000000000000000000000000000, /* 3135 */
128'h00000000000000000000000000000000, /* 3136 */
128'h00000000000000000000000000000000, /* 3137 */
128'h00000000000000000000000000000000, /* 3138 */
128'h00000000000000000000000000000000, /* 3139 */
128'h00000000000000000000000000000000, /* 3140 */
128'h00000000000000000000000000000000, /* 3141 */
128'h00000000000000000000000000000000, /* 3142 */
128'h00000000000000000000000000000000, /* 3143 */
128'h00000000000000000000000000000000, /* 3144 */
128'h00000000000000000000000000000000, /* 3145 */
128'h00000000000000000000000000000000, /* 3146 */
128'h00000000000000000000000000000000, /* 3147 */
128'h00000000000000000000000000000000, /* 3148 */
128'h00000000000000000000000000000000, /* 3149 */
128'h00000000000000000000000000000000, /* 3150 */
128'h00000000000000000000000000000000, /* 3151 */
128'h00000000000000000000000000000000, /* 3152 */
128'h00000000000000000000000000000000, /* 3153 */
128'h00000000000000000000000000000000, /* 3154 */
128'h00000000000000000000000000000000, /* 3155 */
128'h00000000000000000000000000000000, /* 3156 */
128'h00000000000000000000000000000000, /* 3157 */
128'h00000000000000000000000000000000, /* 3158 */
128'h00000000000000000000000000000000, /* 3159 */
128'h00000000000000000000000000000000, /* 3160 */
128'h00000000000000000000000000000000, /* 3161 */
128'h00000000000000000000000000000000, /* 3162 */
128'h00000000000000000000000000000000, /* 3163 */
128'h00000000000000000000000000000000, /* 3164 */
128'h00000000000000000000000000000000, /* 3165 */
128'h00000000000000000000000000000000, /* 3166 */
128'h00000000000000000000000000000000, /* 3167 */
128'h00000000000000000000000000000000, /* 3168 */
128'h00000000000000000000000000000000, /* 3169 */
128'h00000000000000000000000000000000, /* 3170 */
128'h00000000000000000000000000000000, /* 3171 */
128'h00000000000000000000000000000000, /* 3172 */
128'h00000000000000000000000000000000, /* 3173 */
128'h00000000000000000000000000000000, /* 3174 */
128'h00000000000000000000000000000000, /* 3175 */
128'h00000000000000000000000000000000, /* 3176 */
128'h00000000000000000000000000000000, /* 3177 */
128'h00000000000000000000000000000000, /* 3178 */
128'h00000000000000000000000000000000, /* 3179 */
128'h00000000000000000000000000000000, /* 3180 */
128'h00000000000000000000000000000000, /* 3181 */
128'h00000000000000000000000000000000, /* 3182 */
128'h00000000000000000000000000000000, /* 3183 */
128'h00000000000000000000000000000000, /* 3184 */
128'h00000000000000000000000000000000, /* 3185 */
128'h00000000000000000000000000000000, /* 3186 */
128'h00000000000000000000000000000000, /* 3187 */
128'h00000000000000000000000000000000, /* 3188 */
128'h00000000000000000000000000000000, /* 3189 */
128'h00000000000000000000000000000000, /* 3190 */
128'h00000000000000000000000000000000, /* 3191 */
128'h00000000000000000000000000000000, /* 3192 */
128'h00000000000000000000000000000000, /* 3193 */
128'h00000000000000000000000000000000, /* 3194 */
128'h00000000000000000000000000000000, /* 3195 */
128'h00000000000000000000000000000000, /* 3196 */
128'h00000000000000000000000000000000, /* 3197 */
128'h00000000000000000000000000000000, /* 3198 */
128'h00000000000000000000000000000000, /* 3199 */
128'h00000000000000000000000000000000, /* 3200 */
128'h00000000000000000000000000000000, /* 3201 */
128'h00000000000000000000000000000000, /* 3202 */
128'h00000000000000000000000000000000, /* 3203 */
128'h00000000000000000000000000000000, /* 3204 */
128'h00000000000000000000000000000000, /* 3205 */
128'h00000000000000000000000000000000, /* 3206 */
128'h00000000000000000000000000000000, /* 3207 */
128'h00000000000000000000000000000000, /* 3208 */
128'h00000000000000000000000000000000, /* 3209 */
128'h00000000000000000000000000000000, /* 3210 */
128'h00000000000000000000000000000000, /* 3211 */
128'h00000000000000000000000000000000, /* 3212 */
128'h00000000000000000000000000000000, /* 3213 */
128'h00000000000000000000000000000000, /* 3214 */
128'h00000000000000000000000000000000, /* 3215 */
128'h00000000000000000000000000000000, /* 3216 */
128'h00000000000000000000000000000000, /* 3217 */
128'h00000000000000000000000000000000, /* 3218 */
128'h00000000000000000000000000000000, /* 3219 */
128'h00000000000000000000000000000000, /* 3220 */
128'h00000000000000000000000000000000, /* 3221 */
128'h00000000000000000000000000000000, /* 3222 */
128'h00000000000000000000000000000000, /* 3223 */
128'h00000000000000000000000000000000, /* 3224 */
128'h00000000000000000000000000000000, /* 3225 */
128'h00000000000000000000000000000000, /* 3226 */
128'h00000000000000000000000000000000, /* 3227 */
128'h00000000000000000000000000000000, /* 3228 */
128'h00000000000000000000000000000000, /* 3229 */
128'h00000000000000000000000000000000, /* 3230 */
128'h00000000000000000000000000000000, /* 3231 */
128'h00000000000000000000000000000000, /* 3232 */
128'h00000000000000000000000000000000, /* 3233 */
128'h00000000000000000000000000000000, /* 3234 */
128'h00000000000000000000000000000000, /* 3235 */
128'h00000000000000000000000000000000, /* 3236 */
128'h00000000000000000000000000000000, /* 3237 */
128'h00000000000000000000000000000000, /* 3238 */
128'h00000000000000000000000000000000, /* 3239 */
128'h00000000000000000000000000000000, /* 3240 */
128'h00000000000000000000000000000000, /* 3241 */
128'h00000000000000000000000000000000, /* 3242 */
128'h00000000000000000000000000000000, /* 3243 */
128'h00000000000000000000000000000000, /* 3244 */
128'h00000000000000000000000000000000, /* 3245 */
128'h00000000000000000000000000000000, /* 3246 */
128'h00000000000000000000000000000000, /* 3247 */
128'h00000000000000000000000000000000, /* 3248 */
128'h00000000000000000000000000000000, /* 3249 */
128'h00000000000000000000000000000000, /* 3250 */
128'h00000000000000000000000000000000, /* 3251 */
128'h00000000000000000000000000000000, /* 3252 */
128'h00000000000000000000000000000000, /* 3253 */
128'h00000000000000000000000000000000, /* 3254 */
128'h00000000000000000000000000000000, /* 3255 */
128'h00000000000000000000000000000000, /* 3256 */
128'h00000000000000000000000000000000, /* 3257 */
128'h00000000000000000000000000000000, /* 3258 */
128'h00000000000000000000000000000000, /* 3259 */
128'h00000000000000000000000000000000, /* 3260 */
128'h00000000000000000000000000000000, /* 3261 */
128'h00000000000000000000000000000000, /* 3262 */
128'h00000000000000000000000000000000, /* 3263 */
128'h00000000000000000000000000000000, /* 3264 */
128'h00000000000000000000000000000000, /* 3265 */
128'h00000000000000000000000000000000, /* 3266 */
128'h00000000000000000000000000000000, /* 3267 */
128'h00000000000000000000000000000000, /* 3268 */
128'h00000000000000000000000000000000, /* 3269 */
128'h00000000000000000000000000000000, /* 3270 */
128'h00000000000000000000000000000000, /* 3271 */
128'h00000000000000000000000000000000, /* 3272 */
128'h00000000000000000000000000000000, /* 3273 */
128'h00000000000000000000000000000000, /* 3274 */
128'h00000000000000000000000000000000, /* 3275 */
128'h00000000000000000000000000000000, /* 3276 */
128'h00000000000000000000000000000000, /* 3277 */
128'h00000000000000000000000000000000, /* 3278 */
128'h00000000000000000000000000000000, /* 3279 */
128'h00000000000000000000000000000000, /* 3280 */
128'h00000000000000000000000000000000, /* 3281 */
128'h00000000000000000000000000000000, /* 3282 */
128'h00000000000000000000000000000000, /* 3283 */
128'h00000000000000000000000000000000, /* 3284 */
128'h00000000000000000000000000000000, /* 3285 */
128'h00000000000000000000000000000000, /* 3286 */
128'h00000000000000000000000000000000, /* 3287 */
128'h00000000000000000000000000000000, /* 3288 */
128'h00000000000000000000000000000000, /* 3289 */
128'h00000000000000000000000000000000, /* 3290 */
128'h00000000000000000000000000000000, /* 3291 */
128'h00000000000000000000000000000000, /* 3292 */
128'h00000000000000000000000000000000, /* 3293 */
128'h00000000000000000000000000000000, /* 3294 */
128'h00000000000000000000000000000000, /* 3295 */
128'h00000000000000000000000000000000, /* 3296 */
128'h00000000000000000000000000000000, /* 3297 */
128'h00000000000000000000000000000000, /* 3298 */
128'h00000000000000000000000000000000, /* 3299 */
128'h00000000000000000000000000000000, /* 3300 */
128'h00000000000000000000000000000000, /* 3301 */
128'h00000000000000000000000000000000, /* 3302 */
128'h00000000000000000000000000000000, /* 3303 */
128'h00000000000000000000000000000000, /* 3304 */
128'h00000000000000000000000000000000, /* 3305 */
128'h00000000000000000000000000000000, /* 3306 */
128'h00000000000000000000000000000000, /* 3307 */
128'h00000000000000000000000000000000, /* 3308 */
128'h00000000000000000000000000000000, /* 3309 */
128'h00000000000000000000000000000000, /* 3310 */
128'h00000000000000000000000000000000, /* 3311 */
128'h00000000000000000000000000000000, /* 3312 */
128'h00000000000000000000000000000000, /* 3313 */
128'h00000000000000000000000000000000, /* 3314 */
128'h00000000000000000000000000000000, /* 3315 */
128'h00000000000000000000000000000000, /* 3316 */
128'h00000000000000000000000000000000, /* 3317 */
128'h00000000000000000000000000000000, /* 3318 */
128'h00000000000000000000000000000000, /* 3319 */
128'h00000000000000000000000000000000, /* 3320 */
128'h00000000000000000000000000000000, /* 3321 */
128'h00000000000000000000000000000000, /* 3322 */
128'h00000000000000000000000000000000, /* 3323 */
128'h00000000000000000000000000000000, /* 3324 */
128'h00000000000000000000000000000000, /* 3325 */
128'h00000000000000000000000000000000, /* 3326 */
128'h00000000000000000000000000000000, /* 3327 */
128'h00000000000000000000000000000000, /* 3328 */
128'h00000000000000000000000000000000, /* 3329 */
128'h00000000000000000000000000000000, /* 3330 */
128'h00000000000000000000000000000000, /* 3331 */
128'h00000000000000000000000000000000, /* 3332 */
128'h00000000000000000000000000000000, /* 3333 */
128'h00000000000000000000000000000000, /* 3334 */
128'h00000000000000000000000000000000, /* 3335 */
128'h00000000000000000000000000000000, /* 3336 */
128'h00000000000000000000000000000000, /* 3337 */
128'h00000000000000000000000000000000, /* 3338 */
128'h00000000000000000000000000000000, /* 3339 */
128'h00000000000000000000000000000000, /* 3340 */
128'h00000000000000000000000000000000, /* 3341 */
128'h00000000000000000000000000000000, /* 3342 */
128'h00000000000000000000000000000000, /* 3343 */
128'h00000000000000000000000000000000, /* 3344 */
128'h00000000000000000000000000000000, /* 3345 */
128'h00000000000000000000000000000000, /* 3346 */
128'h00000000000000000000000000000000, /* 3347 */
128'h00000000000000000000000000000000, /* 3348 */
128'h00000000000000000000000000000000, /* 3349 */
128'h00000000000000000000000000000000, /* 3350 */
128'h00000000000000000000000000000000, /* 3351 */
128'h00000000000000000000000000000000, /* 3352 */
128'h00000000000000000000000000000000, /* 3353 */
128'h00000000000000000000000000000000, /* 3354 */
128'h00000000000000000000000000000000, /* 3355 */
128'h00000000000000000000000000000000, /* 3356 */
128'h00000000000000000000000000000000, /* 3357 */
128'h00000000000000000000000000000000, /* 3358 */
128'h00000000000000000000000000000000, /* 3359 */
128'h00000000000000000000000000000000, /* 3360 */
128'h00000000000000000000000000000000, /* 3361 */
128'h00000000000000000000000000000000, /* 3362 */
128'h00000000000000000000000000000000, /* 3363 */
128'h00000000000000000000000000000000, /* 3364 */
128'h00000000000000000000000000000000, /* 3365 */
128'h00000000000000000000000000000000, /* 3366 */
128'h00000000000000000000000000000000, /* 3367 */
128'h00000000000000000000000000000000, /* 3368 */
128'h00000000000000000000000000000000, /* 3369 */
128'h00000000000000000000000000000000, /* 3370 */
128'h00000000000000000000000000000000, /* 3371 */
128'h00000000000000000000000000000000, /* 3372 */
128'h00000000000000000000000000000000, /* 3373 */
128'h00000000000000000000000000000000, /* 3374 */
128'h00000000000000000000000000000000, /* 3375 */
128'h00000000000000000000000000000000, /* 3376 */
128'h00000000000000000000000000000000, /* 3377 */
128'h00000000000000000000000000000000, /* 3378 */
128'h00000000000000000000000000000000, /* 3379 */
128'h00000000000000000000000000000000, /* 3380 */
128'h00000000000000000000000000000000, /* 3381 */
128'h00000000000000000000000000000000, /* 3382 */
128'h00000000000000000000000000000000, /* 3383 */
128'h00000000000000000000000000000000, /* 3384 */
128'h00000000000000000000000000000000, /* 3385 */
128'h00000000000000000000000000000000, /* 3386 */
128'h00000000000000000000000000000000, /* 3387 */
128'h00000000000000000000000000000000, /* 3388 */
128'h00000000000000000000000000000000, /* 3389 */
128'h00000000000000000000000000000000, /* 3390 */
128'h00000000000000000000000000000000, /* 3391 */
128'h00000000000000000000000000000000, /* 3392 */
128'h00000000000000000000000000000000, /* 3393 */
128'h00000000000000000000000000000000, /* 3394 */
128'h00000000000000000000000000000000, /* 3395 */
128'h00000000000000000000000000000000, /* 3396 */
128'h00000000000000000000000000000000, /* 3397 */
128'h00000000000000000000000000000000, /* 3398 */
128'h00000000000000000000000000000000, /* 3399 */
128'h00000000000000000000000000000000, /* 3400 */
128'h00000000000000000000000000000000, /* 3401 */
128'h00000000000000000000000000000000, /* 3402 */
128'h00000000000000000000000000000000, /* 3403 */
128'h00000000000000000000000000000000, /* 3404 */
128'h00000000000000000000000000000000, /* 3405 */
128'h00000000000000000000000000000000, /* 3406 */
128'h00000000000000000000000000000000, /* 3407 */
128'h00000000000000000000000000000000, /* 3408 */
128'h00000000000000000000000000000000, /* 3409 */
128'h00000000000000000000000000000000, /* 3410 */
128'h00000000000000000000000000000000, /* 3411 */
128'h00000000000000000000000000000000, /* 3412 */
128'h00000000000000000000000000000000, /* 3413 */
128'h00000000000000000000000000000000, /* 3414 */
128'h00000000000000000000000000000000, /* 3415 */
128'h00000000000000000000000000000000, /* 3416 */
128'h00000000000000000000000000000000, /* 3417 */
128'h00000000000000000000000000000000, /* 3418 */
128'h00000000000000000000000000000000, /* 3419 */
128'h00000000000000000000000000000000, /* 3420 */
128'h00000000000000000000000000000000, /* 3421 */
128'h00000000000000000000000000000000, /* 3422 */
128'h00000000000000000000000000000000, /* 3423 */
128'h00000000000000000000000000000000, /* 3424 */
128'h00000000000000000000000000000000, /* 3425 */
128'h00000000000000000000000000000000, /* 3426 */
128'h00000000000000000000000000000000, /* 3427 */
128'h00000000000000000000000000000000, /* 3428 */
128'h00000000000000000000000000000000, /* 3429 */
128'h00000000000000000000000000000000, /* 3430 */
128'h00000000000000000000000000000000, /* 3431 */
128'h00000000000000000000000000000000, /* 3432 */
128'h00000000000000000000000000000000, /* 3433 */
128'h00000000000000000000000000000000, /* 3434 */
128'h00000000000000000000000000000000, /* 3435 */
128'h00000000000000000000000000000000, /* 3436 */
128'h00000000000000000000000000000000, /* 3437 */
128'h00000000000000000000000000000000, /* 3438 */
128'h00000000000000000000000000000000, /* 3439 */
128'h00000000000000000000000000000000, /* 3440 */
128'h00000000000000000000000000000000, /* 3441 */
128'h00000000000000000000000000000000, /* 3442 */
128'h00000000000000000000000000000000, /* 3443 */
128'h00000000000000000000000000000000, /* 3444 */
128'h00000000000000000000000000000000, /* 3445 */
128'h00000000000000000000000000000000, /* 3446 */
128'h00000000000000000000000000000000, /* 3447 */
128'h00000000000000000000000000000000, /* 3448 */
128'h00000000000000000000000000000000, /* 3449 */
128'h00000000000000000000000000000000, /* 3450 */
128'h00000000000000000000000000000000, /* 3451 */
128'h00000000000000000000000000000000, /* 3452 */
128'h00000000000000000000000000000000, /* 3453 */
128'h00000000000000000000000000000000, /* 3454 */
128'h00000000000000000000000000000000, /* 3455 */
128'h00000000000000000000000000000000, /* 3456 */
128'h00000000000000000000000000000000, /* 3457 */
128'h00000000000000000000000000000000, /* 3458 */
128'h00000000000000000000000000000000, /* 3459 */
128'h00000000000000000000000000000000, /* 3460 */
128'h00000000000000000000000000000000, /* 3461 */
128'h00000000000000000000000000000000, /* 3462 */
128'h00000000000000000000000000000000, /* 3463 */
128'h00000000000000000000000000000000, /* 3464 */
128'h00000000000000000000000000000000, /* 3465 */
128'h00000000000000000000000000000000, /* 3466 */
128'h00000000000000000000000000000000, /* 3467 */
128'h00000000000000000000000000000000, /* 3468 */
128'h00000000000000000000000000000000, /* 3469 */
128'h00000000000000000000000000000000, /* 3470 */
128'h00000000000000000000000000000000, /* 3471 */
128'h00000000000000000000000000000000, /* 3472 */
128'h00000000000000000000000000000000, /* 3473 */
128'h00000000000000000000000000000000, /* 3474 */
128'h00000000000000000000000000000000, /* 3475 */
128'h00000000000000000000000000000000, /* 3476 */
128'h00000000000000000000000000000000, /* 3477 */
128'h00000000000000000000000000000000, /* 3478 */
128'h00000000000000000000000000000000, /* 3479 */
128'h00000000000000000000000000000000, /* 3480 */
128'h00000000000000000000000000000000, /* 3481 */
128'h00000000000000000000000000000000, /* 3482 */
128'h00000000000000000000000000000000, /* 3483 */
128'h00000000000000000000000000000000, /* 3484 */
128'h00000000000000000000000000000000, /* 3485 */
128'h00000000000000000000000000000000, /* 3486 */
128'h00000000000000000000000000000000, /* 3487 */
128'h00000000000000000000000000000000, /* 3488 */
128'h00000000000000000000000000000000, /* 3489 */
128'h00000000000000000000000000000000, /* 3490 */
128'h00000000000000000000000000000000, /* 3491 */
128'h00000000000000000000000000000000, /* 3492 */
128'h00000000000000000000000000000000, /* 3493 */
128'h00000000000000000000000000000000, /* 3494 */
128'h00000000000000000000000000000000, /* 3495 */
128'h00000000000000000000000000000000, /* 3496 */
128'h00000000000000000000000000000000, /* 3497 */
128'h00000000000000000000000000000000, /* 3498 */
128'h00000000000000000000000000000000, /* 3499 */
128'h00000000000000000000000000000000, /* 3500 */
128'h00000000000000000000000000000000, /* 3501 */
128'h00000000000000000000000000000000, /* 3502 */
128'h00000000000000000000000000000000, /* 3503 */
128'h00000000000000000000000000000000, /* 3504 */
128'h00000000000000000000000000000000, /* 3505 */
128'h00000000000000000000000000000000, /* 3506 */
128'h00000000000000000000000000000000, /* 3507 */
128'h00000000000000000000000000000000, /* 3508 */
128'h00000000000000000000000000000000, /* 3509 */
128'h00000000000000000000000000000000, /* 3510 */
128'h00000000000000000000000000000000, /* 3511 */
128'h00000000000000000000000000000000, /* 3512 */
128'h00000000000000000000000000000000, /* 3513 */
128'h00000000000000000000000000000000, /* 3514 */
128'h00000000000000000000000000000000, /* 3515 */
128'h00000000000000000000000000000000, /* 3516 */
128'h00000000000000000000000000000000, /* 3517 */
128'h00000000000000000000000000000000, /* 3518 */
128'h00000000000000000000000000000000, /* 3519 */
128'h00000000000000000000000000000000, /* 3520 */
128'h00000000000000000000000000000000, /* 3521 */
128'h00000000000000000000000000000000, /* 3522 */
128'h00000000000000000000000000000000, /* 3523 */
128'h00000000000000000000000000000000, /* 3524 */
128'h00000000000000000000000000000000, /* 3525 */
128'h00000000000000000000000000000000, /* 3526 */
128'h00000000000000000000000000000000, /* 3527 */
128'h00000000000000000000000000000000, /* 3528 */
128'h00000000000000000000000000000000, /* 3529 */
128'h00000000000000000000000000000000, /* 3530 */
128'h00000000000000000000000000000000, /* 3531 */
128'h00000000000000000000000000000000, /* 3532 */
128'h00000000000000000000000000000000, /* 3533 */
128'h00000000000000000000000000000000, /* 3534 */
128'h00000000000000000000000000000000, /* 3535 */
128'h00000000000000000000000000000000, /* 3536 */
128'h00000000000000000000000000000000, /* 3537 */
128'h00000000000000000000000000000000, /* 3538 */
128'h00000000000000000000000000000000, /* 3539 */
128'h00000000000000000000000000000000, /* 3540 */
128'h00000000000000000000000000000000, /* 3541 */
128'h00000000000000000000000000000000, /* 3542 */
128'h00000000000000000000000000000000, /* 3543 */
128'h00000000000000000000000000000000, /* 3544 */
128'h00000000000000000000000000000000, /* 3545 */
128'h00000000000000000000000000000000, /* 3546 */
128'h00000000000000000000000000000000, /* 3547 */
128'h00000000000000000000000000000000, /* 3548 */
128'h00000000000000000000000000000000, /* 3549 */
128'h00000000000000000000000000000000, /* 3550 */
128'h00000000000000000000000000000000, /* 3551 */
128'h00000000000000000000000000000000, /* 3552 */
128'h00000000000000000000000000000000, /* 3553 */
128'h00000000000000000000000000000000, /* 3554 */
128'h00000000000000000000000000000000, /* 3555 */
128'h00000000000000000000000000000000, /* 3556 */
128'h00000000000000000000000000000000, /* 3557 */
128'h00000000000000000000000000000000, /* 3558 */
128'h00000000000000000000000000000000, /* 3559 */
128'h00000000000000000000000000000000, /* 3560 */
128'h00000000000000000000000000000000, /* 3561 */
128'h00000000000000000000000000000000, /* 3562 */
128'h00000000000000000000000000000000, /* 3563 */
128'h00000000000000000000000000000000, /* 3564 */
128'h00000000000000000000000000000000, /* 3565 */
128'h00000000000000000000000000000000, /* 3566 */
128'h00000000000000000000000000000000, /* 3567 */
128'h00000000000000000000000000000000, /* 3568 */
128'h00000000000000000000000000000000, /* 3569 */
128'h00000000000000000000000000000000, /* 3570 */
128'h00000000000000000000000000000000, /* 3571 */
128'h00000000000000000000000000000000, /* 3572 */
128'h00000000000000000000000000000000, /* 3573 */
128'h00000000000000000000000000000000, /* 3574 */
128'h00000000000000000000000000000000, /* 3575 */
128'h00000000000000000000000000000000, /* 3576 */
128'h00000000000000000000000000000000, /* 3577 */
128'h00000000000000000000000000000000, /* 3578 */
128'h00000000000000000000000000000000, /* 3579 */
128'h00000000000000000000000000000000, /* 3580 */
128'h00000000000000000000000000000000, /* 3581 */
128'h00000000000000000000000000000000, /* 3582 */
128'h00000000000000000000000000000000, /* 3583 */
128'h00000000000000000000000000000000, /* 3584 */
128'h00000000000000000000000000000000, /* 3585 */
128'h00000000000000000000000000000000, /* 3586 */
128'h00000000000000000000000000000000, /* 3587 */
128'h00000000000000000000000000000000, /* 3588 */
128'h00000000000000000000000000000000, /* 3589 */
128'h00000000000000000000000000000000, /* 3590 */
128'h00000000000000000000000000000000, /* 3591 */
128'h00000000000000000000000000000000, /* 3592 */
128'h00000000000000000000000000000000, /* 3593 */
128'h00000000000000000000000000000000, /* 3594 */
128'h00000000000000000000000000000000, /* 3595 */
128'h00000000000000000000000000000000, /* 3596 */
128'h00000000000000000000000000000000, /* 3597 */
128'h00000000000000000000000000000000, /* 3598 */
128'h00000000000000000000000000000000, /* 3599 */
128'h00000000000000000000000000000000, /* 3600 */
128'h00000000000000000000000000000000, /* 3601 */
128'h00000000000000000000000000000000, /* 3602 */
128'h00000000000000000000000000000000, /* 3603 */
128'h00000000000000000000000000000000, /* 3604 */
128'h00000000000000000000000000000000, /* 3605 */
128'h00000000000000000000000000000000, /* 3606 */
128'h00000000000000000000000000000000, /* 3607 */
128'h00000000000000000000000000000000, /* 3608 */
128'h00000000000000000000000000000000, /* 3609 */
128'h00000000000000000000000000000000, /* 3610 */
128'h00000000000000000000000000000000, /* 3611 */
128'h00000000000000000000000000000000, /* 3612 */
128'h00000000000000000000000000000000, /* 3613 */
128'h00000000000000000000000000000000, /* 3614 */
128'h00000000000000000000000000000000, /* 3615 */
128'h00000000000000000000000000000000, /* 3616 */
128'h00000000000000000000000000000000, /* 3617 */
128'h00000000000000000000000000000000, /* 3618 */
128'h00000000000000000000000000000000, /* 3619 */
128'h00000000000000000000000000000000, /* 3620 */
128'h00000000000000000000000000000000, /* 3621 */
128'h00000000000000000000000000000000, /* 3622 */
128'h00000000000000000000000000000000, /* 3623 */
128'h00000000000000000000000000000000, /* 3624 */
128'h00000000000000000000000000000000, /* 3625 */
128'h00000000000000000000000000000000, /* 3626 */
128'h00000000000000000000000000000000, /* 3627 */
128'h00000000000000000000000000000000, /* 3628 */
128'h00000000000000000000000000000000, /* 3629 */
128'h00000000000000000000000000000000, /* 3630 */
128'h00000000000000000000000000000000, /* 3631 */
128'h00000000000000000000000000000000, /* 3632 */
128'h00000000000000000000000000000000, /* 3633 */
128'h00000000000000000000000000000000, /* 3634 */
128'h00000000000000000000000000000000, /* 3635 */
128'h00000000000000000000000000000000, /* 3636 */
128'h00000000000000000000000000000000, /* 3637 */
128'h00000000000000000000000000000000, /* 3638 */
128'h00000000000000000000000000000000, /* 3639 */
128'h00000000000000000000000000000000, /* 3640 */
128'h00000000000000000000000000000000, /* 3641 */
128'h00000000000000000000000000000000, /* 3642 */
128'h00000000000000000000000000000000, /* 3643 */
128'h00000000000000000000000000000000, /* 3644 */
128'h00000000000000000000000000000000, /* 3645 */
128'h00000000000000000000000000000000, /* 3646 */
128'h00000000000000000000000000000000, /* 3647 */
128'h00000000000000000000000000000000, /* 3648 */
128'h00000000000000000000000000000000, /* 3649 */
128'h00000000000000000000000000000000, /* 3650 */
128'h00000000000000000000000000000000, /* 3651 */
128'h00000000000000000000000000000000, /* 3652 */
128'h00000000000000000000000000000000, /* 3653 */
128'h00000000000000000000000000000000, /* 3654 */
128'h00000000000000000000000000000000, /* 3655 */
128'h00000000000000000000000000000000, /* 3656 */
128'h00000000000000000000000000000000, /* 3657 */
128'h00000000000000000000000000000000, /* 3658 */
128'h00000000000000000000000000000000, /* 3659 */
128'h00000000000000000000000000000000, /* 3660 */
128'h00000000000000000000000000000000, /* 3661 */
128'h00000000000000000000000000000000, /* 3662 */
128'h00000000000000000000000000000000, /* 3663 */
128'h00000000000000000000000000000000, /* 3664 */
128'h00000000000000000000000000000000, /* 3665 */
128'h00000000000000000000000000000000, /* 3666 */
128'h00000000000000000000000000000000, /* 3667 */
128'h00000000000000000000000000000000, /* 3668 */
128'h00000000000000000000000000000000, /* 3669 */
128'h00000000000000000000000000000000, /* 3670 */
128'h00000000000000000000000000000000, /* 3671 */
128'h00000000000000000000000000000000, /* 3672 */
128'h00000000000000000000000000000000, /* 3673 */
128'h00000000000000000000000000000000, /* 3674 */
128'h00000000000000000000000000000000, /* 3675 */
128'h00000000000000000000000000000000, /* 3676 */
128'h00000000000000000000000000000000, /* 3677 */
128'h00000000000000000000000000000000, /* 3678 */
128'h00000000000000000000000000000000, /* 3679 */
128'h00000000000000000000000000000000, /* 3680 */
128'h00000000000000000000000000000000, /* 3681 */
128'h00000000000000000000000000000000, /* 3682 */
128'h00000000000000000000000000000000, /* 3683 */
128'h00000000000000000000000000000000, /* 3684 */
128'h00000000000000000000000000000000, /* 3685 */
128'h00000000000000000000000000000000, /* 3686 */
128'h00000000000000000000000000000000, /* 3687 */
128'h00000000000000000000000000000000, /* 3688 */
128'h00000000000000000000000000000000, /* 3689 */
128'h00000000000000000000000000000000, /* 3690 */
128'h00000000000000000000000000000000, /* 3691 */
128'h00000000000000000000000000000000, /* 3692 */
128'h00000000000000000000000000000000, /* 3693 */
128'h00000000000000000000000000000000, /* 3694 */
128'h00000000000000000000000000000000, /* 3695 */
128'h00000000000000000000000000000000, /* 3696 */
128'h00000000000000000000000000000000, /* 3697 */
128'h00000000000000000000000000000000, /* 3698 */
128'h00000000000000000000000000000000, /* 3699 */
128'h00000000000000000000000000000000, /* 3700 */
128'h00000000000000000000000000000000, /* 3701 */
128'h00000000000000000000000000000000, /* 3702 */
128'h00000000000000000000000000000000, /* 3703 */
128'h00000000000000000000000000000000, /* 3704 */
128'h00000000000000000000000000000000, /* 3705 */
128'h00000000000000000000000000000000, /* 3706 */
128'h00000000000000000000000000000000, /* 3707 */
128'h00000000000000000000000000000000, /* 3708 */
128'h00000000000000000000000000000000, /* 3709 */
128'h00000000000000000000000000000000, /* 3710 */
128'h00000000000000000000000000000000, /* 3711 */
128'h00000000000000000000000000000000, /* 3712 */
128'h00000000000000000000000000000000, /* 3713 */
128'h00000000000000000000000000000000, /* 3714 */
128'h00000000000000000000000000000000, /* 3715 */
128'h00000000000000000000000000000000, /* 3716 */
128'h00000000000000000000000000000000, /* 3717 */
128'h00000000000000000000000000000000, /* 3718 */
128'h00000000000000000000000000000000, /* 3719 */
128'h00000000000000000000000000000000, /* 3720 */
128'h00000000000000000000000000000000, /* 3721 */
128'h00000000000000000000000000000000, /* 3722 */
128'h00000000000000000000000000000000, /* 3723 */
128'h00000000000000000000000000000000, /* 3724 */
128'h00000000000000000000000000000000, /* 3725 */
128'h00000000000000000000000000000000, /* 3726 */
128'h00000000000000000000000000000000, /* 3727 */
128'h00000000000000000000000000000000, /* 3728 */
128'h00000000000000000000000000000000, /* 3729 */
128'h00000000000000000000000000000000, /* 3730 */
128'h00000000000000000000000000000000, /* 3731 */
128'h00000000000000000000000000000000, /* 3732 */
128'h00000000000000000000000000000000, /* 3733 */
128'h00000000000000000000000000000000, /* 3734 */
128'h00000000000000000000000000000000, /* 3735 */
128'h00000000000000000000000000000000, /* 3736 */
128'h00000000000000000000000000000000, /* 3737 */
128'h00000000000000000000000000000000, /* 3738 */
128'h00000000000000000000000000000000, /* 3739 */
128'h00000000000000000000000000000000, /* 3740 */
128'h00000000000000000000000000000000, /* 3741 */
128'h00000000000000000000000000000000, /* 3742 */
128'h00000000000000000000000000000000, /* 3743 */
128'h00000000000000000000000000000000, /* 3744 */
128'h00000000000000000000000000000000, /* 3745 */
128'h00000000000000000000000000000000, /* 3746 */
128'h00000000000000000000000000000000, /* 3747 */
128'h00000000000000000000000000000000, /* 3748 */
128'h00000000000000000000000000000000, /* 3749 */
128'h00000000000000000000000000000000, /* 3750 */
128'h00000000000000000000000000000000, /* 3751 */
128'h00000000000000000000000000000000, /* 3752 */
128'h00000000000000000000000000000000, /* 3753 */
128'h00000000000000000000000000000000, /* 3754 */
128'h00000000000000000000000000000000, /* 3755 */
128'h00000000000000000000000000000000, /* 3756 */
128'h00000000000000000000000000000000, /* 3757 */
128'h00000000000000000000000000000000, /* 3758 */
128'h00000000000000000000000000000000, /* 3759 */
128'h00000000000000000000000000000000, /* 3760 */
128'h00000000000000000000000000000000, /* 3761 */
128'h00000000000000000000000000000000, /* 3762 */
128'h00000000000000000000000000000000, /* 3763 */
128'h00000000000000000000000000000000, /* 3764 */
128'h00000000000000000000000000000000, /* 3765 */
128'h00000000000000000000000000000000, /* 3766 */
128'h00000000000000000000000000000000, /* 3767 */
128'h00000000000000000000000000000000, /* 3768 */
128'h00000000000000000000000000000000, /* 3769 */
128'h00000000000000000000000000000000, /* 3770 */
128'h00000000000000000000000000000000, /* 3771 */
128'h00000000000000000000000000000000, /* 3772 */
128'h00000000000000000000000000000000, /* 3773 */
128'h00000000000000000000000000000000, /* 3774 */
128'h00000000000000000000000000000000, /* 3775 */
128'h00000000000000000000000000000000, /* 3776 */
128'h00000000000000000000000000000000, /* 3777 */
128'h00000000000000000000000000000000, /* 3778 */
128'h00000000000000000000000000000000, /* 3779 */
128'h00000000000000000000000000000000, /* 3780 */
128'h00000000000000000000000000000000, /* 3781 */
128'h00000000000000000000000000000000, /* 3782 */
128'h00000000000000000000000000000000, /* 3783 */
128'h00000000000000000000000000000000, /* 3784 */
128'h00000000000000000000000000000000, /* 3785 */
128'h00000000000000000000000000000000, /* 3786 */
128'h00000000000000000000000000000000, /* 3787 */
128'h00000000000000000000000000000000, /* 3788 */
128'h00000000000000000000000000000000, /* 3789 */
128'h00000000000000000000000000000000, /* 3790 */
128'h00000000000000000000000000000000, /* 3791 */
128'h00000000000000000000000000000000, /* 3792 */
128'h00000000000000000000000000000000, /* 3793 */
128'h00000000000000000000000000000000, /* 3794 */
128'h00000000000000000000000000000000, /* 3795 */
128'h00000000000000000000000000000000, /* 3796 */
128'h00000000000000000000000000000000, /* 3797 */
128'h00000000000000000000000000000000, /* 3798 */
128'h00000000000000000000000000000000, /* 3799 */
128'h00000000000000000000000000000000, /* 3800 */
128'h00000000000000000000000000000000, /* 3801 */
128'h00000000000000000000000000000000, /* 3802 */
128'h00000000000000000000000000000000, /* 3803 */
128'h00000000000000000000000000000000, /* 3804 */
128'h00000000000000000000000000000000, /* 3805 */
128'h00000000000000000000000000000000, /* 3806 */
128'h00000000000000000000000000000000, /* 3807 */
128'h00000000000000000000000000000000, /* 3808 */
128'h00000000000000000000000000000000, /* 3809 */
128'h00000000000000000000000000000000, /* 3810 */
128'h00000000000000000000000000000000, /* 3811 */
128'h00000000000000000000000000000000, /* 3812 */
128'h00000000000000000000000000000000, /* 3813 */
128'h00000000000000000000000000000000, /* 3814 */
128'h00000000000000000000000000000000, /* 3815 */
128'h00000000000000000000000000000000, /* 3816 */
128'h00000000000000000000000000000000, /* 3817 */
128'h00000000000000000000000000000000, /* 3818 */
128'h00000000000000000000000000000000, /* 3819 */
128'h00000000000000000000000000000000, /* 3820 */
128'h00000000000000000000000000000000, /* 3821 */
128'h00000000000000000000000000000000, /* 3822 */
128'h00000000000000000000000000000000, /* 3823 */
128'h00000000000000000000000000000000, /* 3824 */
128'h00000000000000000000000000000000, /* 3825 */
128'h00000000000000000000000000000000, /* 3826 */
128'h00000000000000000000000000000000, /* 3827 */
128'h00000000000000000000000000000000, /* 3828 */
128'h00000000000000000000000000000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00000000000000000000000000000000, /* 3840 */
128'h00000000000000000000000000000000, /* 3841 */
128'h00000000000000000000000000000000, /* 3842 */
128'h00000000000000000000000000000000, /* 3843 */
128'h00000000000000000000000000000000, /* 3844 */
128'h00000000000000000000000000000000, /* 3845 */
128'h00000000000000000000000000000000, /* 3846 */
128'h00000000000000000000000000000000, /* 3847 */
128'h00000000000000000000000000000000, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule

